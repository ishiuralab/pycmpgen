module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fcdd498b964295735d78bd0690ffd1bd66b5a806e83e3b53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a44a8b32ee2c2a5d889f0840f0f3f7446324075b9e9fd8aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadd6e9aee72e357ec0d34c7b113dca7216c874f012673c6b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7355cacf108548d52931cb830c4fb88ff0f15023b238ced0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ca00adaa4f54bf7ce35fa99162a8584c2faaa83de31b81a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f727687434a2478b47f908b4ab070707355567517414f8c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf509bbf82b2038e10bc6a643f179f0e0569a4e3b5246839c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bde5b453b0a210dfec2e96f3af4fbaf9ee1bf70bd75d1e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8acddd8bdff955b9e7dfe8be96970e28a47dcfd76c1a2c860;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b658dec18f39122366eb629ff5c1cc39f3559a558518678a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e1e127869655bc68994455b7b404f196c066252168e3dfee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd28e50013d152eafdd8dfbc5b75fb35f0e13c9388e0c3b53e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3df5de7b8b8296bdca67256b00ba5a0c0cdd66a691bab7a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc61fee0fd755ecb3619bc8b785a716e2725867dea6279f0b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10d70ef507ed79af81c3300cc88a8c228fd1a57b630fb36a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47fdbdb9e49274ad6ab28c266c0863295741533923076cdc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc6407aa8b9df059d870a8dc9241267564c991b6ae1b550b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7038d5a3672d00e196944128893a3820405466d1e044ccb8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3549cb78faa476bef65e7bbf0e17fac0d77d1be6663c06fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd5751174cdd3633fa22f83796d1505f27fc30c85144a47e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaac5f3ec733b15c68e7cbe3abd6b5b94ebb47a77b6ecfc12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h878e601b570895aa3b49c7419a4679caca82ff2d5feb0c7ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1db59cbfc817411fbaf0ff181ede446b9ca085664bf765089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9b81978be4cfabb8e49e375ef9e1d18f617362ccaff2bf73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17827b5245184bddb6d416db1831c5e16096dbfa34e3ab711;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d4af746430c9b1a8ccc654de11cf5241f1ce18e2525a81c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3079be402adcecf748677e5d48af4408e5bdfc2e107111e18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72d6d70fc2909ba83fd85312479c969d173262137e0dc3c4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h624de91c7ea91c57828bff7fc55a8d2c39d2f091ba45e0434;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fa4a86028aed19e5075d2a3b39299b9e4257c5b7b44929d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac5fa285fcf7301e7962fed4b2ffcbca8212fa45c8aa221d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5039e7d9dcb3acd194383578f06b317167b0ae20fe37f406;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78967b7bdee6fa04b644071f6ab5a7ab2eb5da204054bfc16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaa36387ae3051a4da965e7aa93ab6f9cf60eb3e1c8a06f03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cbd3adc94ec7bf45e0e3ada4591f782b712e97abb123ed54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37d89f4925a84d1ca36d9c7a8fc2d28452694fb37bfe016a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h105dfd80df06a2bd54724d2c572f15ad2cfed73731bcd6cc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67d48eafc07e62f6cfa2c27551c064c4fb508e50f0959ff62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h762e6806c8912014c002eb42487295241bf34dc71d6b8cfd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77570d8acfbda39045a9a2d2238f2e169a6b4f629d5c497ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88d8801c39372de50f60e778c33047a6b86c203e01f1d6c8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11616b824025f4cafffdf8c9d78b24090ece0b1559caca45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce8e3f89cd8d5593dedf90859a0456a62004396cc68bbea29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf292a4d59c4e978963d088809f7dfe191ea3cba1e09b0670f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9936a5cadbb95d60f30b492c822ee225acf7ebd3304eec8c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63cc9ed01c976c795b05fd559169aa9ca82c5f2d49bc1bd2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h426054df208b8ed3b42e980232a7dfa4eb9479414deba496d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf968583d28c1a6c23de797675c6424d03e0539450cf551981;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74dbf3266d0510dfbf0387e5b3e9eb9b9755835d3927f4a6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8479a02cd14c2bbdbaab49d28472d9078016526dbd9f839a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac28f9bb53753dd67a3ca8128ef2afd70f0415af0043cf816;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91b0dccb28849af1c7b60fbf313c785c1eab40d59deed02f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2bdfab07acd99366847b970bdd9ba585a5d1c497f2c3aa3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h549d0e5e80802ea4ccc7857b17c26a80c9002f494e122036a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf18f9ad32774d51390de70a04400a83499c9341bab2202c4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb83a99bda5a6c20e10496ea97f389f453d2a2566d6e82f24b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdb3afc9f1b1a8762c07cff65414fe47413e630b355823301;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32f0c0258231a016cbcccf0cd9bc651e48502f5864a5dcc50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3799e84c58091be0e370f83a0504591b9ba8bbcae5de365c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha432b935151f3f5849b0bb33a8db2ef8787c739e8ea85b9ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bb8b1c587e49997091cc6fb8fca1621e2490c69c5becdb6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf124f39bfaa6fc8e373d6104f417694bd7683ef3702a1f8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26f227a2d308fad9125ec6b73bb200310cf5971240693055a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45c11cc6e851f40c453ffa989f9ed963fcf9e809ecb626482;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he22bfd70366bcdf2cc32d135eb85b673ba6338c7debc8dad4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72774590fece76f7ddbacf6f6d8a77d7434dd092bfb0d5039;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fa17ad4db5cea9de012fd4d53f9711cac84c69e13765eaad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98bf8f983f38ec139a9f354a09e77532dab7a5e039b2208e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa139ee89eb0b4961bcb77d8dcff44b3583806ffc3596b2fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h826a670775730d60a67118dac24d62447d08597890c08652a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc193d45efa773d2ae91f216a8721cff5162c1e7e9bb85e3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb85c8e64b8815a1aa89b2d6ffaabfe9371e59ad121a4f525;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a757ab5d6ab42f39989e87fe80db857237ca855eb5a297d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63a4b673e652e136afbca9cbe616b30ae5e50ac09e2ad4e29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc57aa3a77c90f6c80ee2f4d3455da0a43631bbcb16142f0cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc59eff7c2904fa4706badb7751be8385e2baffad7cebf9de4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf10ce333f59f83824e4d914eae5a80fb487d6a6e48b41b38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dfed36218dffe6df77f989854f484f487a4f39d185c4128f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa9822a541362f8b2635388d7a880d4c934db691039f513d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4e663212d6acb3955e12048e2e28ee67c6733d55a9fd2f48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11f2d99df44a2524e6addb0afcc19f91ca87e90a59c096c1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha348dfd1452a9133d87e6d5d75f57a96a866827b29bb4f689;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9560a8ba82867244a5947ca15cad40fb3de1ab9849283bfc9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfaff9850f89cfd4aad00c8055b57bc38428d6bc02fb28edf6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc31663093adbe11406ee1da8c32f04b71e6badbf209906169;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6253b376bd9d987d44e610cdfd900da06619e8bc6c298f09f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h990b28f7871ccf3db9bb301129343bcc1e41a221c8ac41c16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26b61ff4f9cc99bd72c54b0b1e168bf19e746e5bd1b8f0cc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d04a2b477d176bcc01f81670ed0d5343e48e18558abebf0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5868e377f2a9ad208a9f3bd53e6ad377aaf9be02d22efca12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78245d5408e98b9d43affba6fca327232d989e6568323387;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1948c984c8b97069c3c5af1ac5a37a02679bcc230ccf01bea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c356c0b889b177728aac2d3e30ed1a30df8c45c62ff0d9c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9af188e1bf0831c1f51a2134e84ddbb7c0a4299b7ffcfdf5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc15ea9a82a014d98ffd297fd41b4b81bc5eca9c053a5567c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ebf6bef235e64583b76fd0c3b778fd3dbaa7779f350fce0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bdeb573e2df0b4ae59277804e8142740dd4997e6660c6b68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h826db3e141e913694a9f0e31588fe3f8b2ef22625ccc6020a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc46de51d652337d1fecb1dd48331eebb12251e691a1a20867;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2755886734ac6a7167f1d403e7391e97fb536587646d66868;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h976bfbec13f649cc8e8f680b53f237a65994b8863e77bfbdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc0edc2b38bb3012243423e37f307ec99d6fe65498f0f63e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h598233187d156d158a34bf09bc27e473f62d5f01337996289;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd51ed480970adea96e87bdb9d61da5672405cf9eb2d655de7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4892c1e81b9cd529762d99542184d104a3fd1648a4567549f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa45163b19ee103e6744f36b38a1273909f6d31bd4531ab66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71eb63fb5f474564438453387c63a2910f1eefcc2efd9b146;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20cb0682c912efd5cb192113c1e9935973c94f56c79304d31;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8a8a01dc971e7428e56c5c11dbf4f9b56e647040433bb864;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f1a140db2f6521549ab007f09069887cbec3d78810927ab8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac3451b99c6ed67bd4efc8a3ef303d5628e6a6b1b1101af6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1faf74c8878d2b90722d59c46177d6460014fa2385a2e15ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39c00517736fb8f9a72e04dbfe46ac643696857809d6de9c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfda9951d4b0aa5619234f3e5387b8613264c367e54ab3eb68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0a231b630010f753b6b6e9749fed8f9eef7d898e2aacc67b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h531886144a7e901c0e6afd429b64ef541bc348438cb45a1ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha135206f528888f2e2380eaf3935b85c8a9074dd9628e3ee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b30f53c4e52c727b6bef31195eac422f10b12716300e3df1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49778ff88ead4f6dc791acebfe955ba4b9338fdced1dc8961;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32c83104e281341156529e74db4310e910d7acb5b6401d7ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h707099f361d1c0604133a75d2e144decb83c2caf64d1a7e00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aa83f5f33f407369da11e1443256336752779025c4b9cbf7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47c51cc9480c4259843061a10db0a22da56e8d1df8e3b575c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76662e930690a6247d0db7097f7425b0c35c0bd370d85e2b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd59e0b33207cd36a5d7501f32d73bed59b06fb1c6866c15bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h953abbc0726044fbaa38d1dfd04c558b0b344ebeb90d0d6d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b2c80f67f9f0416c66a444071e57a2765b497d2d3455e26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88eb7ca9d53539a5ea49424d47fcd1c665d0ab5ac3b86555e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f7c02e2de6de79a6b7ee6836870719c6fe148835733fe822;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd946c8ecd3301c40d2c3ae623241cd50a3c710c40b3fcd343;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd941a4bcd775f847be787eace38877f4fd6b63fcd3d93545f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8262a8ffbe4a4f7eaae653e724fa5887e0ba2fe07d154d3ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33a5c1e3c81a88334e01f58cb712db940be781d5e3ed8f20f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1485f849cc28f9c1b8fd8a08b38e40f9053d0ef9b5cf6bbda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56413dc46d68c0a341c9b510fd9fe77a6d036393beb169754;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99b8a7a1a90f1a259dde1a241ec423a9877937e93cb678855;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac8697b23b7f17dfee2308a04ce2c0f5d3d015915df965aa5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb58ab6edcad031ef4ce66211e46a56cdff32a195f16f28f6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1448a4a93121cd49b2898fbf641114f0716e648a3500d7bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49006d3338de656a292b2825c97e9c2c1964115fdee33643c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77083142b7aef5999f3ef6adfa0a1df26a6908965bbbe8a41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf007c8bc3292940ac687bdbb91e4ff8c3a21a6a993c23ca67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5ac776e324886678cb8fd3d0ce758fc5b65caae0c2750030;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e7184266589bd7106d58aab384d6c5ccc0810a1c86f79c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2152124a0124bb2a0926eaede37d5ea715b1b949fae0fb61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h105f0716fa1de6d4969780862e9cafce7acf1eeeb957ef239;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38d975bd4a5c5542be8546279f2d7888647cae8f4a6d7ec9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8dedc3f22fe2da0f5f3f667c9e3cac0f2d20c03e922139bb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8e84cc698738819a1b59e3cbd15f1ae82cb8462a661c36fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4f8793146483d51a95b458a37a5bf9954aa43a6be5dd9814;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71621bb066b753c74822ec9ff7b4ff0fde3bb01501150a87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae9b069a54f60a357ba64b5d7074be04cba69a89d5b93aed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heef64026d116a050e36bdd84d16453a8e30852863a7174b84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h917bace61f7914d5528ffb99eb3a1be7cf5a5f0b17d03eea0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbaef9e881489b412d83092d8a5d6b0099c95d749b99c4274;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ccf0d6b5d66bacdacd971293dcfd8ea56705e019ab5133f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc699706dd4103ce21f716a4bedb9f661710c3752ff806473;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4615b7abe6083b6ddb918552d4777dc1e059750c2b5cff63c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h651f22e7fc9c2e3605756eb4bef5770dd9b45e5aa76049c82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62b1d1ca23b3f821059836a8575a20a8b20d00a06a5ab4860;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1602cf13aacb85b83d36f8af44b0c58851bbdff3d93257ac8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h507b74a658bac77ad71eb81ea8077f2c01365c3bfe1938569;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1127a5710755e9242366c43c6c9f9272c3d79e833b7bdf935;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b7c2c9f0e88cfdf26b6588108ba7bba9e17a613df7cde77b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf56850c9168f19852df3077d9f7ce29ce538cd0842c87be4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32562c70b79c93536d4ee14d8222a266a0a34efc0ca306474;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf9f0a9d46b49de4ab900fb48a2eb36ba511aa971a8b4ead0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88cdeee52abccab9955170a8a535005708c888f4c72a66082;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89b9ea1eb10658e9010ba543033de423546c3c658cfbf0ede;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca7e342f954ce16ec98d90951419d85b89c6d82ab3b0af9ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cc775b9a47ffad3fcd53c81fceadb3df9d9dcca966d0d071;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81145ebcf2ff2f7b16d57b2449c1fe9302507e6866c6f154d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ef58c968cee211d2114bb070e16f6eadbcdb900dcb33379b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa1c13afddafbcb973b8859af2293162d9255d4b109272f51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cd654e480542b0323eab326497c62d8e583b6cb0593d6a30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bba9240f948448ba584c2f5ef30f5fd79ab08ea8ea72674b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd78e15ca4761a06dd8a0a87f8eb31a3a904818f4a16f80285;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86ca35e52db233e8a7ae2e4f48a600c5a8d64142f16fd1595;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haac20eb869cc0c4723b8c8e160674918298b344c4ecd65cef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc51df93fb1baba5d5cf14d5b38ac0abe1e566bbe9ddeef7dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4d3a14ab4488a3abf0cc4893f61463e73761647f07cf0ea1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5240b261b050237a0dfca95e2d2ac6a6e2bf7d7ef963c2794;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a741154c1875112217fcf5db31f85dc87bc48326f5b5c1fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f734e9ed3da41b1df83a575695c766e62800dd78b23cb3ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcabfd26ceafbffa492631d9aadaae815205eaddf14a8f65d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h359d8e881fe7c3bc4f41b2e0c325f9a3ce2c851a50f02f0c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a299c3910182eca2b27c3183f603d52a30b6a9f65edabd94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63e12cece9bff02924d9fc3e90a21a33fa370565237035173;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9690444b3443094fac69947ce786b2261f02a1b59a4a80b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf03865676b670f1cb2982c17381006f66810a89a757b91aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc078ddc6c5c4d73ca74629f450c783994b3eff0dc09a4363;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35125b95efc155637c494639e2339dd59293e492592ced18e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf3615743fa50b3e1e462399d42940df2f7aa1b9b3362d373;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e58dbccf0824363509d6d41931e5b7ed691372c38f5da936;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39cd27e348373f8d1f6bd49c213603f4685efeb9824d955;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4a9c907d1d3356fb776d835996e917799d8346fbdcb5971e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8121be80c5421c3c4837e744f8296a983aa7ef3c34d37af2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65a8d3f8d7fe09f61e19dbceb05df6d756f5458bade5d01f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1510eeeb2b9c6c735cd467b3b2e076716c8d53718a337dfdb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b7d9e04ab3aea4534bc55b59766a655f97b0a8f204c8af0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2269a862ce301a43b0d5947a67fda8626778749b23d1e240;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf22a5012c02582a59ed9b88c951fe4517e82f7a4c5d71cd01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99f6c4c20eb5ee5b88171389895858d21f82bfb6d3612e2d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9e3fbc5df8d36c263d7d0e826cac9866e8bf7b52d3193c9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2c7bc402d5eb12786f381003ab4c0aca341d6edce520111a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ef24130afd215eb15dc50eb73607d3316b0af8101a8642b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf08430f1b97f8ea4d0e93b7e63539ee4dfd46bc2bb12ffa1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h981ab978c06bdcf5ba0a63cd81a148ca5125c9097556736e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74c7ee2b7751b90adbdbc66d280a85946919b2beb8e29edc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha29731d8c88c626daf0d443efb93558dc0d79c1336667cf6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47f64bb950b409abe2defe3e97d23a9c6e98b97bfe75fa379;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8983f69d90bf487de71ed0098d3ccaa88005bad8519055613;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha881efbd823701337a366e00d345efbe68be74bfc7287073d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed07281597da0916a8aa8ab7e26717ae0ddec063a04a7502d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h965e8174dfba80f11c3e5f44e8ddfd8b44633ec4a09087272;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e297d6f40daf4c2a5c9f27482475924e207d3b12c5d2fc76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9df0afdc14eacf05f935eaecbcfa6a3ea76c8633380acf585;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e8b13c973e2a3455d8b9bc6cf19e7fead0a2b9544b3665fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30224d1b867dc2e5d7120b739ddb1a2a08f7ecb078edc9d94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb406111045dd9ee7a9c0098d5c8426ff67a8cd90245c0e0d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2db4fdc8a77880399baec624ec456208126f61688c8ada5ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b7d03e3fcdf40be52f05d33ad65a804b6aa57f9caef7f098;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53f9def9fc151675c1a93973a776c5209a007ea9ee2efd2ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88822826f1526bb51029aad2a457b84b8581d5dea88496194;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4bcfe252267ec100e02e2c39270eda0c24e5c1a735463683;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9492d155a6459e185147a4351433cf48829ab1f10ed34bd11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8ea1c22a3410130578b3078d1211e8941da1a8f5d1c50f27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc8867fa0bcf4a55167bb6837caa1fb2eba58515c52d61d81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce6d511d142b37fd45131b624584f59c01560f7c3710a7677;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45d8d239acdda9fa8fe87ed51f44c94607d159a6d77e9f5dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70bf24fef0b3351010c5e9b3318053a576462020a62b697e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48680626a770ccc5a3039a8e4d41c4b4b504d1201461e4b18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e5e6ab8d83cf6ada2c5ffd1405023a7325d90700d6f33464;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12663c63fc4f00cda4eb2d2b64d847949362aaa3bf01523cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h261734a1cf48e36db75fc737e54ba37009666db5b1816d176;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h109f3c239eeb9d8f5bdc52712fa3d2374403cb514752a73c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd010b8c5a0918945167148b800c9f338a7d96d3f68905510;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8ea7cd04c64fdb6225f6dd45af6f8b42ea6b929e461e31f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22a12c1c664b26b07d83a4a54181551eb58aa9cb9f82cfd40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27231921aeb59c3e41ed2d4d7c9ad7cf3f15cd593ef194a58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb0be0ef1fee0764bbabbcd45c492af55a62f3af132679c6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36d1f36cf1f0ebe08ef2e9ac4db2edb84566d97e9c0f1fbdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefff6ba9f5295ff324be8d7dd6784d30783363eeea6dcfeab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc43e8a1f1a1ac8a9b74cf5d7bfae613fd4068f56b9ab5c4ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8df7dfa61ee6ac8398c18d7133f7ca3fd86c75a07c51eaa0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c974975502c380a3cc646d965f5798d78882f903f61a196b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b1ee5ac5d7be580f549f27d1f824a1a6e14d42ad8f459834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f3233cdf472a5452e7c003ae53e0c555f1053aaee2410766;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee5662c3c1208c7644edf3ff57b16d29fd5b2a03428b31f0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5f25cf0c757ea99b101eb001ac66ff3fff081c691103f58d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d34f1d4f7de17f86ffbed546573bce3e67c12bed9f4f40d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e2877dfc0d6f178775f56f4718e8798a37a09007d206839b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b081d076c6e0e5f59519a3caaa437836453a2795eef10737;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hced304db8cc7a60ec57144d71c16bd8b5d372c0452fd5f677;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8959e2d79fbe4783442c985c64fcf0b784ce4cb48a5bae1c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cf042f5d3a2058b6e10d8da977f744e5b82e39a31991689d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5865d2ec1be2c3bb4c628dcd8b0dbea85d621bf600081d99f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b5f7d62d21a530798e58b597959c838c6c9912f01db9edd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b702d8cc5ff563abdcdff2f3c123642337a87f988440eb3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf566f2af6d6d7e9c47228c33a213bb4f6e104f32501117db7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd22b189a673b49f21a0feb0a92e19297802add7fef200107;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h565785c52c357c140e0d0c6091a25e50a375332320d408ebd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h883cc703b79e6c987212d03a10814624f698fd2382f415ea6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bcb26346b0df20f4641349577e8983a1031dd39a0d6bed3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc443eb7e5b89b5af574dee38953b4860ef22a1c09e4b719f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2dc6287e268a3133be831e49b363d9990e67416ea40a55b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5405e11cb26cb00fbc45b0cf5a2a76c1f8d92d1a0a9cf2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha42a2b2bd9ffa659d31f481d780c5e25d60cf84b70d671a6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3af0cebfc89a2270d64aff65bf05564e840c6ad572e792d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71d2c50d7b692f2bcfd047db0aca499032de5d92f7c39fa51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58b08d1e0786bf46dc440e2834886734cb13f53f567894fa5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfb3c73e4d000ae067e894c715e9c66ad8682fc9d5d2cc93b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h151b3b259d6c879ff4ee2ba43bfd120d06186d532c15b8b78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcb512150775625a9f6d6e3be9f8b073ff79808a56fc38ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7d144b102ad070681403cf44a3cf5ba18b23f76174ad0925;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8524b7e38e459359534028452cd5e3808fc1d84db72bf2c29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h124a6071167911a74cfbe1594005a47f7829829b176559064;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47485061bcf7dd51bdc94e11d224c0459fb44e7ba829362b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cc29aacf3743a96d8980763e53a98a7d662678f5f8414f9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40351043a658d249b0a77cad0cf077331956b6c61995c0e16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5d262c00cc05b7a49e8e01034f0548c8f7d201913d719a30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd668c98f254a232868b659493ed9314248a6fe8e8792b3d58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fffdf5420d6209ab7152a266e2367860f6be04c52bf6be75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcccbb6517d00059ed386edee3a320b67c4b52780906e28142;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87ec84df07ce309f2f86524a2ecd9f93179f44abe7473c966;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe2c9bb146de5d4da440056369f5165886d169c7214e4d227;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbeca1bb84008ca52761a16f2d02d01548b0d30a2baac535bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fc2a55bec550db42a0468271718ddd20b5f168a7cf2a14fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecdc600ab597ba053495675c7bd53b15139f8669d2a1061ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56a23576d76b4d2bbff0b56f78806a1b57ecab3efb01ec06e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb572e103db4fcf3d1b94f27cf9a04b9ca853d0900df5586ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h533dbd1b9e801236b1190c897e31c72749050877acb5043ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3b4699925efc95b94665355c2af36c490e7b0ee803916a02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab356bd42a9944b1bcb61882a4b4b1918e8d08b117286a245;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74e803b7241b0eb652575590d6ae2ad934282495c1506625f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f3825600da589165f52382fea56e475ca00d1030b6ca37b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ea12b2a24634b1ea3a483da54651c7bfecaa80b206ca3353;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c02718f22c00fa5fc8d421f8c7be64063f53fd58a13e1ebe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h997ed61659b9434aacd7cf2ce42f3fd1be068e05e3fba81e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h258f1f3c1702374027b06ed54cd430a1a9253bb617338ec47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85df0488eb45f13833da6e327bac0c773ffae37f3be1fb097;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71671998fc358e565ccd3d31a9057911fcdaf69289de615e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40cd743cc9005bfc592a7ee44b8f735693ffe92a2583ee1ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40012455ffde74d3ff4dfe452ca303c9f0e1d4331ddf766e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf74ffce9eb87fb91cd1b6eb83cc3ffad340a0b953fb38d19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7def701d8e91cb96eaebbb1e9e3518e220d20948899d8b836;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfd9c265da266d8c80906b35df9e81de1e14db99897abd41c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9b0974a3c850785eb787d97d14af26472708e5cfe995d3fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e24eb9414234d046a6e86993b833716f3e51b7866605814;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha482eee77f6f1f6110f88f5eb171258ff7e0d18362eb27540;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he64372c0e269de9dfce53ef721f626eca506de92b111a70cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b2b550cd4c34a6e5a8966eed3e381eeb966762375d96b711;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf15fdc61be55081122d4fff1c40f6a859a2bd2a1d0a7a534;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h800384392b6e001eb89fae0555c45e2a83cfa06e4e338d3f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h781c2a5e9f5a78a4570d247148024f734ac15bb7c144e755f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c313f1fc84c85b0cd3b4e2f98b7fe48ac4b83f11a85039f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6769e382f20134942615dbc1349ca2283ca4c20635c742759;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9be38b9ecae8f7558b48d4614d48e37d9471401c81f1951a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h367d5e2a965fe69e4a919a4db5495feb3b6fd40c36e7a5bf7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f6149a13ae52ba466b2f78f2c2ca90d9691ffc64781cd07c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb590611988a92a80fd485cf11e1ac6c560757f2a070c4847f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h761efc90cc42e7171b113facf07cc1f8fb5217eb07bae530f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed0017e269960091665f6353840475996a6d5a02443b73878;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b39394e5814ca04530c34ba5e42e973fc918aefde5e71ed7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c1903dfc88964569a94780427b482a2bff933b65bc2a15f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b38e855fa83dba4ef1d78067b9342ef7c4906b379cf3dadb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75232616f2f5ea42451d490fd7c01a77b77dcdb9a85e8a56e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h717bc1de7178f1a295814890ea081b36310e116ff8c188b81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6870b140b4a4db301e1b4490d0209ef4ec9fb63860bfd4a61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd69b51192f14a9351c82a7207621d2cbd60fc19ab9c04053a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dc83de95d2ea01325fefa5f6c579861e59026a654bf17675;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5fba80d2613c1d99ff6a76018e07249f07f3712c986d46fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2d21188f09bdea7e97fbc8d55f5dcc490a8ca157d1af7652;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6345c942fd1aba66eb099af8525372a4c1fd8ba876cf14c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa8cd15106742901073093f17fb106567e23aea6e6d8b4d75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f3cc0add01a89c29606cb642dd7e56f6a0eb67ac06d2bda0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5d361033837cf6461126c5bdcad46872c6f6733305bae775;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70b804457a1c2b5003306764da0378b4c0a3c02c1b16ea786;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49c207136132e6e8fb445354bcbc1a4cda90faeb1198d3ca3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce07a5b6295675b8a87b5d0a2f0a76b11b0a24b788d832d6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ebb151d59e958c747c79fd1e395e514591ad243c536d4efa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4edb17b072b203a962680bb3b1574b47978c239e95ea4e07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86e5eff902c49b523c38e4a9c1613b4c04ee311dbdf09c926;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d001e5ca00f413496d29d3951c23d61e9a67ab13b2d9cc6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f4d143e3e3c9c8068723b4c48383204c1fa5ed58e798d209;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d539359d19aad3b311b69900bd6f4d550e46be26e007b9de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb909900a3fc42740c1d6384435e221c6d22de4ff11dec382d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h300f837b06d64279e178479cf888118b8dbe51f237a57672d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec9041ddb87fee1606a880a70911302a08b39dba3c55e9486;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21f726537ffc7a2c2d2a9618a7c205251d3f31d2934ee1602;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h665e7c2d7814d8e13701c8fa482dab647201a9c27bb67565a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd6d7cb8c6e1704180bca2bd6349d9a5f051fd3f8a215c30a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f936369116f2f6c87e858aca81bdbf308f2c37d82cd62908;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87ab5c7cf9548498eff8d317540d88f6c97b3231e271f0392;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b67aefe5a3c0cca005f4b378878d43d591dfda124fbba2fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb61b2c042121ec82580784bfed7c4ddfb9a3f9e18c6e004dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h537986d475b3e12bfed95012781e2679b0b4603d034b1487b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha08d6ef0850b3625b07852c06ee2e781f41e634421ed867bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cf2d4dfc2ca2dcf1ea661a2a0373ab67c774629dad37a507;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha260fb2ff33c925ba226ed8ee241935533e63031e8f25d284;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4c1e835f7e72e2591304aa9daad77e4d841bc3c86e58e461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha211480107c1825990e40ea95706eb7ef34d1c17be2bcf2de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73d60a26506946096228399bef558d0fd84aec49c9befe030;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd054c13192df6d065729b9af55d0e3a21b8fb0d274a332117;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a1a0a415fa5cad003f0691897797ec2a08e490935c51c706;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95fb4324a94125c7442d7f1cec250c0cf0691dfeaae8ce8d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha790b6a8d800f2463a1b31d274d9a5f1a76778a764933154f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d00f0a5c32867144417b7f9a7c5b9fb738afb9c4893d7461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf62bad87aa803606368fed5e155a11e97fece4e84ade8d972;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcaf3d0f77e73557378fc45bf76da02419fcf8f37b6b5eb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61ab48a595cd7d30d6a0158c84b8ee0e6085a8a425719a2f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c6a81bbdb9441a7b994050f6e1851a7117780d6bcd561dbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d03ad2ccaa3cfa7136dd7f3e048335f634e8438c0d4a95d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69c87b4487492cc1927bdac14cd4e7cf64aa0c4e42b8bd52a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb430f3d2c4a21f1e2f0536199a8a5813d88587a805e39aafb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6376bc0bbc5decedc91f98a7dc9952ea0496684da09c8b64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0024e404512c4ae27a819b5d6870ad8a3058acc1776beb67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab5564c4a0f06e4c8ecfdd5c522a9c2b8cd1a2250033cae22;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd133335ef87a3cf66062624cb713722f75a6e0d66d06b0b57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57c0dddfa9ce742ada040c5543641e182f91cb94dfc25a581;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcfacc9fa89233b435af42bfb6738b65e2316567eb1771291;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b1ffd93ee40bca5353b36c6b9968bc5cb5a479e7025839b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h913c2ec9f942ef144c78e157631bcc36720aa006ee4c3f125;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbd9497f1096f247e3b08fae16490724434d4218b4f0268af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e5a0b84d9ad132b922d3f3ed8bd8bcda4b282dce75dace5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71a04776930fe26468bf4da8faaf711fcf2ec14eb68655fbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cfb851f26e223bfccb6ec584a73994e3f9e4ff596fa1b275;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0d4ebc2f9584f8bc7630a219d7b65435b320f6a97ec9e693;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73e1d2b132ceecb62ce266079804e49b3a7e6af36cc3e5626;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0bacb2bef9c320c52f3a47fd40adfaec3437dc24ed3e6073;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec2c290a35378c0424f3c08e6f2a825baba65d05d139a4d61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3adb5b43294a112e4ad825848c6a67e16769271f35416a1b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68b3d3db11179591fa3502b67032c92235ddd552fa3426700;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c4e5e11082e83dafa3ae2c67d62bbe43f715cb2faeff8aa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4eda59610d7a9708cde8f6c746551d46722be6e70c0b9549;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h774412b8d9d97b8ba96c1269d82bfc8cc4ee0b86761d84ceb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf407caf1f485e065c5befa46d4c54ef7562a03b36d923a4a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf2dc1bef79939ab138f010ede76dcec3d05dbb74bad65ef4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h981c6ccc7f2355c949518843269e2f463f985f094cbc41069;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h327ac279edf86e753cbd001a433ac8df92c6abb8db9fae707;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd5d46a6df9166074bbdee08dbec0d623a1d295a63afc8a1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5c569022a37f27003892e6022fa1cdc663910ac14723153a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde0d41e1ec37ac87be618401ac90e34169ff4f6a5301b1152;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcae4f49fd1a9921207d24dca3fb9434b54b8ec36329082d37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7c6f917ba0f97748cb4ae0c3b9b9b09fee348279da047aff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec17f920521c5d2eaffadafeb4e0ffda67c742311c9f14b60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ecfc0338dabac60d8acb7ec9e7566cfe8580f6703a6a1e67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd011a8cb6fde058e47b2c4fa6d70fde3ac51688df7d8acd7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6d3f32f3bd77490b834c115dcd1ca627a1b0e9b4fd0e32e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99edbab68bd9b542e4042cab0387f44915f964472800cd16a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73d60e1b562c8d2b977992d51121a22fa37be77d1623d48a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29954cc0a548062479e6cf10d2c08586cbdf467ed7bb10a81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb05c97065816e5d657a93f15bffe613a97bf6ea12fd1ca3f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fb24d3a9d7b24ab514815054a2ba25b4da1c5b25cf8d1cc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730a11703995171a1c5e3f757510d294b4eca72be19841b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d1e40d840b2ad4e0a896f8be637a22eb695d5c0fc638cbf8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habea8607df68c2cbe32a87911152d4810878727f3de1233b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef3baad19da80ae272877c11d30b10e604b0eb0c6d1c007f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44860a0a92be15be2a4abe2ed5edfe3441a06b30005472ba7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h190cbda038a4b0a19dba7090765f94d301c523161e584fd4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf6b0ca2ce77295c15165aabed649f3b0dcd514e75ef1a8f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf502fa7de3e8e2112e60982336a7f299c5c8fb57f9040f7b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47d1f80a3bdb396295ea49813c96bb8114308ab36b24f576b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h536de119eda2e8ca92bb19d478cfe12983df589cf6aafac6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb024e1993ddf349db9c0e5b1140255c5b9f6639db4eca00b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80c9e793981351f6b3fb43e655a93c52cd0369f3eff543c33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf98aaf2e5d4ed504d30a0f8db2af9e791ca5eab10d3bfe8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf212bd1357d004bdc38f68c5db543022c17f6b86f05535532;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46c603fdf8146c7d3e1b6624b22cca02af49897dd7a798b3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h858c5ad4e68bedbc048fcf8138a63dfcef9d285e90c118896;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf55214c0bfbefcdbd50882a40c26f1591682aba75ec908316;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h183ac9de980f971c36b289f301be9f095644b905533cb3626;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22ec5941a7f9b5edda601fc6b605aa9e9bc3acbda7d8cce94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6076b4bf7dca63a929141b83da0132ce02c3ce7dff55a320e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h158333fbfd28e89779194d45d712046e9f27400e081d043bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h403ab94f050a69cdf187534398b0f94698d3d8742bead3f74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65c2885e31b03626b58faa877cb7d917232adf1a754708c13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h606b1ab91fe46562c4a2ee036d2bc25b4b08d8be49eed1137;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd10ba1ab9130cab5e1c2a360c455529f8582d5a784b6c857e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h157880a14a0f5a284f1468ce23383cb8cb61b935b7759db15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6fc66b3b50aa95ad0ce611337650f660e2c832094a93bfc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had0140845452cbdd6e19ac818654491d822d04864b72aa4cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hceccec8953ef16da708c8f86b49c64e5e4099c3a54178479c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d3c20cedc663f1030222157bb4c4c7f0703aebd6497e39c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ed5e13f5efcb6a6a25d29853f850c0579e1b8030e838946e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8af06733565809e1546dd65b9f31d3db81f0fba8cc5d4628f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd76b2eeb083b32474025801b4dd3082f1c65d02931be56f41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27d74360219607d2414ca72aeb2c9fb2cf0c2d941de08e821;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2e9eaabcbd8e223a8772382b361ce177a2958aa10816aa76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48f993b12ab67b4aeb560f032bdae702422e3003a542f43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1d94df647edc8e673dcd797b9f90cf6cc8f6949768775a39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9de12fb22cbb928c3f85532c8c36e0de5c3759a79363305a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he094fb65d1e1c61c8edd6b34f696400e1a9901d480ea03141;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h233cf5bfbe2c26810124f1ec2d745b2ad177ab52e81c9e20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24b4237a841117b7ea34859ea709301e934c41438a69fde4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb333259a6ae5d263241940e7637111b913a9986433df01060;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf70a527edf4dc946310600aa6e49e6fa66c9fa81bb2de437d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8851b4aa9eee13ae8a57f1754c4ba4213493b887562ca4663;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf7d76a51dfd9552bed85566b953b2643ffafc21419de0cc9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0d9336888866285998fc2eedae5a368d9dcfe02272a2333e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h690ebde8447e810ac07f819477e448c09b172d4277a515d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbaa3d8e873bf41ec4c6319e68cadc7351b6da5b70159edb0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9c15bf0fef418abe1120b274863fc10a7807b41a57bd74e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b3059eeb89834c07591c67137d65f59864680a7d0afee113;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56744bfe30f3813aadcf7c9bbd7c825b2c800ede05b173d02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e3db7c0aea681ea05ebd416cd383fbcd14aaaccd674f85bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89a03af9530ee563dd9b49df9c51b1f8a2e2ddc6b58203c8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32cb3a9d2d65df579c965722e8b770f01524b467ff35af1a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c5322107821fcc3c6454429fa5cdd594e36d9948509ec217;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b89582c9a828a3db622f3d75ae92eaefbab2d09c95da5b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1e5cef01cdbcbacc3ee26a4a4b479f7b7a3a8dc5ce047a9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cb893971b381fc7520b56c92bf5de8ad3620383e878365bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb8a4a8a8b401b202bf68beed892ee3daa0bd0512978b1c94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bbc070c2a1cf731fb0838d4d2fdb57907a7110ae15cc434f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb235727b64238b368221a4a5e778493d8f31927ed115f3151;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d1ecd03c3b30728fb36a62ddca60fd6d205a4a7a1a9cfa09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5686e5f9ad6cb1f88f8be0b8b79d01f45152599b39a38782;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7798a61cb40748ae28d581e2f2d8684cbffc6c7f37009858;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda4d256905e2f11e43c4ce9a8699dde04586f2eca3ec74304;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e83994327b1c9745113974f9b67970a2d0a68762e240637b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda94db3e6ab935cfb80d25b27be3786cf8b4373d9f01f10b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h252a73a8027f3d2f7cb11ff90e9539a0a6bd6573eefb4c0df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65240955e5b899fb34050348d0d2db347bffa37f0f225b9d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42ea61b32e41985e4f974c2c9ec5fae909ec057a4b224799d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5242be03c71db66ff5b0dadbc7913276012a395157bfc529;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84acf94507325f148b06613d4572091745f21b11aaaaa3c70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecc02264127908338583cda38425f30d6a32acf54ed2579fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd945be1003f20f1f8ae74c91b760b9f56bf9d35d33151ecf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f8456c8e3539d275c1c9e1a6b384cf4fbb36ce523f5f2398;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eabf24db64dc63274a1eeb3df7d4c868c683c029294ddeed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70e5573aabba4538f680fa57eddf439259b7e4247552051f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h856d538862d2f7893ac13a4ccad5dc389721f0e17c20e7121;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30dd7f5a0ff902e7f0fa6c0580a9eeeef5863835b3ff8c9b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he09a52a3bbf9a947309edfb41f3b7571b4f4a3732b26baed1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a8eeaa4c0459d333b6d62c1b8652520ee435694a4b078fdb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h303e7e79d4fbad9dbd9cfe4bcdc080e11b87134b925d0de72;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbc3bb0e010e0c614d7474d76ba8a0446044508c3aba0d111;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bd8df086c5cfee9f6430270fb7069ce7e3bb92681b64a90d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4ab6a4035e662e7cd5d5806509c8df0eb0f370656ae4492;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1762f1147eb4f63159c488712623c61aeec5d6f7f4ae9474d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87680e4e9423b682ab3b0b731379949df7245d8f4afaab23d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdcafe6bd8ecc3ef483bc5edbc6ef2414f17bc3cadb82af6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84da646ec040f000d8d8e74acca2516dfc55e4df539f33569;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h537682ab40cb5716e947000b793f5e300d89ed7327564e7ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefd1e817ca459fa77482767c3a665b7760668c921cd721c8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h283fb80f2f195fcdbb49435045e65aa211bf232ad3e937e70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fa2688e5103a9df9aabf0e7d6c0c20e746807f7d1106f99c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb26f274b6fccd6d4bb935cbc3161799a3f0f1bf73c895195c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e652883619fa0bf132c07749253e051d84d2f37d8bc1a859;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d86fd541422e6737b7d0d1eb525e72bc863e27bfbc70dfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65a1a8d4a359a365bfaf867a70eb4c9ce4ec8db5eee0ba1f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0e6ea0f7e1793e4399d1f2a75365089942676b0d1d71d8b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9813b001015f3ac45635705d585f92e9817814c50dd315834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3dda01df90de906837dd58f8b7aec8de81ca1b6453fdb9c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb078d9da0ddfffb04233cb982a4a5e0c0400ea225e640036;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57f4955fe9752ac64e6f8395f1795b3bb623a107564c29563;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha475e74a8e991853ed7b31f7bdaa327fab8df7998b020f4b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18dc72a355a92a54936361dd4b7f5866fde0bd6b22cb22c0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96abc4f82dc4f0bfc5481a7b95fadc622fe213bf948d5e23e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h464b3f898a40bea10a5ca6f28fb2e75d50fe66d8a55183ffc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb8db9340791c224a4c1d406aba4fb1c4d15a004755c671d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d2cbc97c8aa117962c70ebea36680184b2b51ee3cf5f59a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e503e6089feb95113871fbdfd1f9db4ba76ecee7145a55a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h575ea1ca6ad52b8b3f73800369f625076bd548fb8f30a75d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76de8eb70a005eedff6a4a3fd96b27066f52599995a77790b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd269e59790a12d07fdd72053bde8d82fb379c9085d1b3e28f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93ab7e5b27891355045eab25d254cad520a8cf2c18df9d574;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h802309f579b3e32e567946cda22f29eeff08b2fc63e4e9fb4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5470f756c77516d4444cd300acbc9f0cee71ad15c0dc4e41b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6deda17837c2df84ca1bb3394e63ba318f0777bb6802c3f96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec6ff8487dc5d5efd87d13a367e9b26febeb4a291059ed1b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa399e2c00c1896b6f404c12441a91e5b0bb83350518505ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he92d9cf162b91263c696b9699b3d3fc9cd977ba98126324f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0caf67506a3657056805f5880428261493d9cd6c414f857b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b55ec49839b694d510df1306946031f120fcac12dc9dbf64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29c5dc4464ebbd555d57e60cae6d66b395aed68a7a882b618;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a21c6628567455bef9e14ebe46ccb2c7590893643f6cfd37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h878f770b850e48daebc533372be0317a9319cd80bee2bad9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h295aad58a54324e4cc6347e9245f8151f990ada2af4529dfe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f7adbb9798150b038e73ab0a02b6710a7f093347b22c41be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf638d0997f072363573c0f911fe34b54a3667be0a639c358;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0bcffe4883271b6ba2c83453554204a814107df33155280e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5b14e4d9829e7573ba340e71bf79e16e501f1323a721c4f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfb7b4d1d0f90bfbfa53be5ce9b390d759a015a35ed313c91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d1c66ab4b84f0fedb73f0678bf12d28d4f38fc7d26fd444;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5c22c78a0f6be1147ba7f849d2c637337bc8a2e09c81b23c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d62b5c752faa01dafd2147629eb45192e901aa2c666b9ea9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20a59b6eaa6da6d4261f68993e7fdf0d9682f3ff6fc678be0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75189a700b7675fbf904abc754a8745e3b6e1ab6e45082f37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75582c6251e68da4e6ca169f75ac2d00502e8b4636e3a9a36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h700d6885f98d500da7135db75e8531f569e3ca22a934a9ca4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3215a651e52a3584ec3ac3557e8cd05d482f9b63ee8f57529;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h421357235768a98764972ea9010b0d3f266a86a856af5d1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd2d60aa2e82853b76a467a9595349a188e4a241543b9b549;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19743350580f4e8c030899f2b38e7702a6ca9377ac959a771;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h268a6ab39e2d977727722c82359001d28971a463e2c6cae39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22aa09279f24d0ce74b31ecff12291cb15c436d554bde104c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a9cddd0c398be58fcc95615233f9cc2a5682a929b9667083;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h911b5fd5f2dde9d3beb597ef12f16a6f987e8b25708ec41d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h654821e9fb0bca5b4a561fae2c6fa61f071f1b8a852c173ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b856064f3dcbc0ef84c022f0d2d74aeb2fb8b1320a1c8074;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4df5f1e06b179b0041a2443b4d996f3273770270de337ff1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc35bc4c344b9d97c44de8bf192ca20cfba6c50ff2d8b5c08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf919397b977f01feee0065d7b64b59708455078b0cf044fe8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee23a6fdd8c777b3094da207b13178fd46aa642a77af357d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc674fb264ebdd1520813c55ffa5111250fb20067e2bc5362;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ef88fb5c6c1fab0118c120aa29bf2bcb881ed5598f1e7023;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33ebcdbb49274112094a36eb114b3c49e845202e06dbfd490;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5209d611ff751f698a1c981bfbdc8d7dfd6e32dffe929019;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5c259f9639392e5b58f61f03781d1267d62429c5386334ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c019623f4d0a9a021dd6d7e6a5e52f69f197c5557fea2d09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17d57bcf9fbcfd8fe57a4eb8ecc3a6ff457edf426bcd49e8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e7399346a38d2c17774f0dc0e6dc94a597dc7314bd31b193;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h920b56454038b533bac16177a6c09196e95e24f98e36695f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f4141607ee41984bdaff9e2c5b5540951bb748561c24d94f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab9803b0f3f54966cef2353b227c1a77f3b7c6cea63d854c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36486aef4cd28f4d6522997c18ab572fa508e362b64dc4d6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h794b48e0184dfc0d1f7cabe90fbfca7cb016e34a17f747d1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee9b33af66afb06ab45d8b67db0dd0aa76177d86dc1d97325;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24fd858102a993186178eee9cb5f7bfcb46c41300503be6be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3643f635078b237f91416738bd94b9995d1f274d5e723fdaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b3e0b55f3ec93ef119d24a353620e8cfe1ed19cdf773b89b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c8a100db93bf8eb77f1c433cf9901b798601254e2e12e53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e6bec1e2d1b8c61092255c2ac42808db73a3347f9829180;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfea18c24d9dac7292b25f14932107dba67e8adcee08034144;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35a485d7470af649d39100663ed2f0f96819e8d67977bda0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36d490273a4e95c4610346df078bfe7a094c07c511dba6324;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e6f3d98e7b4065a05a73e5658ae3b240e8c564e19640da63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e635be86bd64b33eb3a9a4cb332ab1be0eb6022732c4dd3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3db5b3f2011971a8ff99aec37f9cc56f2b2995be1325254e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf51801e9a99550e3932ef1b01a3752c4a1a7049ad153401d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf34df7b8165d281593d5989dd9deb19b08d2caf1df3d166ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25c89e0536605c98f8f17dc3215e50d28144a66ef44f2951b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde9b52e9a0cf25980f88ae98dafef89475f0320472043f4a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ff128bea1aa14b1ba1717f052461c02df8b42cc78103dfa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h105998124ac7ba703694bc2386885a85256ab465374ba664c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8eae3cd92b027d1fccbebf07d6a7e21c6041e15aa3fce763f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d88e52fa47479df43c46ee06c87fa202a416c89d24d59b55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38081d97f1a882b13fe1d0f5ca0ea8da9be3badfb55de494f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77bd4c4c8c13a3916aba7aa908c4cf8c3357abc0549381aaa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2c331154b3e3c5454f3c5574e3f203bdcb792339b891cf81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46f8f4cb4a467597132ab14906838388327b9421135a794ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb522f081c3a540d6b1946cb69d63a72761341e7afd387a02f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb278c81bcbc137fc2941cf670d544cc4a169f1aac7e1fbfda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68505bf45804cd1215e9fa055f075f6b1a5c0ead8955c5289;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37583a477459430c3d3e57fae6afb76b92e852be84cb0aba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92f18f19e7d60c420e58edc3508f8e2701d846979145baae6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca7d450371794542100bcd00e1a1b4b52d42aa32f73712aff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h545ab8c8917af7911ceddeda4b1539259b470295cdfca20d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0f06df3ef532a6c1448786ffcab42287e6b888c5ec8d8083;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40b68c89297af7be1739fc9bda0d5cb0fee342180e9b91da1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19dbb33a228a88f0bf6f0231fd2c003b93be72541f0813b26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9cbace6a72b6b60023afc58a2e689bcf9bbd3e4ac823b7d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c39e4ccc9e2a39fc5f0b1b425cd99e2f5ed85b75c57199ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a0b3015e2b8a8be39940f080f633fc2c0293707f96986b72;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8da5b00462692c243ebefa16b483e84422f557b86100d8b14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ed33567243002b17d1f2f3e150f5abe4724462d472a1816d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a85a26a6fb61f68ec56677390e941ba3819616ab16a5359e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4d1db2878956b19ef5c3006f92c33809fd3e843b759b7c50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff22a5ef4903aaa84c242234fef88a3228242de04e2ff6d4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd09e8a81892d0fba84fda45fb447d070713a14566f7b2f527;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1973cdf1e2d11bbbc8897fc9a7097659bf40c970fa72feac0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60b8e3783851cfe85a21bc79ca940bc05fa98622d64107a36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h275c217c5733ccca081e83324b1b7d1103637692df191be55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90329779e4433f712cf82ac3f61d5fa39d2d3188502ccf3ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h258d080b700b6d490dd4150b1fc39909df776764b8039da62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h248fc0c5b9f3bf4b1782022270af7689e0b17bae9e73dcb85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h323502c35928a8b66f3cd0da7407fd64b39c3ba090516f904;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60567f42e5b387c92f8f751aab787b92b8dfbc3212ee4410;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5caedf2a0826a4f3432cebbc2e1a98f2f7f3d3cfe4f0951b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5648874b008322539d2d1e2057989816c87af1e910afe6c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf57616eacd7f2e756855e724fa79fcc054f845f5b2eb2141c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb40761a43ae6d37b34d1908839bcc816ef2757a56061b421d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb686faaffc171f1a93cfa40d336127e3f4e1b64532e41a6b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h175b94a159a5ee653f5e36560d5d2d73b73f8e637e39d8e1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d456c094a4a8aab94be3dbae6325cb4844811eb2339dcf82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bd74a45f177f6bbcee0f78a2b6261485f93ae8fd0e11cc42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3acde585d7ec157435607f73970a662213717bcb16393871;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf9b0fa41210a9ea57f1f874aad1ca31af6e0db60e3702a49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5861cc78c1365048b360d607550cc79533ee349e120efe68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha42ad550f15d1dd31fa775e0e125787eda41e97cc244d5e80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20485e0e13b85fbdbb4f04d27098292701e0e27495d93907e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4cb1245cc4c223859ad4b04555fc861dcac2b9170a1e348f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d5da5b0191fcaee0fc64a4919008488a6cc256c9c01f3c83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5f5fcff4742200dcff8cf3e53a2abab2f4d838761c89ad5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb38e1d6de5d064e4f42db33463665481d7d2b67ce90ccfcdd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h159eaa9ca2e9a4b0ba10980c92c6265a21f49c785310e8d3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62747e0bc5fcc98474099f30bf68e38efaf5bb644d3ffac42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29eb47c5dad962e16fc05b4a6dcde736a690a307c1e8ff965;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafd191e48cf89bb44cd76a99d754010ac5d4209e51b5d70ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87cd8d2101b6bae6c9a955c3de83d246e8051c33ad8cc5e2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h620311100d9972837fb66ccf0e5770d0f995b8c30595fdd30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c0b8909bf6eeb8deedc0d915f04099c817e961bd12525ad0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1177c861e24e253f2d1f4961757f29f435fd63cd493925b41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1532a87dc652d1ec3c37c507a0d99141c1b25e42bef2f552b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cf122b01f5f3889cd66b024bcaede2a582420bf6734aaab8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f4f977b6c569c8aad1af2d8dbe143c9245df9d175558e2e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74eeec923b05007105e176955214ae8d9dbd743e245e64ca5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82ac559360a02cf6d671e715151d054c594e9e5bb6937ddc0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24d4009007a622cf889ace0e1fbf44b88ce2f8ee34b4f90d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8412321fcd5bf1c1c34e68561f650b0b52e361f7133d94c1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9e72c1daae50daff8925aa6c68436bc6b63ff512669757b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bdfb2dd92231baecfe0534947625e360c26b2b7f9cc3f786;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he58a873c4169ec9f8649d63b657eb776a9b455359e6595add;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f3fe518b6b965b8d3b3f6490dfecc9e252571f113093af65;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafabb3827bdc78f24391a0f7893f62d357d5f1c9a25ca1a97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc16ea1f0698e2b9fa6b246ad04c08cc505418c5a6e6f909c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2945ea25b85f5ce85e1c67721815b0794b94544122e82b616;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca318603b020cb79ff593af9feab11e902bc5a7ed58811f61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafc1d3cc92013f8b6384d1f1237fe61b28fd621dc424eab1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a194f568d8fd38b31ff4ca68ffda0a2ec5dabe9178012f23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d77b23a5593971ded9e2d70365fdd61219dce6fc5e0e4626;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h516fedf4724b755c4bcc62b30093331d072b0be9b82af71fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42bc35fde0710357da3ee0fac09b9bb6c6ec0071bfa747c32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he034514a6d9187a79f1957d39659a02a7b37b1969de5e838d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba5678f8458a6b651853ef4ecc2b3d7d5e5dfbabb44cefbde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h449218fd740ad041bc8a0c701c669fdaab260e749b82ea874;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c527ba6d89afd060a3b2004cf15c6b3fc24e7a44628708f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cc550ce7e1096bb7f19a7959cab0fa04617c9090b349696b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdee7af4421506399650f15fcd155f3441b05930aa5810de1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b84224d5d67621cce179c8ef4651e75c404a86db09c85c33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1e964972933ab1cf317c40e590091228409ee2359d7ae8e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f23887d9216a3b4c49530caa458d06da03e8efd3e693912f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd76f4e40ecc3593204f5bb9b752560b51a55cf19123be3c22;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdee19fe7c134c616e6d80e63aa70509c21cf93aaba7e7cf5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h200d8c0cb1ddca5e44660e0b0485a990bf9c7689e9dba2a78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he50cd1de161d2560af9148d1f3d9612337e0470b2f2799319;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc52444187fe0931ee4b8f90749567dd76595ffd5fe64cd8ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h457743c9f39724033e42d13a7f2bb1b1562705ed770873736;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46f1deab0c2b4543732850ee29f90237784dca6b71e701344;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63e005e61acfe68309dc6a07dc59a926bc8ded515cc2d6dd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had9a8aa4df0c555e34f790b4a1ec30c08ea1b968eb64970df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a5558c730e79468ffa432d15c72445ae831a6e8c7a2f04c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3143cf3472d5523117a4af1c4d05e890ed31a16e83e27a71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h804ff3b62de59131613e93df0109e008dd467182f6cbfa55f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccacacc98a6aee4befde716c396ba538ef1d245c8b0b064de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6ded9b808e36f28c5f6c4ee83330edebccafc84da1e5b041;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67aebb76870780c9d7c4fa74654adced89f4d3e160b48d37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha178887ac5354acdcf8908c04304113c72abbaae205208d18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h234176551112bdf77c662a5a97829b5bd9b22e458703b55bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4c10b43481352d9857501703eaeceb381a3e4fbd85fe7fa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20df87761505f77f9a3508c2ecdf9fe3e8213d3e93d9109ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7564cbde34d4b2b477bb9d9c11f7a8b45dce3004a694f551c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h867c3c21b23bdb03df6decb7c2b6e5ad99f44ce0cda55b808;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40eadf6bd81752a17244dd20daf9cd4391e6dd017213fc50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf85999d6add7bdbe4092902e128c5b5d800fb3cd6f26b90f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heafbcf7825da206f15a859f52a373ee9c2831c16f76ac7238;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d7d4ebb341bf0bd4e4dca34284e0c25313c7d7f7c6a7f5e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1c2e73ab97654bec5df3e4f1223256c5adbbf72049a524a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc5f1d45001fd199aa161ed6e1833c7b9bdb4284d9357888f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37f9bb98e7dcb8e8b4b83f0864060915241b18eb65c44c15a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h542c239021ec8371a2606bc02213ab945fb967a8740b94e71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f2cea2ddc74b6ff934d7106f938ac1afaa87e77f3ca9060f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc67c281149ee023f8ebe931e78be83afa5080482eaa0f140b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ac1fed39960ef0a8af75e38627b3806e2e852f9500837a1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fcb368b0ade947f43d220a4aad19c4f9268b82a375b7b3de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde781c0e1a5b23698dfb9219da349f00ba652325c5fd68f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c300e4f73e3a852e91ae88b6142abf987dad962b1d085edc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95d1f85e263071e5649b7519fbcf2c1814a590139ae1cbcef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74ba6f4d17a42e39e41b170311ff6ad4827bf844bb10e6b4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f6d81f468a7ad9a812825146ce95991c661482f20655a625;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0caa1aa0d86027b48a0512b027a40cdb0d9e3cbafdf27933;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1656047248c207b123e29ed311763cd4be50b3a66a977756;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9162d311e560d4365098f13d06e12dd7788e4c232ed3d004;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90658e8482d538536c79efa0bd4a34576468308776c626037;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2814c9100530da60694cccb41e38c0353f18b51e4048313e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf66c70a153b259f2083eeef7c31d72175c47595d4f45b53b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc04af880d2ea1d94d33b56a2d6d50c0ed30043fd81bc7ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90bd5c77164ec7883155905d2062499950ec07aec5ce809d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5c91a3085749c864437dc559585187acd2b6bbcbacd0e95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc9d596fdb5118c566e0600809d9df835ddee0badcc74d4ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cf2f540261be491c5f3e58c30e9c6582ffd89ff3dad1197c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52f46dfc6d5bb2a47a78c589c5accb67b13f5fcc9fa25b2e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd37d7af896e5aa6d3184085e6bf49d420d65990f24fb7e5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ffb5f2ea5a559c1f749a69ac905fa28b62a1b7af4f652edf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35685eea19eed274c8306f0dda903b9702d3bae037de655c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19e4e8b2cd0ca6143e7ea1bc0e83a1e0e702ef46953dde3e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he45837548e185ed06163e1830f7d7a095717f277e82abb802;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc46446d593081f72d5abb9c0e5e584fc380a2e0e97fe38d18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10656b1e897e1becba1698f4ddb9d029c8c828eb6150d3ffa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5158f4ab089b1cf34f50e49d876a9a88df7da4429f2a87a91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8a7aca9f8be59ec7e1851f989507020602d16c53bbd5f7cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he234e7e24ea199520ffd930ff2b39ca1e3feabee095182dba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3779ad52512705b7d1b80ca74bff6538f5c826027cedc891;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41afc37b785056f88bf9b3daf46fb8a0f160b97e1f3464d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5e09a7cfcec07068c6d906d078fd28b21e9fdbf113ac404b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b2ae707496d42d8278139efa8f86ac11441282a36dcc762e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb133d9345df60609a5245679cdacaea7b0a3becc5b8801b15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ec8934a5529e60bf7830730e309b9ea7a7cd9f1b0f43c0ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h145138bb64e97c8e7f6ffb7d1742eb66a0c22065eecde7df2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2955bee816e87721ce1067ac4141a7adab5e27428ce81158f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h383a8ac551c57116c6c64185be81c17760252bad7bdafa87a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89ae615e72269bccfd47877b65c1f08bf9e4a38b3d111bc78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13a4aa9338381d90ba748b5cf159bf987d08780ff40a548dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2c11bd20b9d91bc9ea203bb538a4fcd4a36c162acbb90970;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42fab1c363bd379e68cbaf520c99e641fd557590c5ed23b82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he214f0f3bc0abadaff3e726bc297a4d09e2b2adf0fb0e2445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4ad797c7109c33965a1cbf366d3d38d0a931a1ca3d9e24c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf175dbb90bb72c7a1765400d172571b638463f7fdef50da6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38498374632c65df60d9c26a60bcd4124c9b6788ce7a75dfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b915396cfbefd68d78fbeb4528a71162e39ed7fcdde6473f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4679ae857a2f9f6ee27bfbae03cc71a8aafd34750f8e289d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h147f496f574add05f24ce244f332d251913ff97b59794e69d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8e130cc38e26110ac52c13cf412ce6e438462f4806dcd47e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h379888297bf96904479614cf739259e34526efb5d2d4d4897;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1acafd80961cd022b2a44a8d469f86de1c5aee5acad4481f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bf5a9b4f590d85e72872dc3c7513b68cf2c795725e94dcf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefd3341ce1bdfee706cf59e86ae1b4119db31b3278d587e4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb37ab88f5eda6ddcd7aa746bf5752f7febb4fc365f6ad9c21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d8d341dd06dbe81a9d5779e94eaf31ac597cbd9cc8671e11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e71ea5cfb579f2c950d4abff18e2c5935df3ddff99cc889e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3056b01ed8c4951c326682579537204cec970fdc351f7280;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a8f24ffae23acb65254091e8933868171cd13da13b12038b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4ec304ef4dbd596110e11e4f7a493f919e33550ca4a93276;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b27776a253fb1fdaf9dbe3482a152a3efe8ee1fe7d032c2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab8ee2ec7993402b92e3cdf9d45aa6709224cee26ca48ffdc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fede04b2ad87938ca5ed3cbcd8712f70433dba91989a3553;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7eb8335525b8ef24ca3e7d50ccbd7321465928b5afe58dd9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b12c5bede2dbca70c2322af91d877834d5ef1dc0ce315ee5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb986a25f5bc1e03e2f573c86d80980d577aae215d82bc7f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7077783102bd72cd5f5e2fc3e8f048033fd5f2608db0f4d79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ab94c0d8d80eb21772162dbed6c6d62fc1e147c105ecd948;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha105f6f13835656c3b89cf1592d8c4608322936ecf17e1f79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b62479a6eca54206e4f60c5df826432ab3561cc952e32119;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95cd502dd3220dba75ef68bed93d82ac14d75b3856e58879f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf374d33b0dcc8a1b4df3fa8bf426a1445f5dabae8c8bfa6db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h309ab68bc3930cf6bb46984919739f2fca96edc92478cc081;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48a7f064063de92d8e16a855e965f433fdc849cdc5fc72e4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5d14b324150d37b2ba61582300b587469e1850c7ace21061;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b7cf5894c33068d31b990796e34f6b56e21778f11ef4aad8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbbf644d2a2a2358dd95913c08f186b5aef37a56d68258fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61d6797c99ae5d4330c31106470f189dc85d172e249344d00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h718a78fafeb9d80bdaa159022a33a1d891a3be419d6074c24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94e98ab1c79418999f54c4e1a059c53d7fbbf24c469542e29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8658eae8cc2b9b027608b6608ff9bc88ed763899c29fec1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed4b14b6209ae55391c050cfcc04d67235cf2715d339aecad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48bea22a16218f54a23c4284f478f1c30b8e19b9fd41717a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41d8c6d0f39e4d12caeabd4f224bd780bf80b44ef9e49a6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e28434865e25255e13681f09086a3491af7b8ab95bd76f8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h708ce74f231a0eab9745f6193238f20e0cba3ffaed6e3acf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b5778b57cfbe17cdfee8552ef5e49afe952e4141e5e306fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf954434e9361def3a0d8081b3df32270d0cd1da42ef082e75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b7fc44a42f9d267b0274df09ca0780cd5dd6844b9f447858;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90c8db3b384a146e3be08c7af51964995239bbcd2188dbd53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13e9bde95936d66fd7080eb105438c80924c92a4dd54ba4e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d42aa354d9c5f02f97f830a73f565d33d0f5331c041d6bd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2e236962b60065ebd5b2bd3d274cb6651d7816d506d9b644;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab1811586f71ef22fff43d8c032afd88bdd2b2b31ddae40d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h156673e672bd3987e6b2c02c254ad85a4f9c464dd42127a3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ebbe82da0498f8c58a1c6cc12ed993c2c54886455576e105;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76deafd5b331af38b73899ccb132c5336b2267c6c8c173362;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b66a9c22fc0322f6a7241de5f51024efe6d9abe3fef3e98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h336f49faf2bdd4ad3b8be57d6b8a815a642cdb3a4a1072d10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcf5de35bd995b830ab5384d3bf77389f64298790520f4883;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4a935a98865f522e49f07f081db1573374884d239d411ff7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5674715ab17075a0d0eef402229c1ca0fce04d5ce0d227920;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc18c55417eee8924eb76c4473524b134a5c511c825b4a82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5306ac6ed4349c0d0866b358f7911a3cb7ef4cefb021eb549;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he93a68e351323b76bc606eac4592c224f056b9247f29c327a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h723c344cb5364f85d56b2eb777ebd21a1be1f85bb33fbefd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55083a58aa385a0f38bcc3229a6fde6a9f4937cbbe33af86a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21d99d7c05aa2ae35e97268a2d5d6ed175b8720454052dc86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2ca7bb3eaa94d5d9eb65c5b485a9cb97286de0e51be0a006;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4724ad093cf3083b0a4d814b64cdf453a23e742e0042d16a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h685069c8355b781d13e9a8f45a5b18cd9e106ea8093064653;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf65088ca2cd3027b9ea8db47159a9f3984a6e075bb37f326a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cf1242aa982a4213edcf375fad63cce847e0748ed682c0dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f9cc2226e5774eb1186063aae0aa15521c1b8e3dbde486af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8d64ce4b8ddc5537586384b005fb632b44d77e69148e3b25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87925fbff72c75535e1da3e5e7ae146ac525262eab65cd6be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eeda19511abd3c6da4e7576fe9bc3921506de2d8dec89bd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9284b638948f7af2843c44e520dc90caa907b33b2cf2f4de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he33621cc8d837ac6a47ba0d083f7e185fe2dcaa640f7fe0b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he878cd93fe864ffef796c09c3ef9d15e7f5ac987112bc6ce0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c8da6cf91788ad969ea7642a019a9b355bc070f6431c89a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1ac46966cc66c95aacb19cb59a2c5de0c3066bc5fd20beb2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ca9f1eb2abef5800e8f2b6ed9c6a155be9677ec5d7b3ea4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h311d8143d2820709499ff8ba68b1cfb3f6b754423e89226e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3f6873a127003d4d46942d409e78b5520c4f6ac7130066cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha204751c9d082a998d14292211281f1f458c641d4fef430ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h796f911612aee4c8c26ff2e2bccc725bffa91fbd962db83d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d734490f941847fa4441fc940cd45e3dadf79dcfa1052951;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h588d07ddd61257eeae819d094322e80c3d9faf561827288;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h803e39b994811629a342cd619a3b4f91119ada1378c9f95d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb3691b6c2e7de96d1bf5ac8fb265da73c70f87f49da8d60f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8001c6d7d61319cfcf1cfad409a0394e0eb98b1a13a4a6bf2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e7ea00725bbd69a994b34e3f7251e29fed362d6e6c597ef4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5276b9c841eda02291543995bd0349ca64c4be0a3662d4ccd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda30a5125e4c3845498c05f71a6b40b2546bb1f9bab048552;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b75f1c8c1158d14c3c5ad0f8adc668803755c72f8773af7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf73746cde6947495867f06f5b7cda49d587c84d607708b69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd712fcceea7cc4649a24dce9d2894301766bd0d0cd992a2c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31ea389c34e45d10c651162b6cbdf2fee256e0de46d7f42d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c6a34d7ace420e8f8fdf339ea6312310c1a6b46e70819283;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eccebe47ae4e4c11096073ca2366be763ff1db8d12c0081b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b8d7d356fb5043fe61ea576499c15f684f9082cde27cd7b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbb47ca1f7944a96a581e2681c1143f599dc9da78c2405b37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d11a39d73c43bd2d5d23aeb2f7bd4c046dad8b3cd4fa7eb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h832810af884d19960e76e05d6dc616691065304799fa30565;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d9792cb954195a4324aa33fafdecdcce570da0de9aff4236;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a0bbbb6269b9ac3662fcc7a25b19dfac3864d2c777015db0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf90133cbe7b584be07a528bea1bc8bcdce5ca03a09e6b4ef5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91c006b57e72f511a54fcd49f280db1691a4f93964af0e751;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a2fc12b780f34f7ff731089e94101f55709d485f1567de50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb8ce7e960c34d3e5932b34df624d98e310a50d8311c3a8a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4e1cec74d1c448ecd7c479ef6d191502d40b8984ec7c506a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf33606382c477dd28edfba2fd77b8e3c3bc398fd24bc2f2c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd40cbb6918fadc169a3f1630daf2d337f8ee36231d7e150b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h417379d037920f82e1545514b7ff4367a7db01a9e76b2e033;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d7e479b75ac0b32df2cb705f5c0583a11c738c8b2e5ba0ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf702d5c605eea67b5162182839451f7337060a25bb58651e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86b22c5c97d134bb9a9c52100024cf67286757f219f374241;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16692d920316de9e3cf3708a57ce148cd20fe5a23a04adbf2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72bd3953cabbf784e64a60cf6273b76ed07122d97817d72e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb757831883990c0ca83a66c9ab8cd51d41d419008a610607;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd22bfedcc4e1cf80e197649fbe4c23ad197ea03a8c1572ad0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h811d3ed785f102eee20b96eb6f223f9ad58bdf298c030d129;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h140594d0f9aa64fafdb8a2e7e6503648e450c858b25e9d289;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h278e4d0d93ede77ce523b6c0d89fb94c8a5728c8de7fd55d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h694c933ee943ad88614680b9d9c8f414cb9b1f9103dc9cb9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h136cc610f9e8220c21c5c5b2d3ab988ccfc4a916365587fbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8952a3e44ca081d35ebf0fb5107dfd163dbefa6c9d65533d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6f0543bb6ad3d664fe3b7b0b197d3bd688a23de65381144c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4340140f2d00298c07bbe349e0f7561f0278eec3f5e866809;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3bb1a2a4db9f5aba996a166e40644c461fdd178a5835c3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52f353e1627e806040e0f6e41cdedcbfdc8f8a0e4a7d2e3a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h144c1ac3e6f9fd795978b1cbf7974eea2b4ea0b98b00b3a66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3475793716dcdf8c5711dd71f54e411d5a56aed0fe7f7de3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h196dd0c2e7098a7fc423422c5f9db1430a09395bc2c5f9e06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h931fd963e6bcd48538be7cb09c192ccde0e106c930eae2145;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h359751205e5012be7e148244551c0ca6ccaca8e26fcf31599;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6975012c3e07546c474d5b309fcc9b046edb2c412b6797f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74864b62408d70ef007464344ad0907de70f5d0a99bb18f78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7902e8f651185edd483b250e628b773539f103cd9f612272;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heda70408862eab9fd409424776a76226ff368397e9ddbc6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8cd6ccc489648adc7e122215ffe0c9d57b63e6e490518926;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb30288deb9cf61141f12e0be9d95ff2701d28dc70877adc41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd66599444b788f9797d1190e0e2bff89c02998514c05320be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ea485655e54e1525e216b32d07bdedf5ba34dd02696cd55b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b9e1a3d60cb94f17453156325a0c4fc5ebf90551216d208d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e72729bad5a2d9c3597180ecd5e3d2d0ec2d527c0c15c189;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc63195660447279b134a9d7bfcc5012e64644e5ec3dd1dff4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc98dee44b43023e49026fc14e2868edd6fbe7ff2172c32b0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6484a4b6190623101b86a2782bb495b24a9caaec4e220d5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d98ee003bc8af37b746a066fbf20a8b2a75a71b9ec59db20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3dfcb09dfc85e50a1a955e4cf8a7388bb018816a9bc7230d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6fe0679c7288d599f6a3b362bdac5cc245944c113be6b29d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2da31adbe692ddc0da1745bcc045f62a4ee45365caa32a5a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1624f46605e247ceb182fc0973fdc326f30aec32a90013df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe29215f2a898800a4073b79c65c60cc93222f0be5b60d2af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8443e3624cf2be837a700da00f5a9137b4f6553cc1885deca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f1234cbf9d364da518399757e8f6d3a0a1ad87df2c84849;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b0fe8b5d8a237f0800875f796c1b29f9efef0db591b8f6bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb423d4294d6eb470a7753a6add7e109e8c92b898ae23f468a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c53b394adad6bdd7a89cd6a2d5813a7b052731e2e8ac039e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6d48f6f8fc3da240ab653afbe092595bd4cf84562edcfea9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had595ad8536cb8e11d064a6fff1c034e9ce4dbeb39ae0038f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h513868000ebe4f532e1f483c10287cd88094f03f224f54bc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57d90613aba7fa57baab4693a09954bf0352fcf3ba8afcdc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae63983243094768d5757ccbea4ac56d811d62ca01405cfa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3205e79e98766702e6c53595815ac62a3f8b5bf6b691625fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68b190d63f3432c505d7141e40f2dfaf7be5abf90e0b186df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f9042a4e9cdb5d253803e3c6a381256cbb995b69bb064dee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h163a397e268c8bb93b509f5725d15641cd2aedc15012d89dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1ee27b64b3a336b5ebc0ae235172682df71436c1b3abebc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ad465893a2613b180bf5f9d8fcc350cc0f09deeb6408cd1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a68f7039c6937c059b00b8266bd1d7a2bc202b88de8267fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2005de349718a9578dd5ee58eda889cf0ce380c756261029;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha91c1b269cb9bcf77ae9392d2be3c81620b42e92e82f05353;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b093215eb5d28aa1f7144d5fbd0f89850f0038e8cf4333d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2dec29624ac5e1ab503658983e472278ff4b6e30b122857b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf68cc0d5e1a62db428f64f4203431d95e7c27aa7fa922605d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13656c20e204bb58f7e796a971df25172e37099c8b704a4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf67ffca9423b8f130d41fc84b2659efb4f8a7dfc85f6bd19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fc91c15c8361be4dc38e2c130162c33493b61738085a1b46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a4cf3496435d381b83ef6b2078474f62b94a0c7e535039bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17bae336630fa08a86cb3d7fbc9261fdfecede702e97ffdfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3598d32ce5e541640f472fc213924d4c17654093c454ef7e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bf1ef24af6758c645f65149b90232d2e8d4941dea37efebe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedbca00d63acc4294ca44648f2ccae077e819be6115af55a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6297d09703fd493d3dd2a012146ab4054f749a4db5a0706ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7191f060af03a045ef515a64fab8cea2a3349e899b63d6d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87953c57a184f43163c21c25e124ff68e629cc5c986a652f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfef6442340e28f8aa7c4f4b0e73387b998f59a0361b047834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he12e9f4e6534afade6768cc8eb868a8189fb19625e50c20a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f8ccd709522503c2a91bc8e9d0b463d3a4643dc0cbbaf2bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9f034e0a3b0cbaa866d55b67d7af953cc2d812a832cb2716;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12bc81f8008dcaa651e05f5962374a75494d7337e964b218a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc78e4d16491de6455285c9ea0e7929902f97868a4aac016bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6219f528c264753e9ed3a62e87f278c32465ad736a5753fa9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf64a2d1840c1f9bc7e56554877f5514fb59a71735fee746c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56e63fd8fc2497cc319a0b156c63802f8add87da1e066b69e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha28afd1d61d293ec16fe6ea8b2e61e91593db4a1004a9b3c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h297a648f42892abefec6e99b7860e263f384fd1b6e0888e30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd60b1df485cc1c61d70399c63a6e0c917b9b16624de75f92b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he548e71e652de158435f733fe4cdeac31cf9471437c290859;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64a03779467c8951d36985e47363d4fc2ca4d694f6162ec48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24490b2e2dc696bc660e0692e2c02919b14cdf3b9dffba723;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a0a4fd06edbeee5c212d8cf65e7d9309d7d37f03a253e423;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha04bb8f4cf5c180cf18a7a5278b6dd04eedd260dd2f7d15be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdf29c6ffa9a920d557add8deb2c63178bf70a4d23151e0c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h648383a10ee2cefb5ae1beec9ce4407c5cbd3ce53f1afe6b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc44af6f84646bf5c4b181292172bb4b0f256dbf8f10ed6e58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2eb9fca3e30ebbd061c368dd653fdba80a0cc6a956903f8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f6efd638cecf906f2745a0f0f94e16c729bc8ddd36211fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h855cb2156233995c83ec35a111872316d1cefd009a64181e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76b7edc7cf8b87dad5cb0d897cd334eb4d1d4b11e989660fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30aa3a55ad10afad68586f6ed3aceae06bf5058e0b7bae6e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc19c2659d8770a53897d0cca69772695219f4414a00a02f53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6400216ec9ce4b29584995be411b3b175881f5ca10fcd339;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1008eca620b1e7704659039210b0a8d561508f2f6e75ac905;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha47a3b8264eb9b2260d3b8c63d8ea66830ae9273864523e03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c2f7dda5d22f238b2f208731e1693562f62fd5b6500865af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a6b15e9ab1286bd71b592091478b4aab86fe7d6cc0c27cae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11ca355fe2aa9c7f90b20e4e6ade0107c3ebc9db2afda6ebd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4796f4ca9052f1b769277f39d8ee883ba183736bdf36205da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac3c377f092930ea2d5091788c52f07b5643d87ea2123bbe3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3bf19bb728071e3f28471ca1f5613fca4c979c5bfe9d2ea0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf59c8eb09a84513bb6a43856be04fdaf8c4a1b624434e5742;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf637322fe48db121fe1ac4cd659fdba4731c6400bd8eca2c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a14bc8b70dccba2fe66df6319297178390d51fd22d896a63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a35987f55862c578485fe18a6a99bc2cea329ecd3b9fb19b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44b51a1835d4dc7eb363c27b8c395aca89863375c73c86b82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f3555ffba5e003ada7d48f882d16f6637e277a355ad274c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2734bb4a55756e4ba1883088afee55d71afa553c732b4fe7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb88cba9bdcc5a8163d2d6a6885eaa8ffc3f8bd6f834b95bbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88772d0e8e770e8078cc30e234891b2b2661349791df8327e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h342ffb355652dbf1715036a5674a807502212c2efa29da020;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae3a1b14861755aaaf893bc7f250cc097181a2c50c74122d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd3357ae88c9a3c1a0625277c673f523514e02d7c6fa7f18e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69d931344161cc5aa20f359b2d609a74c6f492cea03aa8493;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd39e4dbfc00c71b64cb017194cf75b052fb599817b851d60f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa3f6471c4afa8b06346f9ce72501fce164e7e99fd7ef0373;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0edcf45853aa6366076951a07d611eccd7c0b845b68e1ef1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd86c871e994507ea98ed845fe704db234bff5488f3ecda2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3c768612e2054878d5891dd379b58691a03bf93bac74d1ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea12ac83d3ef774aed2cf0e235e48df07a8580179cb64ae34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52e3ceba89f8d28277030a8a89bfdbe1fb48fa38421763c81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7140ea4e98d88d84d7e42c8e102467d1e66780cfa49635fbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha76b58b18ccccb168537af3a90310812b2c810c1fbdf6c2ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7bda2716dd443572c8a91677f9fe6e6bdfdaa8eb83c6f07b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7955e6c5341c880155bb20b62a56f1ddd26fc22438f6fdf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4a4c4c02641c008865044fac0578168b00b74bbd69e51cc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h869017eb5279e70bb0349952984177e94d96053bd3af9e473;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9b7f34c62e5605cf5c7a1bb771e81c4cd1b758835263a32c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38019c345af52d9756f582d98735c1bb07603f47983d028b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18cf90f28356d5b62733b66e397599e399889f54e20db3455;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfc1b105c5ac72ad34aca29ea219cfeb9fdc00f0b0e4fcce6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29323fc3b98eab0fd33cb57bbb6a50d63bb4385038432a9ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49e4020ca66f5b4601f5ff7960e7663cf5788146c2786d664;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eefb1be1055aa10de18b8bf53960cdc8239b7765df5af022;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67d6c8b798bd3ae1bf9761ae36f39773ff657eb55fa20534;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58fa642e2e34dd9632eaf96408f74dd75a7237fb6e50b58b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h234317011e5265b2757ce0c5e18bafc436377435be2afde51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba64b3d846f89bc83ede2a861963e8adaa040106035d84f7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heee53041e1a9ff03d621eba941cb46288e037adc321951b2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bc9783f44bb81dc0c9de8c2ab818e09a83f7def8efbd2cee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he683b0826102f8d622b28946cfbf9ae6ed7177442fd3eb29a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h227f8a44e9271e8933e7aae7a2e1ff6780866b5ffd4948c29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1947e2ace59df6243e1e51a6b63558e27142d1f65b72dda3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7503a378d362bd725ee7f39105e03e5b023ea35c8282b574;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf33589976929077a98b3f6675cd82a7e01c6a1d600f53b9f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d5d3ae6b4710cb9ada0d55009995bd0af181cbdcd7f0d751;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e01c01806dc188569602d3a9028c11c3a1e6e99f1f6d49e4;
        #1
        $finish();
    end
endmodule
