module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [31:0] src31;
    reg [30:0] src32;
    reg [29:0] src33;
    reg [28:0] src34;
    reg [27:0] src35;
    reg [26:0] src36;
    reg [25:0] src37;
    reg [24:0] src38;
    reg [23:0] src39;
    reg [22:0] src40;
    reg [21:0] src41;
    reg [20:0] src42;
    reg [19:0] src43;
    reg [18:0] src44;
    reg [17:0] src45;
    reg [16:0] src46;
    reg [15:0] src47;
    reg [14:0] src48;
    reg [13:0] src49;
    reg [12:0] src50;
    reg [11:0] src51;
    reg [10:0] src52;
    reg [9:0] src53;
    reg [8:0] src54;
    reg [7:0] src55;
    reg [6:0] src56;
    reg [5:0] src57;
    reg [4:0] src58;
    reg [3:0] src59;
    reg [2:0] src60;
    reg [1:0] src61;
    reg [0:0] src62;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [63:0] srcsum;
    wire [63:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3])<<59) + ((src60[0] + src60[1] + src60[2])<<60) + ((src61[0] + src61[1])<<61) + ((src62[0])<<62);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he86b22465ed631b1b7479d3c396abe6ad9737ccc7c6ddddf2c0384af2562063a267b252da9e86c5cbae86b6a7cd59b75faff1455ad436f3a096cb90601f7011e7065e6fc3e0384b89ce418ca96b60e6882f4d69b450fcd4eadf16801f781e2b49725510d7d59e953e263ba3195491133d3f56f6e49b8c4dfdae2f352eeb1404;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8200f4d2f7834d67a9e0dee37487c81683a9be824ef326250a5506cf8531c630af9ec1145931e3d93859e7cc9bda1805cfb714b6354749290a621d9626f2d86330538ac5ab818e69cd197e7fa95283ece435207ffcab75091252bb3ff5e5b2993775dfd9243d744f972236cccfb0dca26994f4f43d383087158beaaddb6af260;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb834a0cbc2414a154f41507fbb0b23f7aec83ac760f22f6319c6b0a259527de6143ee82222f79216a941d99ba50d2a404439632a72772a3296d42ee802d70328f4a07bc8809a57f4a776e766163f6d1d600adc8b375dc94578fe894347090cbc9a385c27199e44a67c37f1bb73d096b52cefca8e4bd3bd65fab1a2391c69ac83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e5cabaef47c5e0d245c86f77816db4b45ef5718e96ce681ab8d5e6558de0f47161f77eefef9ede359b62e6f72f623947a9637a67510c5a5b275483df9fbd5a9de0a1f77f96e6922b8d07c0857d5abec269cb984fce4565184f8f01ebac6d16335837cbcc7ca74b30cda32a923e6d2432fb55c2335d204caed9e8c9b0e29e990;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1759d92785500ce66b882b54baa5bc7244d127741f7fa15850f797253abc569e4ca55d05ca41647bf4079288d80ba761ae6d5731e27067087bba30a1fdaecfae8bb0d085243eb40f094e282644c07cb7add98ff8202e130bda4b1975803df825b77d1c951d84accd832272f3af2012755ee7c08f8ecdac4434f5fd079e96dcf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94d50503ead899f4b67a43e395d3a8a54c745ebabe437848741071ffd752133beeaa2a3df9c9e8f61df0c47fcbfc2947f77af004107e631f3988fd4cf468624bc88364c3ebb9c00e713f6d51ad3a937ad6c01f106341f13fa4d37d14aacbcd4b221bb63c39a16473ad78fbbedeebe43b0c069c886eaf1c45f469f6e0600a27b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa3604b53795ef4c1ec9a9d2f1d9f521d68468dd1c754ce5aa40f1dd607504a0d32dda0145836f753b75fc14c304d179ae4901a8afe5d03dd3139f006a0bdf800a6a6b05c2cede6cb785e2d54981d872db0b018bd5ce34ede3191fc610429daacb89da9293a393b4bb60477bc0c9cf105a840ca44302513fe32a7e72be7ba041;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacee229e978ef50360e89d348a75692b0fca3269e259a96dcfa237c19f97fa32a5187e2381a7f213d02bce6eb2ac9569d5108a9a01fd69380a3dcb0abdee1e6ca82c59a2df5a8f588adb75c1fa8f3d073f35263623ea0e5a1a8d681054acc244584064d9226ad68e5703d16bc94c3b7ca39bd0b618ba51eb8ab45ad57a1d45dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6df3e0a3abf52194723e283d8b7d31cf970945068943a241c21da8a932be199136995f17e2302b53bad06d852286d983101eaf5cd181d96ada14145744678326480c7a83a9dcc326a7487db4df574c88572521a0ac5831357a2efb71ec85f86bed38db7b6d3b57457c02a8abe1771d09901eb722afc7f41acca69e2346e090ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f80368d01ba43edef8148edb4078b85536d9845c985a7c006d80acdb2fec7a3d1d050a95de58c8bc30f3c5a77d7861dbc6e694b4551f9a6e07de3a2df9f90649e6b1d0003fc25587f0792151575ab28099f793a75120383d11aa3e988457d5160bf5a3552b321572d1d2730a8c596636c06b5c6246425e844f523602baef1f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaed8609af0d30df5da8a8ee66c4343b9d0d83d3cc752f5f6e30f9437828839fa9b9b3acd32375f61ca32281fca9b1bfdd7e06cfca3098630d6ed166a203792dead37068196b6672c81ce9d19f9fb5cded4065046f4138a3b47e37893b0648e0bc67fd9fdcccd8562d0cd2df15b4f7b5c16380c6538dade20e7c0f9a651950df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec280dc9d7386ed9336eb412e7386225f4b0b07d6ff384f0ae939ac3b4533b3976264216663e2e186f0cc359cf386e85a5da864087f925f91df880e509031d70ef497f9b2b1b70388a6f16de39c1849b16c674bc05939acb0499ba0690fa5c563d1ff1781859149777dfbceee2b2b5dcbda0a01d512d6427d9153ea3355c1e91;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h793f5f0026227b7c897f97a23328e6723687a0a23a985d4401b80e6e91d133d69e09ae555665c88cebde051274533ebbca21ac8046475e37120384210590f120ab3125ecf5118b40bac88a319c8976efcdbea5a70ec1781f29720c31b234045c58ba93e7dc8999d528d6935f48e3504372f24006a77b39723323e873e695057a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2558f29c96e539941209f84d9f30c47dc204d7bfeefe2b0ec71866e365a68b98f42ce9fd2e55d4534cca2e3f5c8d1f6c0ea7ce3e22bd766c75a3428ad6fc98274a3c29d5a756f26b826e772404a41f7853e54916601f136d530390700cb7a8e1008ebb1095c38eeb6fa1ebcf59c93a66474e424e1d9db840065cebb2f4f063eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h800489657e7b7aeb6ba7bb2dab9670891921c8f63bb9d77eb5b3b1b199cfb6dea54f63dfee2202f478705429381e2b90cffc9a86e9427d054f10eb00ec03a05ea66ad97a03a735340f5d16fa5fc4af2011309756e826bde0249dae324431adffac42d9d23df4021f20196fad4d242c65f26fb084d3dc3a650b9afc125974afb8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fe4ce49f2131dc03b246c23d806851b4088b7fc95ceae9b462e84acc92263f5357d2f3b7c7e5d5a73bc67ec2bd19556d8f442fe084ab7e8c2aa1bbba255f820f97e9dbdd7ea21f207d8609f47f2f77353ac82d5e0d812dd5cc7366a6892b78e403d91e45d8088d023bdf294ce7ecd9ccee8bab96d64dd225cf399e3f18db81c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95e1e7600af2328cc30afc3aa8010e9eca8914d1c64850fdc03baef0ae0d26fa33227e66743384df5f7bf77d850c899fae9386c6307ad7c303167a9662e8d2676e8d4121efeac9e13c1cfe2e3fbf8e63c5dad5493233649952aa5b597fd15fe51a71494a97d7aec8b03b9472b502c3c4e1a2901c7b37757a1a92db98964a65ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b8e3de8acbbdb507ec54007716d771e035a3549473ff4f6484721eeb02c8b98a8c66bf8277d15db02849e2b12bb1541daf825ad951b60ca79f71f1d6b9cdb3d87cd75f9bddb081eadb1d06c11090bdbf7f677a8d3e68de8d30c1cafcd8519f065677a1b6a0d74a64c8f44131cd759ed08eb8478fdbf1a5a8963ae6e92dfbfb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h835d5199e9d577e6a8c89ba7fd1bcf8ead7fe2eb2d28e198dc8722d13613116038fa2946406d0917efc3cbdbebca0d4fab9fef1c5cfacb75cea14854343c4968c6190a1e3cbeee7edea1debf4355a3994bffe016bd80fe9401c23b420454b09a2d44fdb8202a9654910fb650151df3705b8d6e0b7e305509ed1c6467ab3203a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6abc159a896c22478f0d0476b2fc44600dca76eda26421606558982cd02b9fd1f7b2ce1907d36e54dadcb34ef4b82b8cae0dacff700b02688ed8156d0b6abd69350d58ed226fde2d824bfb23d69301ced752827659b5d7c460b29fbf7741e6f8c2b1d1af5b39ccbd798be40d66a00527561b1c7e3dd71600647cf071f7d7d115;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0a664233e76a6f9b0153f24963c39b8339dc55e12297cf19f3fa7138b78a63c1be71262871ace2f8914c88121b5a7429751e83c3cc1c8e8efb39382dedac10f0799b69fe1d7406b5239bc99bb70f2d05229dc6c3a807c442cba51656915467c2038b5f7bea616e2c15b3f7cb53e496add19aa4f6144cf25f7603168d76a14af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83b15c25ed7a957f5bb5440f590d1597600703114c9288cc00f56b3617531bd131849211c5369d70c1a5354f225eff729c8455e16a3f97bd7d665b763b4e64a1201e20f3533292f56e80674eadb7c366be3d96e46c1514aaefb110a20d76a0f9e67825477b65964f4b9757a669184454044e99f8d9fcf67782f169634cb416c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26edf36d3d60fb63b9520052a62212518d0714753403656006fb40bf7b2c24847a7e8071fd2c387b45be2f79896a73283ecff8ad68cbaa8459209e66de74bb26ab3b20d7cd6085973c63cb6a0edd91c0a80eaeb52168283038ab28473b7c17495878a052b6e1baaad6012754b22fba041c48e7d944f8474df51bfdef84873905;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h502f84654501584b5687fe3260922f33906d97b3685ec9dc5a9bb109e4aa8359d410669f2104794df41878459ea752b0f5824a65456bc1889c54c7a0f71abdfb88996e7f1ebd7bfd245299c4e12c61395fd7bec0dac20859339b25be9e7222e62d00372d9505003120a96c7a2e0400c17bd7c23ceb8563d38960cbd8798e415b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2430d64f72273021bd32233226ee57719c914df889d30f7525d166703bc2c693530ca680423dfafe621b0a2dbc1e0f5c5cddb3b635d8e895fd17b4d47a886acb7a3a7428bbd890d8422e26b9544167fdc5163d24562f8054a0005c3fa3c665bb3856e9ff68802bb727eab76a5cc2d303b0737a7040fd0aae491d2f2a2d7f047;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8a951d6a8bb04b38fcd857fd3231a23dc10bbf563ce7e6dcec0543ae4fbc4767b4a1db4a8fbda8de3f6b6463b819e5de07c7d8bec1b4018cebc04788457d931bd0e1f1ea6edb8898f38c6c27aa3a5770224f780d4a18298e3867320109490013fddca1c70137554e95e039f22d4437ce4d1cd2c1a1661ff7827ea364438f6f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h632a873f664f82e380980f7ffa64492d36bcdba34a711ec3879367e974678f1d514141a3e2c3c3067c250b906eae7183418ae38034aee6e58e89652d90eec1a02b6f31792938b1c089a81bd694887b80e99af5fc0ad89155ccd8fc0c33c6c141f98b747dedf98c4fd7b83e6025620bacb721d79ff798229a0de8426476f9fcdd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc122d0b4d5efea22e6c8982eb4d1b8f568dab16e34fa62bd7ad090ead9ea28a38f89cbd415707609fa84a3b014777e8644acd220f480817f04395969ec73bee19d11aa6c0bc6a9be35ad388c87ee7bdafd713ed957d04c80cc6c07012d0844871786fa155813141e7706d2e247e58c08be2eab67a6bb82e0cf27b777785aca8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0f3f3e924c9c76524a33b834694b132d5932347b9156c31883dd64aa5f08b4bf1b4383f7a5bc08dbebfcab3c0983231f915b5cc392817fdac09d299b120f1c90049ba4c57a7829b9bf9e6f366f485d5215b0963a8672c1ac6cb40fd634d20a5c79fed2108ae0397b014574b4883af64c2746a575a984e3f99d883d4131058a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfd338805eeb8d1a24038e159b7e0e287385eb1ad421d95beaa9fdc0791540433506129da815d82d4cf0b6d264df90bc12337713382d9104acb4fde45c18fbeb6528acfa79d78474fd1b1f161e8d1b420b597a71eb9767ab6ec045e9902581e37f59dfe048272f4e331e1d7891a233a2e98188c79f288871160dcdfc49c5c963;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h732cf2fc77ebee3dc5fbbdeb14b9ea44bdb6d0efc3bea06c31117623d5673b1fc3cc563672cb3d87de1042163ace3b6bbc0eee3abf1d4d08a098d6dca3130c4ab8486dd0e15416222b7f88bc8a869fe9cd7ba18c465ec933d607a1a986140cee707060e14d64b64e7adf0b52c388522e7e01305321fdb26490da34b32bc80a5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63ac37c51949dd4834415c2db0493063ca51a7cee6736042dfdeffda7b95d02c97acc6a85965b32ee2be42c477c268bdabbfca5bddef6d10dd8b89e3e6e7fb9a4ff30eecd67b080158eae317bc62222ffaf05404f3eea8999c5ca28345b778e071172ae2b9a0ed927b0b9b84eb3e2f76096a648b8c16b2905c4b05dfdecdabbf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1740da8a467b928ef3329792a3159ab95cf400395d4b90ad2405f0e2168126d87bac665bd2f01cf7f9fcebc0e65893c51888af8736adcb41c5e27cddcebf2a5892390e8f57e6c5baaa260819c648a29a7b12c7ba04483ce9885b8cc4f23adba2eb5dc2e6f64d64f32a0366f5c12fbef62a1fb8506f36e741dc41521d3b6a92af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b3aa821ec5f7d625fc3e4f72510124c0f5910c191e5a9d528c8f4d29f409b2720fd73b5eda56cd94ad688452f2cceadf3e2b8481b565e5548c263a73d3927fc517ec9c1bb2d8ab06253da456f8c64ab25f50b1604e6472c084f68e0654636be2515cf9311419b2b47bc8547df23f6e509548505a18318012191bb7dee7cb891;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h624e38fe2355bc31ca78308033a05cbfc70e2ef045bbadb81109be9ea7b41830d080e6bda474422d80a17bd358da2058c7cf9e46109dd3100e2b904179bd031ddc5b8f855e36479d0874b4a9520e97f25cc32492bdb6f8ccce5ab47b421cda9adac2d34543656e5854ad21e22d185fc0ab5f1e5e8da01ab9adde463626a66edf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd51139c7e20eeab593409f2965be9de654c38eb81a51f1c575920645e208ebfbc88b5839410afae07a5edb9631e8b804c5cfc668a0ca636f2edbc08125947212ffd69339efabe3c1cda84e3cce0ee27ba04a9e1310a22f035ba8a68127bb1ac05ff25196100261ea0e07daabb80801b73d7b0f3741391be058a901ae01936d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbdfc46f581ea458c1136c5c2d336454920ea24eb776cf0f68755803139d2f0bbed12bb35b2d88f8d17bcb77291be6efc63e7e351b80fc69a60925bac2db8f921eb011d55f5ee44b2c8bcf7d9a41b7f78d2d6bdf17f61a54ca6402d32ba77f62ea098b4536b9fbdae00b600df5d4ee5034d5f971a003ff622105b8a45a1ad312;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he95908d4da67706967f1546410588a95b776881d5340fde95c05515c27e768c1f2a5589e31cd1d75114f02e881b20f9456c7bc20b518f81534c911c183708c8a03fbbbcec08bb9211ce96a21914270a097170003feb43c5d2f5d594128dd78933855aac9815c332b3bb70ea48d3248d012dfb69faeb66e7131b716bd06b6f2db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ca1ce5f186bd0f659309275ca6fc771558285f59090b6366c498c571bfb7b773683ccfd5b7543daabe3b6cb86323fe25e14e2950a4d72cefed66070838c6330a14363160d49737ae46f31129260504f3431a2cbd9d38d288b8eb48b7b5eea94ff48d92da7e0e3fe8f9ff2dda0a611086d632eff260e773cb79d886cc0dd4726;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d70fb7651f8ce2340a8ee476f5a964d6fe1e174a6fa7398561b1242ffe944799f76195c4b27bfcb5b7f56e65dd05abc3924f09bc897bb53f1736528b523caa65cc84d6ba8c89c8c28eb2fa82e0ee95ff8e57c9a30def3a33c1601d00d4e77564c8314c6a8544b41d1864ee1ba1df1c377fdde249ed7ce134db9fc1760eef622;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1eafaa7d56c75ee40e4f8692f760c2d21739a1d09caa453f0ef8ca412a14725b950152f3e7f75a63622078ea4da7a23f0b8c4aeef591a07e6e9f780dc1213df14087a7fd1015e7aaf1d594cba5cddfa16680ba48b0c49e90d700659f106740cc0e9582cd04f79657e7f175a31f9aeca7bcd57d8c7fd2e14d10745a96833c77d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf011a09b8adaa54adb260d9ecacfb5ae568b2acaa9c1809ae45cf69092317693205659cc682f4c623883613620559423ef78abf290558a42158ebc422c141863aca6e21a332dbc32945aca0e1215b524e8a224d48fedcd8273803da26eb0277b59d3775c49f5f558f63ddf8dbfd57bff55ea9068dd4fdf09013bd8c4b4ee89b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha922df7e7e667acd01086f598696aebb286e662e20733889622e833fe44e9a68cd4f924124f0e0f11f975841ae129b9d37d17e8d20c8354f6ecbfb1278f0846846009b5a252f615231649a30fd7a2f2744dbc24a68a9a88efe5d5cb196394fd6d374a7b18e29eccbb7985fe3f542f24614eb992a3651a6df3373f948e52a01f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h617a34fb66002409356b02ac70c38931a2724225ec8bbe8fe58e4665aee9da6e7de9f1e76b0f5e18f3377a0b1ece65654e81b88222251f6599591b31863b9fb18a2704b87d5a719da244ff7b59d40bfc51dfeb6c4531827e736aafb242dc3ddc60420d9e887f72ecb54c2a55fa40358dad401dbc5e1785159e6b6116c2e80cfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7a47e10fc30edf3f715b85acc743d694aab2c514dbbc282a869db0f6c287299514ede15e00197865d64492b0ba7b083a7b19cc2f0f6c77851f9f914eb7dfa757b253d0e31d3777dc4ab99081157409778a2c87a6c2e1aa311124e075aa5a8958d9a8eba5221cf5aeb1b4b177147c7a68454e16c8f2fc9833cf0d82202b2bb50;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8ec866a9b5c2a782fa55ab11366988e90391b9a3d751cae529be7110080d7dacdf65dba8a5f99f4d610b9fb03f374506414e6409ce68887257f954410738ef56b8e0b9f364a8232345045bec5dc5a7719f5d68f8a4659724af06d17ee1a9dbc10bcab79f1b93fc6b9cbacd45c8d501f3432f2273c2b9e3a39187189a4f5e61c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h120306f8a28fbbb7a71b8e739848c37e30a11a5a70e1a50a03370fb3370a7e696df3a20bd65da3e22c1efa2a99c883b081f691c44464958b1f50942e17c570a4ecca3f8f55dba46d0fbe94ab946515319634c7b50281551defddd8c590d6b49edb6b78a07ef1d8a689d86f768d4a1284fc64b0e78a18071e5d3182f49553ca67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf063c2c1c945c8553615f64905aab6ae89527b96f00a88ad77c8615efadf0918475c939e4d77eea3f2037ad69413f3b5595e8f91480b57d9ed15fd67ed5a8e3ce477d0593373de5de2680467a86b3fd2b60f12ad97425edafa763c4592f6c422a3e150d8ba60ca7554e6856ba098d30416bdb131211439e041b05d51fb87608f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42c6ffc02e02dee87c98cf916cb6d9270025b40374bf023f5ffb9258fcab183bd34c0652d47b7adc5bad7ad5b8f0f41584431785a82fa6f8b084293a6686a7eaadd348fc7e8fa60360ecb0156c1d3ef0f0ca3e71ec27966251b74f4525c796f9c343bb0acf2e0e51954e8388e138ec5186d7f276e03643b7276d4efd00ddf6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h836e824eb5b964f5900dab5e9af2f59b3927812b0ed8faa4f10ce7e533d0a026ecc9fb7e8f9dbad711a55c4f2222572ed5a2c0f59e1409267973f12f1a7d448a6211697027fa774631c697c219ba2e1a7ab4ad68d7b6e08bf4eb67dcee1e1fd3ff1fc0f2c213ee6caef46c078eaa2c4e31301de2cab5f041a0482b61ca34b084;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93132aba6098ca6475c20d951ef02d095d824fe53ff9c5337b81376a40e7e2cf3cb51ce5ab2a9a7684be807c65bed6908e1ba4dff891b300a2cb14b9b6a445492a0c416366ba130218a8d43fff79416a223925019ca3b959f1aa03ab6a294aa0f7110245b6759ee65ec849f5f6236270890c95bc3953e2175bf2b1b0dcce46b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc204b6a29db98e207a432ab4b8a1b474d76527ad77bd34782a7558a6e808f4db4196563f0a29f8a3859c2f4b74d86ec007b65cee7f7c0d894f626466514b26dacf38eed92ce6a8bf853c2d376c4af50d863b6eeb348e22277602257cc972d7df439c13fd69dcbbc916d4a861c2ababd5ccdef9b0fceb931bfbf915649a6155a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bc0c791545bdba2c6e5ec09ddf99eb397992266e37e93cd4c74c7e1a8f77e9c0056f43d4500d9b0c7ff0c6b34933c4ac9981b0a82be8b4acccfaff4ad35657d2c5414e424331b0cb9b451bd2562a85c5a10800cb69261b5dfe4b0b08af1d48c9ad917cba43dc66ba8fb12b4345f82f8411d7a19c6b376ade0d87f1f220a1715;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he11c31e35d24d832cff163b263d24180dcb1c8e65a849b54b0b0d7791a822bf2226f20b821f1a9eaf31774fe2f2ddb4d709de65f5db9fce175bed626b80fe3e79003fd40586ff5b4fa453dd434343a97da6d755a0a64c02ed4bdd9afccfc666eabedd7831c14cbe8a517ce422f4bcd8334068452bb57a0fe64a509f4495305c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6407eb8025daf14379fabc89d9a793b596f627a1bdf1e364ca26411fbe894fb23d6f4c6c0247f766175d7af2c2ab11699897dc464ee971d68a9de3f2bf17c915fcc22b012cfdd427d7bf591e390d2e2e410da9e206adf6f9beca5517589e7a3a69309dae679ab27e6d11fcb1d67e594b73b6db1cfa7e0484e6d44cefcc46694b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52132161339bdc182d96f15c5902432331d00a700fc3d1b1dca0f20e0cff12e3203d516fd1b82eb0b1d44abd22d3d19ce9d8748c6c61ec2b14147cf631986d52b136c4e7a53e99cf1fd7d39ff8bb5222eeaba6d6f066df460ee8a504cf9a9ab1a19caeaeb86521a25a0466ff6fc1ebc494dce8802454710bdcd846188de9de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49b236440f4d26426dab08edad1c095e6082779dd330407314fa39530e2d58a804ea949fbaef72ba18ed7adb8efc32ba82fe17baf45c3c9ac16c8be1281f09a5cc7f08a9ef8f3f466e69efb215f82c44f395f283f9e45d2cf9c1482391a04158d62bf137e0d828fa98cf34c66eaae26b8e5b1fc9c501e89ccaefb3ceb62e2c34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae9e1b62c61554f44028e591ec6a39baf22733dfc9553d6a1211e14019cf8ad549b06bb58056084ddfbf4cf882dcaa449df8cff5684ac65695f4d7e2db0adaf447a418e842d204e5631bbff24f0a81e2f94fc4bee6c1db641f0bfaddb290a65b1bca5709295fae546d5fd76fb211262a89dd8594a24a11e2eac84b4bffe7e7bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7b8169e355137cf1b596394481c649e6f478f4349ab12dd85d21ed60a4fd569c0c97228811aa73536e3bc49b15b3a9592cc5d91dd2c84b14764b5f470b1baf19ccd31dd73b27871dd184a5fc100de71dd8bf495e416a4b10038face8a1f14ed937336bbe4f5bc10e226e84a02ef1a77dea7a363cc81a53045af10a0de7fa783;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5e9fbd1c8b77c5f4dd2fad64885c737c52f98d5286efb65abd93cb084726b76807fe4714666431706ab968d4bbd90d9318222cc7a64514d4969c628b71c854b4d4ce2ae56f33844b41e09dd0138e4edf90307ad69becbae425446a56923b5f146aebc414913356ef6c671e1b4fce1667f20577f536640a7ea7efcd6a8687aeb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc47939debd0a611e1ecb3a03d693e26e6c3c0ccc5284b28ebcb98f8209d8f21754c248c840c3f356a2ea831e693c25bfbb4e069efd04bd428685f8ebd5c6493e7a0499c23090d7d7b5033e8a319baa1bfa87553d24ba9c39fefcb27db85600a3dc84b922a06ea1d48c9dcc94743b97e67b3ade9f5e5e2814b47b76545fd85e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95245af11f0cd32e41004e1853991ba3770d5b61a6a5084fcd6f3af7966222bbe35523226679d7da6ca52c615e5f570d37bb266c7fb72dd51ea63e851d130d0d012b4d1da334fa79c211814dc43d082095e15a7fddcb3eb1dd23bab3ddf17349f112db5a0ae626dfa46405994765795ba3bb98351f73288ef7d3aa3d99e6ebdd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4f608a6ad7d45798f99d24bea2947af6c722cb72d6ac13bcd7d430f6c54bca4e64e414af0a82f58d9b0a9280722ffaafd053774ce0f127f599182d81c084515ad2bc017a69e1b0c8b95b63491849ecc65b9cecba3bbae9ae3e063532338905259186e721994788dc28a5280dce38bcf76f95e6c46480774e05bdafc31fb1604;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h778cba9405800d514c344990b8113baf34ad516c6ada984b32ed9c0d6bf011a6e626e002700a30f6099ecc30151b693fb8594f1bb0c127b1880a59cdf302ba7a7b5e5b9d6fae155a4b6960f5446679bd871a9407bb72a7a06406127ae54759d9987573b03cc834a788873fa1acd113d886514179b7786fd0546d1928eaf52fac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf026dc9d49e0c3881a79aaecbe3c40b79647a34bf861a3fabc266ee4d6db86c3ddad38816f34750f16c59c00027345ca8d27e56c6bc3225bdf3973a545128dae674d8b64745a9aa9dbaa79d3a01d28edce0c7e5cb18fadc144e7d8ab6ac9bea7f4d4d8e516cd47fc7b667e88573e6d04a8e6c8b779cd8e246b7d79965382749;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha01e666e9328fd8f6f1bd0766fa2ff95994e3e94621920014eabf29e22abe052b3af402ec165316d1fb4d4e004f6f97037b81d28be6c05ee61c4f559fae31845b529bec58faf1bd8367e928e283bea2fb810a26b5fd416e30a842a7d4aea97f7ea7e56ad65cc4cf41ac7640ecc6da7d882c1b0de8fd114b2628f4718eaa08d62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1f83e739a8830b3223d2ecfed5eba6ff562930dad113cc48374444d4a942e5ed9ee6d5ec1b88d85257bcf43195b3796185f6279e3af1433dc8e213f9a33134cacff3eb70d5777f6e43aeb077be73691b89e0fad9653154d5449f9a7614b31e6ec266afeda1f7b915564856d1ad7ebcb12fbf067339fc5b3fd96c8f9e3aaacd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1620d0389d102b9b5c3741b6e2f9c0634655eda4900b03d7ed6fcd05b33fb4176b38df9d5b71a1f1c6b3458405da871fd707c0295f20d4e8a706cf04595c477e1a125ee90fb36e08a91f1e215ced5b488e37019c84018376c507555d579bbdd54a278de53c4424ca261ce8a43dd85963b9db75a9f5eeaaa186a90ec0e7db5bb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3742f3adf37960f429aae45a117e28cb5eb8b6521532b2f908af00837e9d54d1c60e980be84cf2e23d91a1baaa48ffdfc5fe734474bf14dc84878536664d2d45b1c202e0c7ee9c2d339bc23efe7e6c24d9055539beff283986124d31e4ffa38f0aa59e3986931812d625ef04b86ae58278fb5c792e8d8531ef3a6b59a5aa3a8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf8666f7cc985c51662ae4cadd45da5cb3965bd757769049f8256d5a6c8a1c4b85a1fcba20c4bebe5ccb4bd0e5be205d7bed44cf177f5e2429856c58d41bf8454fd8a2b175c2f17ee4b8c2ab4ee987f332f60fe309b32681a8d2abb285c1f586e48c1769f4cd68aae34215b4f0a54356f6a83f065b110415db7fa17f23fedfb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19c7f9d826753a15db16338fa4cb3341354a726bad94c9dc05775efbdf69cc9cfff6185d30b233a0d39a4f2f1f24866ee697b801fc5ca2df80f54508c6bc561a3f6be4bb1f9a36a205c59771069be4f293f08a828a499ed16b5d0a279520f7ac8dc8e298a58ff0df07980846e774ca2345a169ab4b7b2c1cefb0d8f051d41c56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55b919807d4ede63ddda868be3224f39d162fd59eb5ec268e048e231c6abb5dc37e57b8ea45ba49cfeda954766c2312faacb096554b6a9de72f2cacba91b77d8ac78a87245e84106ce7c589d3d02cb25f1f8a6edbeb67df96a129cd013f72a270aba2f7ea03384d38bd4df8a90a87edf6660139d6de0860bfbd198bc9b20727d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d771fe975e8f2d17b01b4acfe7c71b9b630d5bb6b9a00de51efb756b0a7454153d0492d7b445b111e6d9e18171ead96b1455736cda66dbd3c43d02c74c638ab1c6f464141c740663c0e08827c7b9a9d70c6585b1f18dee959db5f9df881cbe5d10f71ca3045d8ec6bbf7da2a6f991fd41e51c63d6fefe81c18e92f56b761d10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb57fc481b645a7de158eec62ae9992a3c586e76095d2c373f23cbd73594bd5be2f8c0c8f03c7b4e3d8a83e3dcb21ebbb0cc7fbe96c08aacdabd9d764450bb4fc38fee9e90dea8a7159125c79d72ca0a1c02c603f7bb05b9aa08fe079bc5a7cb235193186c0cd5f69c976963a52b2e27df58b5bc5946726ad12935731fea1d67c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h245aba2c6cac6aa52f1693961c46d4abd264a51715c849fd8268345ff2a37ffa140249fcf238bce750ce99f36aa8c7f35e26b29af718b1e90f18479e92a10bd467ce8d7d122b37168f127a7b11684740506c4316f091094881e0ed5a35eaaf35debfd61448315bc257efe243baca28e4c28248087158fde694d2a7f58fe671eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae6a36b9e2e14d56417130af4f3ca04ae1aa9513b5df956392060bade5e128bc1e9f53b9eeae49d98bcd13cc4dd7884d17b6903f8082f4e78128c52334ba4d6dd962d4428fcd25ac4d7f18bdde02e729620678c5c66f53f2045cabc9fe0a4843f969cacf6c3d65325ecf88e990dc39f2586c99d2c1cc770b2345950156d24825;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c7920c68a467442044489d2716d8023cb5e0abd2330e0522735fc81e2094c3fbaeef39390c313d6dd79dcc0b44723223f7ed37f2eb7fd70cdf1e92e5ec0127faad9795ece35f3aaccae430f3b2ff6d2ab1feea90147ebef39b40bbf539ea2c8d1a44d8fddce8303bd5ffb2f24c2766e49d81b5dee52428ae0376525a0d39571;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8eb75ab15a7e71843a861eed2295ad57e67f8c71001c4520af23a9b275d9eacbdb5ee4f01be6b79be1ea64d0358cf214d764853fdcb687786f7a2011f8c7e6215e86fa3cfc4be2bcd264b27681d0392fc3249d8db1ab53e3413da1c41d4be266aa757bcb33b66915890101e194614ab17ff8b7a093f089cafc651b30799cd097;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3238429f5d54b173dea8a554d2ccd21fe030714e951489f9721d38150a9f4be6aa8975e4fcf8d87143e1eb7f78e861201c3b0fba1cde0acd34ef6ae78d1ec866dae294f9c79127f72aa8caee54f1870429e18fdce31969a2582df9111f2d42840eb77d6073f7e3b580896693a15a3cc92bcf5acd3df1e197c84684a52d371870;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h417c3a92eabb4f88613223c616986a7ee8a7eceaa0abaf798d87f534187d04199921350f11451d8bcf9e29677f65646d5478ab38221bd31229d6465c31f19c2ac6e1ed9469219268ce8c852743d98839e3161d776e9f572a220f38bc40bb308687655009f347a0ea218ca5abc1f4d732480cb4528268a114d83f639ad29aa110;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf138310a7927aadccd42067c956eee578fa95997c0d719af1f6121d29f634187c0f3bdd9f3939312b3330175207e898ba7d8951012da67907af643d2758f5570c514f059daa87e9325be9512aebf70eded9deb67796b089b954d3be5c2b60808cd97ac23fa571160a1074b9572ca55e1b6c6d10e99fcf1f08fd8f46dcf6ea29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9296134eb08d11f544ee9b5bf58ae77c494ab3dc3919d6e1abdb3a9e05b443feb23663b4a05ac9645efd68721b4811f1334179fe3baa59f3d2e6a7cb8045c4769a7a9542e5377c918569e8450f6f7e3e84405702c5f97884cc12ee63f8881888da7c9d08711a4cf9b6f73d73c1d771f18af2592ecad293942557b937997ab49c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83e6bf33413d5a426d8076c57a50eedfaaff7d99bbdeb29fdd173e6883c7773a9e70645e39627cb23b7c212add053af114042ec1033ed286e4f39085466ae883254e249313f8c3ead4744a9800f2f28b3c3301ece3c554771307a4f16c97becbe1a3ab53dbd8fbfd617aacf715e1755dc7afe0a7bdc6c9d7c2feb0c76c35c388;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1524dd669a41a52fc037d8644849b5cd381c4dcf7f28658d178e4686fa7083c5cfcb5ddb0ce2392307759d2a940783ea1fb5d21bb78b9161bfd299139718b57a6aa9ff635668e0f52c7f7472c9be7823b351222fee73ec5becfbdfb287e6623da56a36ad635a3b680f068cf04ab5c19b98725d297cce8cef7b7c773e02596436;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22949b4a50901ea940d601e90101214e7c0b144cd6c5e2874e8ecd6254121d267f27baf266c690d90a78b950fd85caec4cfb7a930cc200317291266fab2a437944ebf70d6c6ca22cf9605483b8d34c3d30366e252bdb53b0fca7c7240956a7fc8d3eaeea0602056c91235a0f6521987c16c5eb55b0ceeffd5e73242733692771;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf157e1db8684d88689ff830063d43d64879bba0d92eaaf0a5ab9beb380598d656679273dc2574b047892eba1164c8c07ca3492fe28b3dbf0d5198e0bba3a11c6b2119b815260478abd0173cff62f3805bd40f02c5047f1511b48ba5a546123334a94f1d6c02c1df1ad0e694cde77fa3771bfff1100538166a755f32c65cef70;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93e7bff8e8d69a946573d3e4cbe1ad0ceeb49397c55a1da7b4ed41a76a42ace4dba519dc38c7bcf4977651de64565a73d52e5853858f794cf6e463d281866704fdcd5b784c8d557a2b9de5157f259223d75d566104db5f8d8c5c2b2a3a4eb7c2843e3301b045385bdfb2534182926fc0826f23cb2d564a0884ceb637978c36d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92abc623d5d1e945d46eeca211ac29e75d3ecc28151509204ca15af7bd26d2c08fc1c15028bd0b368d6303bd85bd48d69943631315ff3d0319d62681422dcd6d061f7d2b6c8d08945508654b69359721536890738f6bac352712078b0e7d5986c5b89447a1ee0e0e830ca20b88ae67c11f1d635ffd13b35ecd7e1376276a002a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34bae4b5fb6c93b8c4f5da3eb353a6f88509b68b5f1cee598ab54e342e6b69780388f00d50f3a12a2b77df3f35fa5096637990cff9859a2d3d0599cf428fe0bd79ac2155fe48b459db67d70fd5205419a7a028c9a541893ef9a8fbba917c9bf102d6c98de1b01365dbe2ae634e2cdb3f7ba85fa752c827ca36f7551e21ba8b3d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5d9523d41e329e3d8b6cfcfd31e176e8a9e655c6eb6f492cd2e593c8a87f7e955cfb0ded081cede8bda9f4702fa6552060af4cef541391ffc695ca6e1c92ea7c7ccc5932979d0dad5f4bcebf115cdb110985057c13b61fe7eb3540e6d07918adb8a9b9523fb9c55fc4c96ee5c2c2265357d4bdb4a38bfa77e423ca7fd7c2e8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heca8f3cf11c5c40aba4573edae5b9f5d916fad3cb27e91423fda5ccf2956611946a76108acfb9235c436b6ac8b0bd9e6a69fdd6b19d8fd7d704beb19984ea9277c328fa052e99cd8629ee38712cddfe34d4e549a3e2726ce85f5d6695126446f553bfe4f922d37b17a9c891d1302f035f630e0efd2e2731f79e630d9dad59289;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h404d9b9939e57d47a1a4388af6026b7742b761c37492e785c42a798f158ac74edf68641e8e24ca1acd6ffc52b6581ea3fda9ea67830420351bba2f14edfbdc329134c836d62a59d3a6d10791e8eddc9314c380f19726ddbe297523e1a590b19cf7b538847291984aab76dd33307034fc6bd82151633c0a873b7a35b09db643ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3110e2b3d5a855619205968cf21be47068a64f50053bd5ef61445c919a57058e79607d7c87bb59c675fbbb9e91b3a8ae675ca6e2434257e3db5ea993f5fd7939465a6cd85ec83b93ecde2d04a3ba9abff3363ca5dca45b3c8a18f79be681b5a7de39cf8757c2780790ecb3af08355cb286961fa0619ebc106cae45db071fddc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20e526678e709908bccda6956831ae3fcbe511ffdd8410c8f8468ac92830ef7232221635f20ab4cbf27db7e4905a12e28fb22d1ac8fbcc8637cf8fa3b8a9b6285a352aa3bc052ab863f7a9a658064bde89d92cac29bd5e9639db628fb1dcf2955e34c62e20355af3509ae92bb4822ff1086b626d91313528c26fadfbeb57c9cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85165ff38e4ef7cb8617f03254e5a987b1048e1ad5e7564a558b3334a09025aa2d3e757e6b2cdff3913a972a9584790efbdc8cb59644202a7c0bfd6399f2d13bf14f1260efd53523e7041eddf47ce2d296bf86acc54fa62bc8689b8f9724b145676b5c506412e629ae1dbeddf83925edcffe250c65032a47e61bdc0c359f9f1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he84b79ee6b9121286a3ea718f590ecfbeb0df9688e0952baa9af3543002b4193fd0ec1b00492a52102ef1fb25e70e85ca50376c5a678e45e8b2c12d433d38f85f868f8e858dff962cbf9e88484e504f27f631b5a5482a2c7e4bb5126ac300188b464cc866694579aa2e656492312df1a193ead532dbe4474143998fad59a15d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he14bc347390bee39447a8bf51c524883a78076f754c7ccd7382babf92f9caa015efd92cb41c142b1d998eabe14560111d7791b0e3983ea954c48e597a816bdb54ae65b474757d6a1952bedaa05881ac853d15071ead99011b0d64185e80acf7cbdf67986a674946f53977deb8cd9c48f3cc999bc44fe96a4ccdc212442edda1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35f071599bf2da59b7e960094d27f9a80ba9ffd42591cc30e86d66705cae4585abfcbc99f535eb825d327d95b6ba1f015c7359fc12b358d3d51aea8a1503fcdc960abbcf5b58b31f91a00f919acba4f2b06938b90f533e09536f653d56cba25fc605f2abbe9a81394db41f286f2b5dc295964a748b0fadd733c802bf46e65cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b6f87a7bb016900e56fddcf6881540abbdb5bfdcf346b91cad57239ef05670c480c0e8476204162b4e2c026d1567be3085735abaf1c2e52f7ef2598614ef603c42a00e2aaa05109959012270a3c31f02bcafde33b581548eec4a39777a6d2a8c1cfbd889463691768a932d6685515246be4c8943980638b8104efd1d39ceba7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedaf6cc0ffe24905ffb66d6e9001d2e954fbcad9c61d38be1506bbd8037ddf6c6e1b103cdae0f0cf7cbc0719fbce972053c5f5d665b826bd510b3e55d4bd1f9d59a7b5b732e9eb9bbdf843ba5c4e533040e8b175e6d9a779a9f75f2b35c5cadba4ff25df155ea5b2d46bacd04d331a5a68935ca057dd202e8ddee6404bb56f03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h801e54c86e7a9039d0f7d97dd525e8bb468fbe1a9931f17b294b4933fca07a6a4a69c57338e909c130e79c2330fa8db2705c7161cf4323b03440282d5fc2c101b89600e45f32da076894209c1bd01bf758773be605ab6b870878dc78bef42a3189861dc62f3df9714066a8c4ec2695e4695fefa516bb465a23569e05c9eec121;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd12731b9fe03e78d8f399fbf2e494616b9254662682984ecfa267fe12d4f85644d03665e8a4238cd763d4681ab7349411bf91158d252dadbfee49da382f15f3bfd79af2a31eeb7b20f6255ace431fde658ed029e4bc4eaa34a5fc594df5f3dc9ff2f622b1ff25c9cfd111e9fdf3d2ba2037c1e44e801325e2fcecdac1bbc2ed3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c0358953ddf1d6975d6e14d0e15a464d92ae05565198c5b35c417820472659d7851435ed6377e2056832a88472ba9444d6ceed820528f4b18676cdcf9c396ebbe06bae283f68deebc5273c3e6dec7d8c8008827cdf455d24a713620d560e9a2c8155e8279e123dce1093f277ec1106e510b1cef48aaa7ffc6667f513f7a0369;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h295b70cc46c49eb8a03f72619848347b1ee11995c97c84c341e359ea3fceadec3245ef568cb4dbced23a8c28289566c74a5928ec5b3249b8969e2f78c58838e99e368e69de881d40e81c25f8b0824466b796744d81c56bf47524f82813efc5349b6e5498db249b7ff4f71125e646203dca2017d471db5ce425d0095d4fbc6660;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20166cdd83daf81c5016db8c419820ffd47c795252f1be1f9d6f178226f22a8cf1780d8946f46fc90b5ac708a408826314dedd1663643adcee19665c3ce657382cb6350523954c2b1cf22b1d9792a742c3ac5fe0fa3eda683351a48eccada9e4808fe4008c8c9a2eec95208af84cc7cc20b60ddc138e1c3bbb5167b2447bce6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65105ef6ab832c0359f5c69b38e8c9dcb4c13a39e603aa7314431581e28870f61cb2517983e83ab7aeb999551eb0c636027a4fc1b73e385995d37c1ffa6a91e6bc6626fca17308e5e48bd52c6abc6585a9f03c3f84506dc60a912f9f338c9823dbe1862fd81da764906b5bc2931912677ce8dc0306168fefdacd23764e03f04f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae0ad661c65546ce95b39cc06dd11503c1681edf9c8282bd3b3ff165dea34b182f4eeee37080ec86a3624d6ee1df519e96874480eb0dcc2b300534bf26a1815c4f17a2f6c8c692208417aefd42e2121f560fa0112ba4ddb25e3e40994fdc4f1a025d05c76e0c6cb63d320ee14b304061bd842abe36b50e1bdbe4ddc250a1e7c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17a3a64c59d55cdbaf181e5bab00d93f870ca838b5e15714d1daf6fe3c5dcce0d7edf5b6cfd0e34b93f6a345aa4c67d0df7eb662278614b40a70242c045f2ba9404b8b9fc146bc062d2bac6bca93a1eaa902631fe47fddd3b2e1f4914ce8f92777608d1c5b0556a34b42dbbe4236cb7d539d8f747547be9a2c33a476c300ae15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f68b6333f9063572284671338076cbd0f9327cb4ce5cd7abf24370a5d1d5d0264518f1cd2eb727eec2c8a9460dc51683f82e4fd358e65e2fbd4c824c2db04c5ba0000fec1c755fe31a3300a08f73914478c9a762160ec4f4efd81b60c4e30833ce57ffa3f7a563f5458f8df4bd49fdacfae6df5b8e9c5b90efeb16e82efe7f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1e04ef361e5ed96926edb3700ed84a320ff1bc3f5d72fe5adf84e0022431d0a8efa0a29156740967a3d72a7e4bfd5f4a6ed1f9ce0ff103c09381647af385ac97b8320bde04b291c73ba876f12c64729d7765ddf858801c2288c59b9bac06ab57a5e86883e6badc53ac35f9ba61ed248721d073d42424882f52238e520dd6636;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81e6fa45b0e53b4892ad12ae7fc70e69916fa3824c6e324c62ec7ca0a8c7da372bd6df00b16448f06882ced3dff6d555e2a89da5a61dbc3d905fd59a255c6d1b67f29822eb5c65986c5b7313465bf1cbabd2c46b6033406ba3a24eb28b03555826d47182e9d9bf9df9cb387198a00f33fc9d1f4f92029134a2f7e75a68dd3f83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a20a0f0b004fc13ff94595411851645be2d317d1486810ded90ab49a4c1c47314c69d871c924a6596a55446eb4be57b2eb507c091958a38a7ec989fbcf646fdd404cd73d0205c80115f8c221281358deb86faf4f99205a53757500629050237c10aa4b794832cdc158f6817e37eef67e20756e8dfbddca1054a69d3f0f97ad1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b388d1ca4f50e69ed31830602a25ed9d755bdd68b2b6477a7d9bacb2fd46a73e552fe7a3583241e6df70005be559e43735eba67c257ea5ea5f6b701d5a859efc507dbc7e63861a26d4d423d0bbd8a20b6356469fc92501fb8d84d420eb62beba4dfaa55588e8b90b9ae80f1b7aba43135d71eebfe417e646afe9aff593156c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h469a0d52ea2069ca989384727d918908cb6e9349d0b8161da405bebe64636302cbe93a6d218395a1c06bfb8b0b9df0aa78cb9a6d046bcfd59b040bb423171a7e52dcb19113360d50b122c1904c67e3dcfe98c900cb164819630fcc67a66946e5bf7b29c8b7d1f10c7455b530cd16894909b8c398506f5988d1ac5af354c47f89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc837f90554269ba29fe9c75257e311f4861058d955b444c34c9287582e6d05b36187c4b8f2b46510df1cfe8f31ab69f874881df6fdff5004aec54d31987dd4461cef9a4fbd36b152be8e44aada98866f754a277db71c03e1be2b4ce6310e80f4b11abb16c55c6125fc91a25a6c8f1abb6e3290e13bfe3ac528317626280ff494;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc4a793d0165b39ae0ae728da036867e2cbf4ff64a8fc6eeaa587078ece9c539ce8d28aed57b4e6ff868c6e1292bec028730128c1d874659856561144fa2f788ec9082b7693bf88062ea6b802b04b407d16b1e740c6291f46cebe09f928aaf6ffa96aee68bfb5bf1139afb05cdcdb93635a0c41f276592e8aec5c16f47626d02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h889f51efc3958e6849dfc1d065ddc3076b906abd69b0d064e11691a3e51af6042f89e6de948b348fd3bce720d2429edf90b716e18e33d6664d58b2773406bf000136be93c2c9916b90f405f53994e2bdd96dbda3efd147734f8a546be5f51a8ad6f6b60861d9e416f3d1df50224f214228d2c4b715834914e96f6327b8bc502e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f3f3aff6d74e82e9a77a1f6c8e06966433104c0921bdb40e0fcd619d8f08d03f929a3eb204c4f57304c8e2b3225a199ba82e127935d24dff8ae409fd70f1f48a8863b504080fba3d606f5574b2df731752566c931da3152549e25020cec1ad383f07c3827691dbe974396fed4a5391eb337a5be91344c6700df0de9748bfc41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf99af8ad855f89c1cd5204c71798a61a038761fa4db5e4c573739cc9f07b21fdc35cbfe6308f6e11f50b324713a8b4de9ca441d4c85b9cbb535bd14c0c98416501f18173fd996534919c6297cd649a092a586294ea0c9c4ed208335ef146b097d2a336d7daf8395d2dca8cdde77b3126289ab2ad6aca5d5c10943b6e0889fb1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16d27bf7b119fe39a1d4292170b6c32bff62dca07bda9c7eca58aefff121b2fc7c7f3fa3209081cf86821c4e073df559100c924bd6ef2554e656c58935988a03db88039919863b19bada910b517a7077fb76e09dd3b62e1846bbcfa3e6f1517734a5c8317b97aedad5931b8e9602aae269f3a65212b07a7417eba7c90f227bf8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ed44e9e6bdef85ba50f7e890c5cd57ee861730d3d32e4b89a7e86060aaec71c296eeef4c0ba7ad0201c02521b80bba40644c8822feb04d2c0c80c593c0dda957697aa3e75b8449b39aa70312f7096905a70522a56094aa5f4425518ad9c68d7c63e85027ce7bf5abced3a6ea841b059947090504c610de1cfc67fe3c172de44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb079460c51e57eaebf9d751ffea552df3fcc66feebb8918269d1963ae196945b2a908e80f308a24e8be2a521eaadd16292043c17959e8ac41a9416cb8a91f7007d34b33cc7333b488c606083e3ae50d2209be3b19d87e960e02c367c37977023452ac2a058116b3bf86786510c55a86f367ab0da884a623f8ef8aecec70311ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7ab8a81fb27a1147bf7af2d5222f7b0e947c13ec5ce330ee2395dd95546268adda0aa4dd87359aa23c0820979837a7c7a241ab79a682438753b408e6af912e5074781a517356b7575bca0b8c0075c44247eb675ac0ddf618f6e5219ecca1e9557a7c735f8c05efbea5f4681a2f024160aad670ce131fc559768cad66cd7de9e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce184cb55aa15681aa06e834a02d341931c9e38b4418fec6f39cb1c0d7384f66250bcc56fcabbe8c240b9f746393766c87c52946ce29ba35ba568c96248090cd754c8c8dddd970e891452efeea3e9c07861be2b12ea51cfb286f3cd7fc5ae15a5e0af9834a90f7a9f35159f26451dc97a394cb3acc76af64b9fd4e890fdadb4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86f137602b8f2cb2cbc9293cf3aada32cb1ee4694f61ea046ad185bd6cf6203dfbcf9342eee2b20e9e3cb7112534db8bad0730e4e53dc1520c25616f8ad5c4ee97b5749fe404f5f583227fb7b139d2a56e46d0a3d0ce3831247c668ee48c58621f11027387fc0125f67f4c20d6a7ed3f4dbf6240f69adc4e3bd2fe1d9156ad2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c778d5531392a9399a22950aacf785d09b44e9943ed84ce562cf3a7bc3c886bc7bcdc2abdf317b0c587996169121a43b73ab243a888bfa300e750f588b09176e4e250786f4cef13733310d0d61b9685de8ebaa82a5b798947ca3720f3deb641e371886c61608cb6f8db5e1e4e6c6c0c88192c0695e22107aea2d901f754276f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd768532214e54358a3d0711cda6b93d9ab616c975cabbf188203bf8d020ebb3178d0716c5dc7864242f29ddf577de1d376e31d8dec3a3d66e334bc875e6043c572919b90a8f85eef7f85346836d5995c30a13b30c406e105c15147333e2a29a7c95a220e0155498b6926cb59bed73afa7f33aa9f9e263f69f0ca03b95b6ea2c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96513bc309cc29bf7501b40bf673e3252ecbae3f8b4acfb4d7b4074a68a004be47eb5cfa4c189d2fac9eb8bb488306b3882b04eee7b848e2289c1fc057a91b265d4e056efe3f024368cdd5d85a01110f0d73a808f57d167f767d46c310d300f26eb9d616d8e7f3cc36e6376d882258becb5b159d2c04ea49ceea2c2d3d2987e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4acc66e67d6c89b7adfe9291d288ce1decad44e5cec9e5a0ee589ff11fefe8bfcdcb4a1fb510bc049d2176a87f2e4f49744df3efc2ddcad51bbc253851f46102cff39f3b6cf8adeac9bcad41f200e73270f9db6d30cf043bf30863df284c94b3c02a66e240aaf8435d6fd8890bc2b70368d79b3717947789515f73a2fda8d4e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6a2773f5fd2471a198ad6aa389ef484a286faf13fe4b87d8121447852ad44c6f03f8a5e56dfc11f05fe0d3906cec61af00a65e37c9894d96630c6da3a702abf1238cba125ffd0f137f34fbbbf15f1027f0b54ead6f7076b4e2b8c152e3d0bc4977634bea928689d2333cc4e946d7a916478b56947fd1aec90594c03d9c8ba72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha55b3d0c22ed7ae8ea6f0d127615006aa46e42ae0a5e84adb4d10018ffb879c1138d2ffc8f1e3d835af1cdf9f130eea6fae66fb22703dbf522eb8b2281be8e327a2503a9e9a7286b4816fd7102f3d6be6db13d65f551982c069f951ab3507648b6ee0b2bc9a987712e9ddb4fe2c3f2006afc57d18bc71e6df4e5367f1d7b60e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7b9bb45fabbcd29cfaa9e2616aca29289e6873b5b7fbbfcd1a01cb6b5e9a40221b2675e83dc22c4c367fc7592c8c1bb87f3ec3a248af84c9f6dc6a577decca8374ce70a3f131c82e4b6487b43a07eec1fffd1e67fd744dbe90542c7cc2ff22e0d557a5e21a412ca246c96b039bfb1e090fb0415d3701dc94439c12b20e86213;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56306eb66d0d660e9be541cb5cfe6edef1ad8da5154538ce47fe8fe3eb3af131f63e41ee706151b2e6e1c13d0a804986e1a1f249426469c51780c63eabd46fa04bd15139da7cdf46d83fcb902dec7830c6475561c26c489a44b5aa9947e1d77f8d591ce2b21b4d033dafb1629c06422ca93d6fbe2048a023d64d18aedb0c611f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8ea4babaac513667d676aed213a01199785c203a159375f41e56c592c33cc334951913a43969b1ffee749ab6675d194bbdcbf747d96c4df9818737ca59a59c14d55452bb1d48e5b750f1cf52dc54af676a1daf467435b02c1f5ac584f9d4a425ade5aaa5381c4873874d9e30a268c98cab72ae97eafa89018cb793b79f8ba68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd32720382ddfd4e6d60fdc203172c3203c01c0c809f7c0bbd5ef720825231a215203b7c67b33fa1d41ae857448df7c379f073d1aab94b88708349eaac9cd58c10a0bb50ba2d9582dcfa0cf14b24939c79643a7867c753e0849fce1a4c70bffabfaf9fc428f941b6ffcb8f377e8ea3bd07fc847276df703aaff508cbf79596a1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73e75ce79fc8600f24ae5d26fdc2897d4786eadf3e7d540890c4fcabbf4817cce2d2e9b7cec4becadd63ef276d7429b3055ef55faf792c459d43614ed9dc88041202961e76401496531a2100bea93903348d69c0b58cd2a206ce2829ab06eaf8a7730ad4b6edded94dca8af59d1da9d9bea1e751998c3204cfc99db994d8acc4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e2f9b1ba9f820fecaa138b192f3838eece010f5507159183016c2298eef5026c156f363d057f5b4d1a973951ab0ab85386c9e8e5c690f8b28edf992d96d09cba04c0760a820d2fbc2ef2615832fa5b6c9572dec7f833432da62fcc3a1a64bfb6dba04de16540ac7b2fbd820f1574eba78912ce0a06db8fec862b9cd038d61fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd5f5cfd34911b341fdc953aac7d4dffc334c9b6df06ff5949eb270c3d2b8e426f63978708f48afc50cc90f544c64287acc4d2247e13a1a568300171799f63d6b6447d14e74f4904968ff7a27ba316f35c72d2967e888f62496f511ff757467dbfff41bcd2352956c0b367b09cf0e9788a4c7ac295ed6fcf2f9d63840911293;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c09b274e16fb887edec392e297d87ea75f0c5ce03b420188ace12f232defe0b709827643941dd1a89bef357d45b8df82f619865cc6577f59f108787cfb117a43710fc01ee6dcb6f5ec0600e9e33539f99886567df2d295dc8f51862746591221f1987d83c35c614a95ca425e7684c0963767f9fb3ede5d316f35fa6d0b8ed32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd51c1a5561294dc9d83c4bbdc0065a55f6d38224564ad8733d5ac34327b099a8ece79b06d8a9fde578d765cec300883b76178aa9eba815b17829b7918d88cfc94c3707e11dd8779c93cdd575db86b6e0f17cd120e9cb48c83f908c3e0a1e45649343655270f6e73bccadd0ef77a4225c1eae77de790be356d55dcc72f546411;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h698220844290706a8539b495e192d2fe2791fcfd8fdf5944fb7ce2eafb1fdb57efd6a4a4e58641fdcfe4f0393840c6aa000a648c842cacc9d990a591237b8a93e5d424a856438959dbda2fbc5593f553624410cd0344120350223fcda2b87bd0d3aaa5916c6bb8a1434fd4d1ac455f8fbcdf744996a2db29084c6c076f20c1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc13d835d3ffaf3ab1513d946f13f9f19a3800e3d490c31c613649aacca613e69f799418f77f4cdf2853489837ea82a7cc38558469d5c2d2dde966bdf84368aed3799c55cedc72fc0f622a5e5a94e65567ad4543132fe2553b4d08b22845e842b0309b9e0a3939dea36fb94b98680c1a66f6774babf57ad5a78c6622c7746bb5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9158da320bdb28a8533e793763de8e774c48add22635f4f86ed4b8ce45b9f8daa1ec10bb879a374a2c5269647c0f2461eba2dad99730faf8f1f969f922db54c563470722c76c6f80d88abf9f0dbd41d1d569a3363feef6d0dcd505eec55eab0e75b3118c31ed1b8b70857aed21fc5638d59309ede0c42ec0662e3b6d5074f31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha058bd1267dcce9f718b111fd82f4034f14eef2592b3e72b2af0371b6bba1a76815b380d46eb3f42bb90b1f0b43f1d04dad8e35ab87765672fa292bdfd09bb12dad5c66d876a832f5e086d4414de837e2489e479ca8dabd2dbfb9ee40d1c6bd800e03428bba84a86323f5aa837dbfe48aefe6fa930fcef06627f979cef9467d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fdc59e45da6fff64e86ca199908ea5568ac1cabd681b2de740d7351ac0297f81658bb6cb03a0f921fd2657c68e3c94f660032b8429da9535d7221d1883cc9e04cec4b8b980aa38cf84607ddeb9dc68978218b00786f15f2e2f48e847ed8508b3de4da3a0ff4896d569c07c46e18b0bedbb5c574598e016235306b0df599cc1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacd159170428712135014d2b62e4055ffa56bf6fcecc7dd996cddd886553e6112f8ec7e59b0f7533191664208ef383f69f93d9465e598218082d5575d71dcbfe08323b851976d49e359ed00e2588cc182eeedd36db82f1d2820c7b9d74ffe8620745bbe262f3527b65a3ed1d8966f33307ab52f989faba4ce09a393adcddae23;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea55a565b0c93bacdc719b54ef9c200b315f44353b6ffba2223543c5d664541dffd9a30ea4f53873795dc79659633f6dadb382e2c43c55491f05c80e6d078b78c162afe0acb64053f8ef0335f5ce80f5742a37ce80c9c340ebdf2bef368ab864cb6c2d375c4c2eaf0714fb35e45ff9ee52abde6c69a7738a4a67d4836a8a76a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha766089b083da0b2abda46eba60b0100d6281feb218c1592a56dc489abb16d61bf8dbcf3c276bad924fa4f0c69e0f2deb1c90ae0797d51afabb16cf8fa82dd69ac2a51e53e862d23681d9922eae4537231757d4ffe397f7a2c436483c6d7865b7c7b1f9d81868143af4ee84c2f0b7b6b330d1c0f22c802eed85c7fcdd54f250b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ca5385ce43500fc0c0934973a2bcf4ae294fba1d747eecd3c7e52068cf21da6c2bdd3f00b03792eba0d5cd651410f0b56e1de361850e4e140d6cb53df8d251d77d0742f37b7bfd9cf2fde029c6524b344f9b552184c1bc3ff85b85d8614813ae7f8c88bba5340bafd977cf2fb53156ff60523761bc7321bdbdf8b6b9c26d15a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h485a6e3b011c085a59b0082d644c0947c5d00a1b775290dea4d3158d902b638663bca6a96f5d2d2751eb1881895c974a964bc42b8fc33d68902ac47cc9397cde336a9c691764694dc5f73a3a9f85f8d89d0f66ada37721899aba85a8e153f59a2b6d235f6b2be440ac301b1e5a19f408713973ff01c3b01f723a726e4e9f1be6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf74dca7f95bc7b8259dbc920c529377eeba07a9fd3cf0ee233711d6c854aa83c6e7108b333e35d18efc3ba20997b9a4476d0abb02ad242e3e2ac87bbbef719f1d542ae0ef8596c7467f4feb9b296972b2a6088884550294f6e886613fe38435915bedaa2cf01e69cba6e823bf14c7ec98045250b146a47ca2c159c3cb7ac1fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h468e270792ce83e9808277bea1c74f91af87a7fc04e1d5459a7ed099e474e1566464384326b9cbb2b473a2fa4147b1292997915ef5438a42a2be6a728a7e080380189132122d367cad2d723bd45112492d5673aa3ec313d349e49f74deb6513b1867cf744dc5cd5ba4abb0881c461aeba9ef332311f7991471c95cb842b707f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84b040a5d0c4bb1baf193020499774dee00bbb862963b2ae73d31ae1084106f99b6cc1e4b97be9a937bd1bde7de6deca70ea55b365f5a15782f622fac83d32f49958994a4e2ffccc315c15fd83c92b5c820d130cb34233b251c68b5006089b7505858363d761b0732fabdc7e4b3fceb83a0143e30eff44e314c56b725c8be27f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had0e507eccae1465ad57eea506242591fd3fc857ad6fa8dd00ad5c302f1ea711651fbc5bdb9cedb3598ee1cfea71a08bd5c678003819df40716f4b38f37d8747c27547f6234dc8647b6b167dbd4d28d4849a57d14e07680a500804127bf5958670da300c14f249f0b29aba8825f4eeffbe9cb11506054759530c9a282ecc004;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h368549b604fea567b926e86e1f6e9983ce3c43e757769b9277d7bbda4ed4bd56ecd879a509cc4316b30b85c8625d76587f57af3681c1fed5ada47f8871072e80876f9c2130b161527589746ee5e0930b8c230e91855c7a9ad20b06f0f34a4d94b115aab4148f041d9f8217ef13441a45e8762a0147856712317748b22cf94dfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87e4c450ec223bccfde35085992fc4a3e2228ef5717960394dd7aefc275d7f879e452b1b70b7c6f43937ec44a150197a4fa1546e8281251cddc6a25ad9ef440ba79a09a9d40ea32b1b78a98d0fda0de8cc85556aebd85b014e0d66a66035da325ee2c65c21681b418ea7367b80b9ff1f6bd4e198bee3c99cc04b0dd3042aa544;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4eb9c90572acacf0d624a101a3d24554e4f5aa4e2e6f9140d738f0a2849d0235e4789a18a77f39a7f0fda5affc59d57b70c0aa295c191486c3297fd89387c976d1462cd6475f108ece6e05ef0519600b50cecb029e511cc94fce79b4ef83d91b0bcf2f03afcd9b30608efc955d47d0395254936d809b1b1a369d3e381e7002f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3cc4ca6f7a0744539e0401e8ad341055ee132146d53e06eb917797a03de9ed577f757b2b595cf58cccd40ee57d2e8b6197363e78f2b6507138b7d2580343a6277723cde7a41fd811df69fb06a8d62529fc1fd560d3e0147e309b962e7385e6a94b89e7ffbd49ce746bca8ad514206c9e21fa2cf7818d50f557da0b45a8d7d55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12b17fd852425d7fa3b44bc158b17e637fbd5a7d7693df04bf6c7b9697dea93db8070a68f5bfecb3a6bd2892bffc3d2792c40e6888a1b81d2bab2dd96b35c1b92af2d2070ad4c34bbe421a45e4b1abd03ddf1d0f5eeef2100dda861f13ec48cf8204097db7926851cb9fff780e0d47a693aa691a5a4d8010ff197204d68be17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65ec7d4b9dd520d7904b5ef86fcc536236e5d933d2a22ccd57d5339918a4ad8ee571322937b62e5ca295ba4b3656797877d5deeba9ce9854101de7805315c8490f231ca6a80d50d427f070ef99dad055ca6aa5662948fae8a9aca5692b3b89867719bb3d49f9ff85d3e64de1cfb29fa5faab6c39e4aec08c19438053a87f11cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7b8d7cfc1806cd30f97593c4febcfcf3375657b6491d80dff7378c8ab2b609818ac895b777de6984b75aee58c0aecaa69c73d0e150070878ae266e40743355be1c831e7a77c593ba68c66df39627506010183696a6fbfa446f0fdadda73477f0db7b3678309bcdce4d4463490fe4e5f8f7d77095ccdf7b55e7c5d55faa28af2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59616dc892d4555f3d0e1aa5441fd3bb34d46668e3a789662b007a8f3a15d8aaa28cfde92b378b8dc32aa7ff222c67986c72392f40260be319d8b951672c656923a98875c040cf27fab7c908f54678c6f28ddb115815ccaa85361507e16aca419a6334f4c0407910284befd1d08f0ff83151e4c04a3840ce254bb130e46096a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4272d28ff838ec6115c2c645ab94199c4301be8b075655051636c06638303ecce681d9cff046b3b2288a249ac0371ce9618a60ddf25cd70038fe4bbad77864afc3f72138851b59bbc3c6138d6ede886dd6b885b28d125fa8531358d30b7af5906036da590db33f0c19b7de9ca671e24d3ae7843e95b86800dac41db4317d9194;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h918edf1d635d23cd10123cf3fb95c476346b24ed854f73a1c210091ed3f364c8381ca10b91d09211860f6437de98992c754dc227157ee66ae26c32ad2ec38d7001c0a1f9d04c853a468d593f48a5247e519ed8b0e42b36a626ff2f812811086fac6119ddfb4e9ce66a200c2dea57a948e820267d30f95ee131b34e108a97992f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34d9dfb97f46d9a56a1fed6d55e7c182bb90ab5fbc8b1adbdc2cb1841a627ddbab9ca9b0a175baaf5371679572f0a6882de0a054f71b51562e102edb7c0a1ddfdb338205fb92ee823cb9aacfdbf8fb85ec078d818a3d50579980e4e6b8153dfba0ac1b19457e53efa45640c72697526092a86d71cb95eaf25faa9e7f46ff6af2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbfcd70f56a710945f160b49f7476d413d755559d1cd2ea40ffbeb3fcd0438ac22fee61aa8059664a0d58e5cbfe271fbd79c6a0f744d83ab4ad89c0069c1dc29d8fae30448fd949690f3bac75f412e72e97133c781ea84836c00a191a247b99af238d16ddbd6cb52f57180af40e689722149d26052d8fc954e50c082460614cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5a54a60c1375ce33e857e5afea3970874130d75fa52121d9f2529b66d5adc03e1ad057c2fd9618a31e66bcdfe4091e4ac3dba5e87bc673222cd99b60cf11604af1e3d134b7039d8fe945cc295d975285d9b33817891f94c6318f236aa2beaa1125c25c95b3be62d7d4ac7834851c66c50ecbcd96f173cbdfabd18d61247c5cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24cafe7e1a2d41bec703092afc7fea8ef501174a4f4e20e28eb13c9ebcd7f8f92a61e8b1e26ecafeb639da147cd767510614f9c29a867c9a60fa56ac5a4801cba00ffd2801d4656b67af575b532646cf249e58c0acfe90bdbcc7c9fe2170e07c0e5074129c3db34f5c2d8e00c00700a01812e7323c9a3dd5487f296549bab734;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e7805d9829ae4b2e7aa6e1f28ece328fdd9b44ad7250ce85bcc4b1cc88c0035e49056a0ff8a9d5be3f75495ac53691c7437292e2d5a63e357a0c02c020c9bcb410475cf4ec24bb0ab898ed07de207a816c7ae9f5014a3dade0081d9f1863ac977dbc57e75cd816a797e68beb588ae56d52b43d35bf4f8355b193707501a809b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc485fe86b8378f3e21341979e009e7e990ba1579f05589a61d5f5b6d189caebd1acd219cf0b8838a3e6cfe425c6809b0dbf8e6747dfbb39c967dcd8536142d7ec72e3ad39bb6fd8e3dcceb51047132172025cc6e155038cc7bd5f7e2b64745894e11d330e26a2bfc28ce2d5727a2582084a8b96a2ad52218aef88fd0fc98b06f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c994dc82f307fc61f7cd70a1c0e60046fda347f0a136de38afa2377a654e372915da176fcccc0ae6393078c18e0ac0626bc8709e46c6e5b2d4faedfce0c2191d8e41e8c9b71dc215d6270ba21a4870fbf15806fabf2034f45d53ff780eff7dfc1c3b5576db9f494ac1608d6ed6e1cc50ec98e23c4dea076272cea0af6ef9764;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a822801c236afda26b29df7ecf4cb129bfcba0e189c2c416feb69dd5d8d962a249f04a4bd4623fe47400d8938c54460f77ab45b1b8af6bd2577a002494dc947467f5d545e331b427a659cbeba860e904b4d601affd0efedc83526f7f742ede4d7dd4aa268f1aaaca5b32f274e289ab25bc99b13cfedc3472f31087c97f99282;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c24fa2a4a9b52082b625a292f49de874ffd7c40dd7b7971bc1227c1dcd042d4b84bd7c29971fd0b34edb67ee5955c6e6d1aec9d8f029000105520f7c4f4e90ea26725b4a8e058146b54089c6e650da982083813446480f62870b50e9cbd69546c4276e2387945983049b309dc251793851701eab004f986b3a80f5551ac842b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4840f7821816c0a86744b76e5780ef5e12052e4e08866988a0403de7b44d070eeedd8b5e0ef2c834c7d9eb95f7bbf7a32baae0c4e4f905c2a4f04fd84b90a582e65e8ed5532f4c49e027a26e219ec8892a6075be85cc514d02aba44dccfaac0ee1175b556f08a7483d048d2a819a3831ca3fcebe56ea3795bc2c9edf251eb3ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c714a3eecff6656878c7993a849a46e8b07367e365eebf8285b304d0cd8328526e3be3804f615dc89c58d83cf6dedbc4c16d1e70a3e12aa4a76befc0422761f36cfcdf0e9fc0d6814a90a73dc7b48ebae4195bcf5060ba74ccca5406e0598dbd36879c34b39df92f82d9a19561d251b360d73a5967c9a5deb5386dffac9387d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d608cf40c0c800cf0eba58535c32d175bb0455a2b5dcc4280450c508b270b346a7278ba1fdcf605d2ecffcd8696bc25ef5bda49191bad7312be559d7d957b09049dd720b820a392a32edd42dd4a5d4fca542cfd167bcec87d81e8ff4e755b5ea14bf7b974da91ed6a21c4f63ec7ed0af3b38938b8f904c42a8adef30f070696;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1cdf30df6f0634d88e7b9fabf1b246c2cd39727e017efd7d3462ca2c85d02e48cc68f4240ee7916bfe6c73f2bf5c96cb6696e09c9f7e48971421315a4423583125aa4a500b05aacbe312f16ece235bfcbc86ee308ecd9a469782c498863072ec5c0707a2ec0f2d335e18683ecdf148df43de2d434164f1369010230036ae88e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda5b410f3089bc944ca7586a1f9e7d8e21f67918a49111c5f5c2378b70bb6a872e7c497130bc135d97fa35664d5deee0b1f2b9e3688d8c4a2b6fcfbd73099ac719b6135b24c548dbbbefbce6e084509d77088732526f996b2d284a67a5c4a7ec02c54d7be14cff36a4bf49c624cd44284569141880daea21c113dda71c4ac0a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa06575ddcde270271dcda660dfcbaafa452f2d654634a9ea5507de7963bc209d6bb5c465aad41cfeabda420c3ad298f465f5b3cd8ee311e5a94f61cc00edf051c9f3ef6cf540a63374fac83056d12ee832663e0177b327b1c839b72020011f5636ef7171c34f9839ed4d85bcd9d0fbe918222e872c2a1c68fbbbb0676d13226;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc47822a6ff07fe5499963b0e0a282d9831c072c6a24574fab5f3d41011bbcf7f0f872345ede46fa4521ed93b552c4a96a40a8e61f694c7adfb324e7e2801ec30356c2df5224209e25e1c070714097020c54524aa1a44b393a7f85e8ee049052535a6c2bc6e6bf727b325295e288dfaee47dc2cf605e2c581c38c51ed9255754b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h115f12dde343d7e75635e505e1d12580c9b4b08e613385b921d16849dcf59897668ce2465190647f405501fdc10efac3ab55bc9c6b1bf838135fd444b3450f398dae0b1db9fe748686d4db6634a759947753f6d8226e9e36f52f50c881cfe4ba3c296413e4dface984f163f22036581c78bad8071c571fd637d8eece7f1cfaf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d14f348acb5ee6284d6281a67c6d70bbe741a81b921d7501638aaf25ce198b70af494feedd96550a48014f555b6ecbe29a8236d331376b17f50257ae08ade4940719b7cf09258950543f38961e79f7050f5a8e99320733714f4589062d8482f2e6c90737cd3289163e526009d2fe660e7a607891b1b934bc55d63d0b6378296;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7eca99490a366108dc288a90066eb0a27029fcaa1ead0731b3edcd3285b507a563e26ad398d24a1edf90f292f34e13b1ac1730ab4d1a4093218981a5c4c6a9c00e1ccf4ac5269af272af727e50772650be4d12805c3af9d055558404170749bfe588b79bf3839a2531b5ed85974760a2ead996fc4fd7a222f6bff01f95091b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9a4d082261cc133778ebf3c747a31ae1e1c0276359da6e4677b5e2a6fa7642493360b95f72bc97c752166562c15a513007635c424888d724007dd05b452a6af97bb2b533e4083afbf635518e9a0de6b093cfc890b378f7e62fcfcccf298c53a39266da12a685f4eb264905ab392124bbeb115f145bd83175d40be7b679fd0c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff8ed6dab023f5ae24f684044ac0cc3cdfa01c3a4021fc8237721825efdafc3cdad233c83ef5d8bf1dbd1bf64c6a3de0df6577fca4d49e571a766945d244fdabfc0925f3530a02271e496c38f306942bdd29cfddb65d0925209e0118eb2d8cccf850030e33836df7423d1af55ca946ce8f04df5dc3ebc3c3718b8825eb9a02f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d3d344914fd7bfe2597b330438d5e9038082a48c944c59ebd9ec5f499a36e0d967c7bcf89bf2fc95de78d4a0316796f3c727688a16be787ce8e716ec7e7256c5bcebb9d3564b74e31d7553ab5f4f0fbac1c6d3b7792ddda6ce40beb80b5841d831814fc5dbc689b2af5e93f718e68c52adce2e9374fb474c4a8701aa0017412;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5657d18e416add7dd509c1211beecff76328e4eb7da737ce6d148f98150fe0d22517fc0ef602dd9a6ad3d864d3b84ccb0afa213df74947f5d9d8fd270fc834b9fef4b38fa9f5218beba96346395bf538e88d1fd18d61a28607fc93b4eedaf12bf5c04587e5d3212a9b889d50e0a90fd018fba5ac87e41af06cf895e58c774e3d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1716387f0359775dd53520d5d2c36c763f64601e0f9e17d2059992fa8c9c53ea192b0ec7f02c51073cb10546ad4294e98bc6f84214562cc93d1033e7e66567a46769b6e71002b8854c8e3c1a917853e07975325fb2342ceed1347e110f9f629108196f507c981e4d198700f79a3c96a648e30f86ce5d1dfc1dab69831d079b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71c9962ebe8459ce016f0b4083349f697a4caa830f6b7877f2dc27082fcab33cb3c92801d1101f0fe62742694e32c68640a178d255422db96615de1ee700aa437d56c9598e9d132a06df7845c40c055a1f31536ca7634f65934f2b85d15d68d920450066815f61700174c7e068d8f88b94765d5230b3b53f03d73069d2ef8fe6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bc6086307688110779877561c08f482713f266b54074c43c159f62d08d2cf7e77162c54dd3ef29f1ad3d52614c094cab180fc27668ec8a02eb48a79118a289dfd95183a44444c1239d9c09b710762879d8e126a4f46d57d8dbf48419a35c73edcb75df1d171cd1d085faee2f2dd10cfab5ec208285f23c7ea1956ae1848e818;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5305e531b61c8d57d24c74e0a8bc567b0cacc8618e3af295854994469ed582f66b6af2aaf2b13c27c04810c8186f1faa16bddfe041ebaf904ad1a7633395ddcb1a35a94bce09985689effeb7ae43affa502ab9102006103f9a895b44f406cae3a470777fdeb643f9d90bd0de9391bccdebf4e1fdb4a8c47dead0f020d36c371;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a35b27f99c8c054c72da6e1b31138787f92b5c084e234c01c2e2f52eed106463024507b3d67da615be093be772befd0509a003290d5097262059d0d9afa5ccf7f6d080ccbfb96b4a80882424c4942ecc1ab606c67bde0ede1a674bfc1259cdb9228200d073fc40f0912cc08819e251b01b10a66f04cd01987e25128b346ab28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6201eff19b18dc589d19af9af2f86a15a46a79e6b61d123b5d8d332cb687134aaf291138a78f2e9b74a6a9150a1df638cf2bd0188d0516abb8f2a2c92cde0032002b1bdb65783be9ea393aff8632a8bd63d8054b08a5e75f930b3832df6cf7a140e5e42d6d6c3bf03f1a0cfeb8047ff9ca0c4d6becc8515acce54dde36128764;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he63b632ed03db2f811471ba924bd44cb2f3a4bbf717da96d1a522e32b2354b02cd3cd7d42fa8572d00c873f4b5b54ace7a31c7b8aaaafd84a8c161173ecfe278015e4530702e9f49f444149f05650f701212b4595f9edc7bf7e35ecdac3108395af9d1016cc3799e5f1611f3ac50470f0a4262efa528bf340868bddf09cd2626;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc03cd5e9e93e84393e922d9de3ed1b0d044e03928d282990127e57a33819ad634957f8ce4cb1817013371338c973b4e36b7fbeb860122892f4e941b904204ff4f120aabe5b93566ccb93b9a5037e38824ae15221ef7c96d53cef58d43b03d677e8f21af74430335d146f7cb6640d603bd82404b47efbb79bc72d305767c96459;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70acfb6428bee3a5be35fb3eb6af7da7a34da00c9b215bd978be98a4d98b3988010573be71a2ecb8229ae28b6fa244d0f7eef0bd344db7ddc4a21018c43292258b037a755293468ef793e95101a85ddca934845df6152e9b14404d924c233f1e615ed87a374c4633e9cc58a1f1fdf7568e02a4bc58b3e2df705bf80bd3dcda2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c7bee3411f45012e36c43b5170ea21776ec1754e339ad36bdb67d560f61fc9e2dda165d3c2ddfb876d1d3b3f5493bbee1a686718e20360279f103fc55a25ec6d40d7fe5dd7ac00f4588a2abd507348364bd0f7f9bcc26e6d81dc92653c1cc339a17c370f6e686243f604c826dce5a7953b6fb68812a4b4f1dec74395c235e1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc58b6839a44fc28458b9403b7e8a3867f9f02aa4cdb4de8239b78983c7a46c6828b116373f5107cbfc5725986f40950605a7472d46a81630fe118cb6eb0d78d4e5ab7fe32cba687e49643012857d7fbf6161e18337da0742656fb4ab523313843a8877d53229e83ea7ecdab1795efa67cb2a9e20bbca371a098f920cd1b226e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c2898a6125d90935b0a7d7e3d51c4fed73db3a3edb8fdf7f19c5b65177e6b09159e79dc7c1003c33c78df1f9069b628a3d3573e1c5d2b5ccbd9ef152325b7a4a18b3e1e605aa02e58c250c35d2b0dd311eada6cffacf2dfd680b151e50db6258eaf2e582cd179fd238d74e0ad522feeb9d1fa934ff64adeca4aef3d2c0ba350;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc1a872f4303c47bc9a6140928e3c0165c127a67a72de8b2e708a36ff899c0db70eb34b1a6d6d6189639840c88919dbc951125dd9651d6b988ae163bc2b8b875ec606ae6df1704e3579b0cf1e31e42f21f67d95d6c5b3b4fa1d415956d266c2ecd7a7fafcb905065fb884be3aa824d14fa495c6d261fc5ae8c7ab3b61ad4c705;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb231c4e83f13ba33c7ff30f20ccf0d965f064e5d0f23fc7f8a771b370ea9c02e67839cad642dc333a3710f01dfb943b01eb003fd55e5a181d97c0c4c3bc9b5375cf0b4a6ef9268d91ef0db2ceb86b918d1fa4cb6b7ab412a3fe729dd558206b9e4153153a2b4e1e2099801da46084e613b65f815756385623c60d834427846f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf2be7ab9b14dae2f75672eb31ab1853a3836a20bb73004f5ce1b625b2c5d102a9fe037c96aef7b346e38431a61664a6a1c29fa5f414aac9d521cce632dc7e6b39cf8235504520b887bce74ded2be96f20e2f423ce66749d53fe337a9d8bdf74302e63639e2d5869c981b2dc1257409ce37740bae5c99e0b13a6eb56e7eb8de1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3931917a4bb89c69c2cc39b0f787e2006920ad637cee98cc7c19841f09f1df29a8f14f5cef03ae63b51d4a99be703e0acae0604776928ca596cfd731cf2b94e686d3d68e62894059efb4916aca277d1d08b0791b16f9fcb10035711fcabc2e9bf3740ca91f6e7041e6dfe11383f181e45bf7ecaa1d83d944a3f1831e1d7004d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haaeda4c78a8ca4d62563b2c8e3d4fa182490c87ae56a7b07ad0b7651eee282bfd370e128b1ecab020581b445632dc5bf149cba288ae43dc3f8683ca785ee2beaf1fff8ac9ec9bcf3ed9abed0fab1594b32ad3ec4dfa0ad78cbe31dbedecbcd95303ce88e44266b5b0683f4f1c46ea40bb239205bf646fdefa1c596857e181ecb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4880ae94c18dcea81b0bfc5a49da6b669113a00328afa5f2145804b493f8c56b4bbd3181add957c9233f3a030386aa3d020b942508bc2a2def2136aa1fe39ec9a4f4497737189c3682f5fe6693c71e850b8adc66793017020027531579a2f54a6038e4d29c72c9827100977cdab98c1d6d89c6a071a5458a7fdd54b9e8cd23a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcb6adf28fc51488a6ed8c582f26e1aad0c0fe41cbda04b87d990c9473eea5ce1bd7c398e020df70f934942dcb79adec285cee2ee1ebcd34b8b9d9db00a7d9feb59e15c980fb1c9268c88bf490af47fa3717b388d9e6e308906f3143c75a6ff5cdcfe0ca727cc72584f9a793c465810ceb7a9f8e689b05f9fe9a58c3a61f4b92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18ff3724e2d2621328fdc2c743c66b4faec1771fa0009b1f8ac1a217cbf5bca0748f0ae681d9a7bcb149557714548ae3002f8141d5b2d8af7fcdd604e87aa5712f4ca8b9b996a4797831cead10c0f6158e089802ea3998e98d374441814659806dd9b7eded9cadbdc62ff54a0e1902e4d7a1f555030adb35541e4ce9529fb7fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb38085f922e8cd0a509fdd7fa6044c16af7c5d117d20f07caa0d59757a33379ef998e8f6998e910a0e4c4ce5811e226ff1aedf238d7363bbf75dd3e32e32b2c23d7ffc1c1f6177b593038f74d8461ba5e0f900f153c2292e3e66e8fd5f37eef84aeb59f747390e49f9b51d23bfeaa21cab393590ef30c71557fec03bb6e01eb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h693bebdea34ee81beccacb144ceca2e559af5792599eea43cb8f7fa673739a504dd7cdd2741be1f5366524e91b3fb3a483c1cebbf4172a5939ee61d0fcca8d7b606192c5d285b8d076eb8082bc4480da6ee8fae522636fdd9ff6b82838da53e7690ddc6aae283872ca872bae77f7b67cc9ae07dcfb4746b27e3066c79050e8b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaac644443e06e013febb9475e0fe8fc02c599fcb1fe2aa2fcce9c410ad03e76e842636e8fc9fee7146724355cd39e448e8ea8a85e6e0a2648891444bbabcc4db36e34ec9692fa3787c9ceb30cd147ac39008cb27ee32643d932c1cec33089b06c116f6a74540cbe61ee530dd0733190d68df8bae454aadaf5e0079c85cc7f14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h299d38ead65380040e8e3c7074c6cee2417593513451db4c5417189a15e395a4bf079534ecbcdba19e18027974e5d9f899499ffc1e049fa054560b38e81a85f7a781e25c2dd217f9122aa675a8f872b6b7b3e3d8e807db39c3c662cb3ae3cd31d8c8541f108f2dc0901afe272496deac1250b19796e560a84490b61b9ff1166b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfed42791bfe06c4d4066207a306527a6f04362172af8bb0b2b6b694af3ae905be592a468bc14d5d1ec2ff3b504720845d6568f669f08b83080374bdfafec5858d3a16e60e93fb57ff35c531f78983c5e26d65e58818e92a8aea211a66efa36b8ce84de1da56e61b273f11d1977f54ccfe1f4353c35ce45ec5c51069fa541750;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20ac94ee37e50173c12202d42b8e008502a294580e1fd6ee5aeb1969260893057e24d83ff0f81435ad006977050f948af9992c26a1bc12394abc1b18d22df6c99f353db67bb5cdcb2a178b9a72bc956ed87b24949a24465297281efd34ed13ec2ab2d1033b890a4f22a839581ca1ba7b6d0f247fb3095340c9d95f70530c8f87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f1a558723c165c3b3c6a7e14c1d5932b310817cf081c48cc9fcc31fa8589b6dc55c13ea13a50546db154ab7ba939a39e7b5d1d20098b3b23621ceb1b098b9cb81b06d657dcb91de704104e4a75641f2e8d9b91ab241408f4137e05ca4c679ddac9c3788d5d422e0c97546ca6b8b36744e13062503e2c6022115f2bdcaf65a5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdefc165eb3b51f91488c555560a7fea1a2b1510498548d7304c3ec3e28198f14f5f43f532c81bb4617d3c8e636c27620823abda9b30d8021e6b8bec725c8f7a5a7ac5329c856b43d39d237b2e5961fd4dfa8991da51f9a858a8c7beaca82c372a9f5c0bd4e715beeac492bf04cd0e164be48cf19f85b498857f6c34504169ed0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1cca283cc350b7c6469f3f996f7963a4f85dbbafd3f84d6dd2820340c198bc4181b5cef1a107aeaf311857440c0c7e73df7be87608c2fd3d5f7c58faa2bddddc14c3fb6600aafbf2edc016fb1f819494c71cbcf3b44eccbc7b899e1b6bf1f6a066f574dad5e3a27f7b4e0a7b7bd2172c3dad5d54cb72f04a847f14b45bd822e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1002faff8d8dea369d370520f46473d95abb0b34b19e3da24b9d76174ae34789e213299042269653c81f9cacbb25a311494376f68f4ae8e120d722d5dea12d076ee0aa5d39a759fad03f31ca43f0e4e42b32c6abf9993b8fb60d23db5433c7afbb2f7937aa9b5a6a43cfc306a78f8a49b6237bcfcac3248351adb03678c764c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h997e70cd40ffaba4902c1b765a73d3140b7671d3bff334b1cc8eda97cc1f02ff8f4b8326d3f24c02ae3ce481b0945f4f06e52a6f444c33fe7d34aa22d7077aae1d4a93ed2e147febb9fa443f7b27110df6b3c6db300a45fff48d655260bcab54b2325cef62db3a917b7678da4b97f4d7653eec2e4d83974ce9949f147e35f0d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fbdb89af994287cae5025063f32027e17d58f71fea0733d8002a72f8da0d65651cdf31428f339532e5c20e447afb2833b1dafe560756abbda33b5d6212b119c7fe90befbadf8e00a2878bff3dd826d7ecc7f82e69ecf0fb14ccae9540b3e9dc786397b5786d60334898da41ede5adda4f9be1a015490e20ef9423cee8025dea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3db831ef392e75bd0a0e2c70161332bd94e3a20f26c2ce0f212e0604f4ea70cf7c59f17650d66bf457befd26e3c8a684264f27251017c863fa206a07e1c2f698a94839592ef4f88fc05ac4232e765c0468b39c01e968d69cc110c7f50bddb7e0df74b50ce0b010ed04d1eb5022b024de9b68893d4c6d54eb24004ec32fd04dc4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6bd2055bd509bd125d389bf87759920fff3c3220913180d151fbfcb2ebfe58b96a51939265a8bfd9c80e1a37e32d844ae0c44ab7893f552be8bff57c16b5990ad0bd2a2207f6656fa7e433d64812b27f030ee6924c8ca7f6e5201ad3d405ee780fb391701d452a11c30eb5b0f0e8140f00269c30a613f68aaccefb293e3a506;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc1e17dcc7bd1d3ad698af72abf8be874294341b96a6c02104e549575086be351b0375aad4aa5eeb517811f256ae313fd103d3bcf9fd46339da4f547a034ef961a8a9413ea6031ddaf63b7268e20083aad5a3d2ec3af5288e8aaff91f74f3f18b753128cf731c1fad7c8527adf45d953692d6e1a11793d556d009473c7fc4e1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ae6e8e1dc2d9b2a83fbbe680c99c4bc56ec8700c2c6843aff61012dae72664e6ae853684fb0ddf775d70138e9472fd499574ff6ec418af92f77b323f45091706850e81d008acb4c6d97f69ff04a60cbe998e81d2efd44ceb07a226c18d0c16a8d6185f05df21807b32d7dbb6a76b8904d88b1df97839c04f82632cc27ad5c12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc94040f3e158ed5f042c381736aa7d5f0979a12642f1aff45515458d945714212d995885dc83fcac8bb49ba5048acade2e753823c6f78fcfbba9642a7b980c1140a119cd59c334e75ed3ad86a0798c5d7af40057a2e845d505d74d6a011148c56ab70372b4a8bdc4795cb502f0c75006211b9abe0ed693cd1a8d5436ba73ba8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8cfd221b81a8f4d945a47b69332f936637856a02034541891e0cc26824eb1c1cb5e05949dc67a71e4a79a08c25e0cfc19a1d6a23f143646645eeff124e83cfbd4cefbff0b30406463b4c17004cd2e0e0e9f44239417f0c4f295e32c05e1b83c675be63aa0bc3bf546ec9aed3b107372b4bfd1e2c5b7197a1c67de0a94b558dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5acf4431aa49480ff2399c67adae26707a718276a7b9a543f5fe4a1ab1d5f546fa38cadda9288307433c0e9e4dd84d83672b0addf36ea5e493e6918df404f2f7692459c88618eb7b249b1ff13d5393ed5207d88227e814218fac5b30ea816649d63cdb5eeeeef91c810d903f39b18485ab898b51a685546629f78699af23930d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72173f888aabf6570950b823337aa0ab70f6b1bd36cab5a1491d384f1a6e03c2528d120feb4d4d8a9854e667c23008d2c421347829595839295a228ac55d451b8155c075995851c74312b666b9de4fee0f84ea5100041fc65e10e679ad0d905ec2085cb80ad467e3436f6ab8334cea12ab631be837e8588cfb12ea3d0a5c7b40;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86d83485f07ecfe2a480739b9cfc6337ff143b2b605399bd2569b763e1fda4a086fbb7ad5a85e69d76c1add94bc5c406bed13983dff18d098caf3554bf135d131fc3d89ee505a9798a3d4d68dbb88145b79f75177e6b3288021eaf194de2ff19e06345b4f1e201f46f5ad065018c2f02b890b76103d4e9afa807f7d3eae22a6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h720a934c8e13c8b044a6396a75c4d2b639327760dd7138669b3781730359a2b95a3a5001d2373ba19b3b68a5cbb0a1bda351439d1f9c4728c5eb0dccd38f35e31eb1070ab1bee67c1ba3125f0eb97062ce43ede73a22807b6c7ba8268d423831e0285df21d3d522814a6dfca79f904437248e0aefdeb29789c89b51fb0fd3fa0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47e5a728469666f0a75f127f29000e77cf7035e021c2931e65b6be9a14a63b27117278307764005418a102ac39f80df79c0407e1dd31c5188a10bd253a82e5fdfc49bc65e28c8d725d02ae124fb5c9d1369af0038fd770f9a85cf650c85b70ddeaf787daf837d10b37b7d6a78108414b054a08a09187b3a45f5f7c433c662522;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haaf2a032456ab682e737ba4b39ad54ffff30d54c459ff8e05871820df75e5def4187e01092c3923579f2c5ae5e2926550a36b6dfa21ef418be93fdfce7d4e1a47d800d245926f81775fa9ffa2a86b80a8f0ca7ab0ab8a76bdf0933808ccde51c9446b128fe970e4c8a006c4a0da85c1d1f1ef2f9771a18a916ca3b2534ed2284;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11e2813592a5a0357da6941430502728726e9e2737d98a9123dfc2cd87ec83c15431d89330cc786f27af49c6235f00285901a2c4cdf2d5b3e6d13d24f06cca56cd59d66e011e2841333dd5664cc963c083b95f9f29d7a74b209fc11082d70b188fe4721ac2a4d7520280dde7e1f9b1431719b2ea43750fc509661e42e9bee6f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h402503c46a31fa9f58da5400a66e6ca8d59d61f17d43956a4c1ebcb9a9c43b512d46a12cd880b810e0fcfd6813afcb43ab2931d469ae078dd6c6a8323661ae2f81204c78b2780b5531d115a81ed0e1ebb6ec4016c49c4ed954b8211d7f50c3e803ea4ae9653cc6aa69a6de3e4614efc0091e8e43436e6604253993c2917eba48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc5b04c56afa3e15bafdd109d28ca5fd05fd29514ffe853257e129364291213fc1a9cba09141c7b347d8ba6518a15b8a0ac13c62a910f88ec466a8596c1db3adab5d56d300fd417784d92b7c9f8b881078e3dec6d2f7cb4831fe5bbe4ebb783803c9c8322ae614ac91d671f8d8cf480859097861a4a665ea2328e9d6a103e0a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d7fa5c78ae0fc74df2bf58c88e947753ee7af7b9e6d543950e62af680c5b53edc18563389d50892f2ccb6c4724fc84553d9a676236eb36bdc6edec6fc9feb3e97154ff9521762bd085cf2a0284482333c5cc7760919808132fb7b8f560dc4b42c7d6cb6a9290c1e688af6ab3f6e9cb80e29bdbd9e0c721a9b6aab2515d03a20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf424d17408a69d26ec0449826251a29640107f5547b3f6f9dfedbc82612d6721dd148c1ba3a9cc43f63c647c4213dbcc9613d7e54682fd0e17954e23e7bf6bb5a531354106f1452321f0af248d4621ea07fd348d1b00e501ddef218617ef9d87bae231a62fe95bb9cbfb05a393d636a5320f242462414f96a0228bcce8d581d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h209464dccdc5dbbbb25482c4b506d9069c4c2ebfc6604a28de50553f482cadaa99b7a9ac51418a5d8f00824596cbff5ca56ca4104011d1b2420aa3de96ec7ede0c84e5069303d50c5c53584e9d8784380579d115b43a046d4029d4b690aaf7227cad905ddf7175edb66293017e1aa756f8f506145b43aa7ff71891fd830f5b0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4d3037879399f1aefbbb213e39946a879835f4d84b654e8738ec0b050a225519fefa29bc5d5a914c90c3f0f83f41fcb2a5aebc790acde2e758700a1c57017722b9329aaf81140c1bd774e86b6e280da2edbb932e4a0a353d482e5b397ba6eb4e5374cded462f936d825908d4fd9fa6fe04a6865263bc565c17e53ed3b6c8a13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2f5abcecb99be74d823a3fa52e803abff607a583e1e47712026b7ddc7d19c17a9bec3bf50ae599500f5797a63a4272019537e5f0992a781da7e9fdaf2f8b59862fffd4d83b4217ad87b70a07beda7ce826effe094dfa74812085a479714f6169f743e75c6bb4c79378f24f5c78a10e1cd3d733f20b9666fc94d9372a96b3914;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc90aa304728cca3bfcd768ad27bacc42595f74edaa40c730817fbee817bfc5f1bad253493d0678dc240a3aced0a43f155d03d3b0e611fe01a47cbe97f2af32aa3c00442b084502a019abe8cf8bb75e97ebccb76a5b81f0071cfc804dccf351e6ee86d8d9fa941d4ab0e38ed7f40dd366f785905b04adc0fe36bf6146ebe99979;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h858d2cfe169a37c447eaabd942c41ad8b216e6a0757ebf5a408ac44cd24c08195db30560f34da6191cd907c1efd602a94aa912a77a7fbeb4e946cb02e102d7029bc357aae527aa0c1b77e4d02d921c2ac05801c5137a21aa99ea08e1d1d9a28c1551d1bb8f0d1efde068ca2ed8d2d8993a7af67333aa780712a992f7528f5706;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4825add7e5b731be31b1188b5412527e99bf2a3d44bfb6e947488df7534760a26f9145b284ffc53164f2475fe379bfa9f243ff1ccba9f92a571bcffdeb6e63f029ba22b18f18cb0ca7812e56c005427280de88feb783ac77ec8f049987bc468a5b4ed24387c99f89d8ec87bf3e8eb60ff729a72880c9b9b618376882de1b28cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5a7c7477a5786d788785c7961f55a96dccfb0c9f310f3947ac511a4d8f733c0ff9425318c9e15bf19ceb9d5b451f8f894766158fede5ed841ee869dbebc1b29207841cf9ba09191069945c1f1e3a585f7b758a6bc6ed955e8a6bd2e89544c2e3754a30dc378ec8c57ce96c4e1c83fd97c683811bd487af46707491eb639b4dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd970b4f66fd2383ea0998a83914607b2ada6d9b87376a590f686772121f1c172a8b500e9c520421cab12f00da457bed8772d875471cc0a0a855f8c12cd34d5faeb5dc39af9c17acab6eefd46337ef89873c100fd52b030f5789b5cf92fd2502b2cc3b3da89bfd7b86813e347712ddaa345c8eb409b949df160204971b895f1f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a11087ece252c38cba6843be512953c64cccabca250366d4bf21e5ebb59813695758077379c8f02d47935f8137247866f1498b7dde1d45409baa1d755a164451de947ecb01d2f9e5c8af7ddbe1f72202f86ee393704ceae637d891f03450578e86a4792e020fc2542dd059b988742fc6a7b29b817aba7531ca84ee91b3495c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe4ec4cc460140c6897b4f4b3e9ff0fca2f29c1788faa06670a728ed5bcbb30dff56bf189735fe7d97e2e0af9e1c66c150a233377f67fb7a7d5b5ca22c414eb94a0b806d2ff24999db5f7c650f7b60210966361559685e0d8c6011c1f19259b91bd310d6d24f33c4c8ae92a6316cebf9053561a4e342581c144d9837b472b7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaccbe5bbb7b22feef339674234b5d40e4ee791d84cb4a3f568f55c7ec7141df5e56eadd3cbae609f07e44cbf0a42d20bc8a3738c4d57c30b6dc016d6042d9e4ea3a23abc6fc640ef677b508446840386cc270d4ea76c6b22c312b127f2b6a52372ec271ca699058f8522559edc7aa81a61b514c875b2e60d58d2648d9b07154;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90f501e4413ee15cccdfad5c01acda3fdb923068fb6b88bad754db878a4e7a9e5c79f950d69ce74811af140254a36d93e07d5d22056f53365e084fa45fead22c02ac9edca1b16257c12663ec4a5a3bff1b553fbf786521c8a43ec8969fe5dd8fac35cf426e964e01d20e1ad5e24ec72833ac4a082175921de38fe6abead74cd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1058112cf9bafc9bf3b9e1d0001a2a9f9817c554569a4f22c4444b71645a24616c07838727d54b82b98324bd892a1b84a693757f63af2da4ed21652ecfbe691ce9c8697e9f8b88f7d469b0fa24a57a3bab67c0e57f9d7fcbb8979f364dc4d1b8972ce10c60ae194e49e36f42569e7912ff94aff7488ac02a900fa4ed5a949f28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8c2ce87af41b51fa67ec244691c81a48692d9d68ded07deea0f34caf7060609458746795989d2059cb63fd64b77770eb6a5f9a3871074d3e7e0695f7f85ae5b8dd8710852398e1136929df2dd28d978060aa5c8314271dd5caf17c6a9f7d265ac41d53490392e78dcdd1397bea9fa0a3cdb3caa3d72e17f0a1c59dcd1e49c15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3e08c390241c645bb111a6d7b6a937a6fc1fdf9cac02095dc16ef211eb5a5642f62c70f605e576e9030c119c4db3e7a141a296e0809e3c73208680961f3d561b3d976899b96b3e471583ca89660b2c69add2dc232cbde1901c4d2e4c9da09ed70b1492734b9e36281bee8897fad59c47fef8995073471f0bec992ec712db9d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45fd93bb303d7eafe8d2048465e6c46f29f8d557f572e6779cad36f406e2bed5e3e150d411f89e4f2272be5d51e9d7a11130ef7864db170e674bd5a477b7e3d28ad2fcd83ca2e05040d9d4dcab96d3290e4b64b7b1968bdce5b425687d6ae34a3857f00847b42c2a9a390c4c5d42b02d564748dee4909108ef8f976870604d4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1ec9b2742be4ae1232988474abd63de623f7dff6c97cc760d427e1e0355ccdd6c91f747d5aebf3929fc6d86101d414e7b54e07841a131a42e5aef66303293a6e9841f6576fa41e4f3bce5fe07f74956e94d244bee6f97e035836560d46f199558bf9ce42faec872acebb6470901a4cf81e345dcce9b3a82dcba7447054f0c05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72dbf689d36786b3854d440b20959d123671f7bb593e672b6123007be34376b525f56a600a61797cfc29d891934104578776c6c97f677f1b7eb76ecbc16c8a9a47d3aa10ca99aab3171d2036f2a043dd1a61dd397e3c2dfdbaffa5a763b4b00619cdc5311df99506e76fb9beefa442784a337dc96dd879d673e60338f5c52f10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h359dec6bc97e1b83997262598a8ebe9ef9f4b9a8c292c4b063b2a148872907bcbd8fb8625f7f2f336a13293b36e0ccf44616bb678c0b6ea82c2632b8c56de4e6824d50dba6f56fc4d545784cfab2fa8268810e40979401e0b473705fe5ecb5cb0d5e9eaa53e99e12cb2c3f017cde524db82b4fe56624fe58d528af2d3af329b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6001a60fb9fe409a4a91ba8382d44e1d002144ab8b972eaefc156c0c20d86d46b210ee0b8cafbb7786644d92e6653bbca8477f06f3d472d3e81f0b369ac5ffe1f166138c64a50669c970934c917478c14b061f9a294edc6a389afa98a8ebb2ae0a997ff1e159f976d8a4edeb2ae1437e0ff46069094cef91d174ed0e253a3f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h536db9fa2170146aa519715e374a61e2832abda8bd58d0fc6a3b294738c009ab55d5802fb97af25491ee2f7203859e2e81e6d303cb049a0c3932beda4942386c20e3c1f467ea7b91ed6b19565442da3163c21221fbbd2aad0fe733d8857e848e1766db9ce591b7cc2917be0706e9818dc465fe817333b9915f36bf0cb0a0f7b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d2233d404b8205d40eeb3f4e303d3d6b03d8b5a9eafa7eb581a369b7d23f2113611f9fd5ce346a808a039edc9cef5765279ac226911eef367d51791c29a822cafc03ee775791cfc9594b4108bdcbad2d48d4e6f7b46d6058c05b71110ba146950dfd93edb724f8d96a5c2f50cf307582b9fe28ed1f4b14a846f428b153cd55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ad9b45f5e31f699815e91ee67b9905f3b28bba0aa9989ddf8559e95298999ec90b14e666bb7a529eb72dd634d66c8ef0bfae34d162e1ce93527be67531deef77db343d0535c0f079242bf837b3c3c11568d431a189917544c10e595e513bdd2b2f6ca7b650d3bb884ee97d738e1cdd6e0f74f680018c2b18491584499c21c3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb37cf1a395341132fe1df258faa634e9f182c4077c39ad3650a1a85ef46f25b6303948ab642b4ca142de89bb56d3d5eadd77bd397087ecf23bcced036d9d2ea43c723f2145ef397133fabbb383b1f2ffeeefae26f80e20b49146a903cb6478615ef8d3fb96c9c42f7b36898dc1cea0917b4a4b11c5275b3e04a67b6fa89b90c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd17e88ebacb5716acbc86659b1173d7e47acaf2f4494c413661b6322133cc59c01c56a1ce8d2d3e703ef509b02f3df2879926d99dc659ba4ad3645795db5ec769fd50b51c7320977bff26fb05a7a2bc9adc29047677cf269a849688cbf6a59469b22e82c27a1d602f16c38f68cf36656ab8ae20909ec1a48ba404d308e1890ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h457ed766d6f2b225b03329f4ce84e1eec11fc5c8cc1d648922603c9a16deca958059a22bdf9c9016db3baab6b86331151ebe258fce56718df92acb9b1952cfc57a7e6a3c19c91964a5361d84d56bee2063dca4102ec05665cb55a6cb072a2e9e7c32be0fae9ea9aaa0fb5a6f8ea457376cd4ab1326c26dedacf2f4dcddb4af6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30479ee462334e0132c8acb86301d2d944a09e7d05cd67c41ba512d4ac2162fc253dca15fe196676a79fb02286946e5aa698249ac2668eb792559714bc8cd8877c02de39c54d980059ea4e556950f55bc02f0c3a2535367788b4336faad9b4cbf14f4c141d36657489f8969852c52af563531feb001e0eb87b6cd57af8a243d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b1882aaecd25b58e4e22270857d89d35accfba76c76bad27e65216b15ec4e0a4fb6933d42d16418eb8102e50036458a515dbb6c8ffef001d1bd22ee7fa1d2b817a0e4193969672efe1d8be1a67a9ab607a4dccac727802925d72c3d69ca897b047e2f83dabdd0560e4355c8bde7b6e5de62d5fad223401a36c84285b128e1d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ed20c5bec35af0c9f50eb5d634827657f3a0810d0e95a4db2a6e857e449faec43940bd23d2512e782127ba1124e2db565735590833a03dfc3661654f4fa259efe0f6bb5a1285efd7c83a4897191f2a027b52eccac6a0ea16ac626b0856a56b5c07407f6709e7e46f291c9f35c795ac43538aca19dd580f4b4ae39cd976583c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91787a926f378867317e5eb974b0e92e4d58b973f594fad89067703a6ebe7fda5cc904248233d5f0768a88359f1185264ba01afa180b6a5b4d3b03e482cbeede61ef0993460332708d02b5c04950baa7fc35325dc831aef93760c92d6af336e7e24a797651f68515b8a2e0d253a1fde840d5179ebd06390223719581d094f6bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dff0e4ddfd2eed641294d1887128628f162ee253f537b73540e722bc4264f290e92b7c0688c7b1119c31a0083feb08e2a496f10c6d3ba75fa476b1c39df95b30571911dcbd77e2fc9c2574df47e42f88a29b0a71a575f93ec19550f0f328007bff98ff3f8ed001adbe3d4241b98b4c76d8370f8a01caa76be52d18b06702cba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ad60baee6cfa90649c57542439d56bfbf4e7bf29e02ab27e1cd946c01dc66aa4977f67a86a53c2de09fe1917c3f9d1d87ca8808dcaa274a6ee68a2bc8d1d2c2930e0afd0971ff8eea776ea627008e4dc1c2bd69d52c9eb28b619abc806617709a902c14fac4a6575e22b169cfee337040f6e6c9a65ed0ad9beead90bcd6e043;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha04ccf9ee6ecc0b049cddd12b2b83c0f0df5b8cf2a1a1958356087a063986840426d5e7849b374063bba4c147811593aed7027e96710b20c20d344e9308aebdcff9001cf90cdf8891cbb5930e2eba31b8adc3fc78581aa60132c6d44eaf5e2dfbd75d2d3774a0fa5a8c2cf81f6f93f8d8ad401b367d160635c6e18b129509eb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1836819b1ae7d8b6053cedd476d2a3e1e8f26e6ca0310c67bca7c9006cee84cce2d586c409608f416a0d52b2fcd66871acb3ac266ddc48f1ad55140ec5494ea739679c8adc0569c1aae5d201c4c82478d4af2f2394caac0111ff1803cadac1c1081e1b8d6a1d6d192b3d6474de1380966c9c504f195233af0c85204b30ff1cab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6e82eb011095f5534b8965ede7ee997311393466afce29df66c13c11855491241a5eb496ceef21b6681da6c16576c92af98a6c5390411690efa2592a33b8343dec0a1f74f1a174b4df3a622889193bf6a320d32bb924b6b8d782e1fd82ab917d73c93a1ce3b82eb7f6a752e8031742568595695dde570b6e1215f3c5334e902;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7062a11c7dfe46f4f2f83604b25c0842291dcfec4d952b02a82d9ed14999634baa0388ae4792335f28ee6e2aec92857f160fc840642b24b1f64d1ce14c659ff78357c04dbf1eefefbf6a35befd04a9c755df3836fca444b32247f042caca39c977b3117e82ac68866986bd196554e07ff80bf407d2c127d26d5ed26ea28ffaa8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2bac2fa0e824a72aef87c02956839b0d748bef313cb41338d2a89c4c3d2a60c02afbcb42e645825eca0c8528e439c9037ece0a0ab336bd7ad3b52470d97cc9775351c71e5ee69a4ced4896b6a6318117e3fe5d50c3f8a01a13da91d5003d5c51da07057ed39af5a6d50f1924b2a8f4ffdebc105c77f988b59e32afbcca6ae74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heeb15d334334289af1108b6cf65c682f097de4a19444761c715e56fa5516c4a80492887ccd1e4b4b4030e8e3d8af9f772c8ff0eddf9181766e6111892cb3e364a6acabc91fc0faaf7c661f0dbf520fb1caa2d5167c82b6ba881aac8640bf4880a65586bdc6c2bce4383e3fa19931d919841b556b5bcacc90ea67bcdb4d909f75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc285d0bfe544a098a71c38e64a3cf5ed4690866a243a2a0c409f2f4cf521e8481c33a6664135ec9db3faabb58f034b1264124db13ff8401de4ec4b59bb293946fd26a20f21b56479d04ea3e935c016979a3774490b9148e9fea367e07b4cd97fedb8e8c56c44041af7d037e1e3b9c4d18afd947f6eedee9a925226fade5d805f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e91c22ddafb0b95b6bc51ff2eda1bed36d969dccc12ed24c273a8891594824ca019a037077d58808d528a3711a09715dfea80c2e4e5f4353f5d98a97e49f222f52a33a16c505409edb482108f39ac9ee7962f8778116750a1d6132ee06ab85237be906ded8609caddb18bc501db0476d0d07070a32db9e63592f88b1006ac3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cbcc82a41dfc4afd3844b4bd50874d0c4d2fc8b39b9217b4b6eac172c4281d9b12e4227b415583c1b1badf63fbed298f0c365a49de926634a04c4100f89a86596f2752551d8cad7f109636645ea2761fc319655cf441209dfefbcf5a55212b2e226f153960dac59393d2b93f46fa3c9f7e54df2d0d7f683b8f8ebd08f6af287;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccd05814f3eaf1c9efc806b37e072555921045132fc0cb850482cf0317462709c46f29d18695ab82cdad39716346ca78bac4c58b579bd906fefcdfc0e64e26e50e802ccf421e8ffd42e67bbd23fc31bcf610af6684052a4e5ab4723d8394c78e37de7e64d0f81ade85d0e13abebafa7335b9c6aa37506b550733a8e477b2f66a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a70a99113a41428a1c6ace250cab98ceab11b93de772aaed29271b68efe515d1432c86d05011c827df6d94d494045d9348d825e491366baa0a80f2f1bad1234ceeb79ec09f1b0c168be03a32b5a4252abc73d801f63d1664cb3eccb0e2d05974d0bf43db19c90eabb2a9bdcaa98ab6848aa4efc682b1660f78bc5623426aaa7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21e392b4d2cb4784f502244e4e6359512c8d20125898fbf3a04229c2ae14b66607983f337eed12270964bfe36f6c14e83a8db68b3791568aba7aa6deec4c6f79381b8f73277bc451ab162d3bb6ffc4056361756a8c9777807ec03643102e5755f4b468088a116efa8791d3df2674b995643493544280ca56e34f693bcdc4ae87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h317a66d915a14f003711838aed6f5b5ccc6190e97fbe336b36b0f0845bbd424aec2e2f54c1561cf960431524d8c3fb823f45cc881ea168bb7a06bcdec2c6dfae9fc498dbd7013345f92cb1d3cf141983036bd120766980c3145f1edfd0224cc008075b90ebbc641fe326d17a44077cc80ad71b57da692dc010f0b36b0790b35f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4f3d3df46f6162486460764420f3cbab0851d3d4fcce33ab2d97c7c5f8fa9cef7cea432847e68d019f9c326e8545285b2ce01edfb0737e1087c3b1763f5b1f29b87ad34d702a179bf09c79c816ae276ce7a9b6751428d5578651ee3c92e6263048b9d6460bcd4f473e900b09f030d03e2eb00268efec87cc741d062890c1888;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d3fc5c18cd1af4936fc8cc54ecb782cb582aaa53e89ab208329c3778a13cafa5682d48e2c1d2f0c40615e8a72d4568954ca712dd1f2c69914204f74d54b18702d55fafbd7fd3dec16bf516d4305e8f535cae295eebd1adec4a81370a456e0c3fa1b3004f61ae830a4d00f5082fb5e57e8f66ff5fe3d33ab50e5dc48d4a36469;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha498b637d1388335e645ed1b3235eda2a279add05dc60842b49fc8bd28f79297985ba732be0167a6dc970d53cb46abad9d70c11e00c81033549fbed55dd373aa25cfd23387fd7dc58887b3117bba603a27345cf46c44be8a2f28180621b35e5cc18b6e799bab2b027b35df97b50ad2281893f1c8da4c77bbd7fec87879a49a74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccb424be462b77bf42ed72a3c1d1d8b5548e48a32a515d642017682e7c56d0909084eda4020ed7a3aa9f0eaab5fae42fb96e4c55a569244b18d5e65050d7e32572c9e6c863cd00d7e66bdc564df0210a4110560f459f6d3827ab5c124b6c84ba1c0c931e8a29ebc1419f84b4c9bed3e5cf892cb2500d17d26a9d9747718aec6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h304dfd77289bd931485b60d6258f06e654bcd71bfb780489a3360ea60673b59739afbd4a1b765c939304e0e34c2bab17c13a72251734ad2a8afb5ad41021e438794dc2192f9e9e91154fbfc33417cae829d3cc663ec6554fb9300010bfbd8db99d2628d4f81a979dc30945368346edefef0955eb238899404fa38a32621ec93f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96aa41c48cbcc6eeff05ed8b3a71a04b58ed9de8eb5353c3e6e5ba66824a50bd30cfa2622805e7f86e24453cf25cf119efc841a9a4906297042b77adec76b11a6e29e14b3f28fb077481d9dadfcb1266c19512607c0b24287987bc8a469b50bf7b12eb11e9dafb01b734ba06ec7edc15db5e78a12df3b6f9ed09c8bf7f74ce17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he902dfd8fd31fb71e398dcadfe6ea2167afd6bb1f3bb6146439a3d650c64c8ab357582c1af6277067c5083c1a5b4ade4e3b9625ab96a2420a9f1400cf208a23f757231d3f9845bafaec4a8a406f29d4fc571400ff07ab1bbb0538bcb735dcd31598b465da41ab7deaa54dd5dc9886f0aa83c19d4ae1fc042ec9ba711a82c6268;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbdcebf13a2c6f662b2b977db4b185d35e0b9ba7930c11941fd48e79b0529e60e52138fddea5db592085565dbdecd67559b191a62d02656f0810ad587af16829f1b4494ea7f96eff59d792c43b7f46b6556073b38be925ac4f34ce7be61f3f47536b33f2ec351804ec9cd5d4fe71a345d786a341b68e51656ed3647626dea5d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97c39f372bc0eb9af151d5009c3dbd27d4b8ed6517bcf7aaea86d02f5e04ad2068ec21d70cb4cf995deb457893ac539853d378b67fa87323c27713abf7543bd8e9c979448e38aa17c86c1e5116c0027cf16a88a30af830cf82a6310faa39a0779b9aefe4fd3cc6a367367fa88977fc2428e2933edbdaf19be13a4d2eb0cb6c41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd03f407d6e7c477906b65585ad38569a9c9c7fb1f3f44bf9071c08fe90e030b3e8a26c75a632fdf662e10382a236aef463aaaa1b15c19dae3173310c62cf103cc36809ae0106522b7d1735665e68fd9323f2b7de8725931881e5d065205090dfa42e4332d98ef5c249c10c66b49c4c2a4a2bedb5ae454d02928a2dcc488aa5c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d6d91d163a42f033c0f3dc00e57ec7f8106f91c705adff35741a42752041c2ca5b91cda984a30e8297ac15acdf40afde50bd2ca3e89c54119309d3da59475640028da17dc1aadf5be4742c606accf7c4161b75b4c8aa08819cc2348de30b5ce1fa1b338bd340cea13062f6ea51bbdf80c8c4034af823ad2e0e0f92ebffccf86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3553036a2844fbca55e1c2f2c5c8e8f513f506e6b7b396f138fbf3b96246e63aa7d02a164a0ad3b24d5eabf9e5be0715b9b3df76a804f676abaae598fde837115a7f38fdfae11474c8fda257030a47af07b3bbbae30bb994283bbf267256c3c7ff93009d9b22e230843476b7bc6fb22f47a90915536a1ecdf4cf71ec2a65fbfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87350acf21e76e434b3ff58252215c0bad3212ae46c5e02cbb9cc10343dcc5486530ea0d8ba21be43368e9f2e035d704e38073ba2fa0ee850ca909d1a592dafd59f0612a68d0a5bca82d710d3816a5ecb9ad1ec6526447bd42aa0c4a2a66b2b4fc24814c5c47a60c83fe55a0bd26069af2ed318dbd78cdd7f9f0561875e394b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4ae41c78b18b20b4f49a798e59c68b647012abbed732ca95543213d9ccabec6927132ca98f886c2734058751a50349dbe64890f1085f3cb87a85cdfaffa6826cb5365eb0cfcac60be38dbacd987542f7a7ac65762ebcfc279a3b7ad14423eeb64ad60a5322d35b5850bd2eb5edefc0c5282c49e62f04f7872cadc0dc0149404;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4251f9f9148c911c675cac7f5e57785e274bcc38578f1eaab78e07aae85281d08a04b44d5461804f94b24ba2aac3296abd2e83f4b2ba639a6a606b97efa0d5ee6a3db43e4b59e46f8066a6197b1b93d8990b672c4d2a11128634b3c09ec49be6fe6de4cad312668ef4a0c7ba26617c90707885d0bed6f6226c7667c84b754c97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a69ed95ebc8ce40817900a8730fa7d3553914e07fb02e18f3d2bc6698f11f8b8dceaaa63637d7c79661c4d77a81b0f7d464a5a57f5133127ad601c60b02e2795e45d1e121bac7031a8f4ca68990ae777263c342da0cb8309e571855c67d2d65de48d950c646512a28a9aa18c47e0944c3bbd1a1c9fa9001b3dc5e198324f331;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9a6e63620d92d1b86235490fafe11b703c58a600b2f8a9246977e4b05f1482d628918847846094d739b7e118f3de42e763cb58bba9d15072d28559341c84941e5ca82e133d904c8031cb5a495fff2382f15e906f15113fb537d95240d08756a00d09ba9a2c003e8c588500584ec3d183777051b7209f0cc3746aafd0a2cc926;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he57aef2a166263658cb03356fc806047ad38be8b8c8fd058bce30614ab8cc4c377b3e61f509bb6015080d59ce11bdc6ee76ebb089140a169b8e801e214eeda06263bd74cff6fdc413b505bc5f542010ef0bff710ea5451733f9a1cc0e27b35cc4022a387ed17c25c85831182a3c883264581501e32ec7d99adb15ab0cd6a9cc6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb9f0fea4b5da6ccea112cada3fc433d60590f3129abf7e3bd91cc9e2ed778880dfd29c707cbb09967e0c33e18412ca74cb1487a7b3541e2657010a55d4e298e9239ee1d3af05f5ff6d89b5ef07ab95b11382de77ead2ad2579e88b6d1b9f04d9e5c98054a0413bb07e990ec88ecf84590cff1bf778f6b24ba276aeb515fbb73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ea3d44c1868f3e763ec3ad0ae298fc5aa5e4020a4c79c42892d55594fae3f9046e53799141b30f419e40c5496a46fbc874cfe6d6192158105957e96388a987c021bc15c4f1b1d3c31cdd71e62affdd9965f216306c790f91b796bbc4b959470680d59b115a31de7fc66376a821dd1296b996338048d403512beb9dbdd672a95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80c0aebe685f3545e626041c7fef1fbe270621400e877ecc6a3e36b533f87f5fb8a39b501ca8117eaa70a09f28c2dbd0b3af4604ff0dc6b2cfc5bce8e239b99547a137468f9ae4b9a62bb695d612ddb536f9ffb4bacec448de230274f6a9b490b059a4e07b3dfcb6c7e061e767e65732ce9f27d30a4074793c9f52b640e719c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e134c3c123b1d610b0e7ccf7bbba73f40dfa28dd7f64c36d83aecd27d6ffc18eb279d84ae5f90e6ff1994c04ac6ef2995d2cb595a1ca2c3da3a4b9ed65ea25d0f9785dbd0c0573b2d97ec44aebd5e92dadb7ffa4699de5c5342eab26359332983ffbe1df4d10b05d2c05146a14bf512ee879c87a5d854c1a56373699470706;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h317a8f1b1dbff0a2a50d0616c1ad486bab940554a957fa94035f990cf6fe38e4d014b82e36a413294f996ab86f322db3a3cdf1935542808a678efcdd574458703b6919cdbdc182b19b4638f19426f474f000aa8cb63b4ae4b82b6d39c4dcaa8b2c7f7361c956bdaf89284f3145034db3e179b0f04ce4b23389749be19e0fbec1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6901dd732de788135066f154c42eb74d12f98300cd5e0f96082adbc4be38b2bc06e01701e05d514b7b98bc7cd7a42a402df89e452f8efc32167b3bf6cc8651eaf9f63f98735c87cc4e59139d1b6bb2a2d297b0aaf456c4a25dd66db68ddffe7475da4349151315c75b6e9b50c83bdbc8f4266144011d585b9a1a50b17209a39c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0ce7019a4007a3acd990cc364778eeba18b13b169650b44f28d4a0c24076ef615e409f4cb40d667b92e0f0bedfde4abab0f258ac9d10567a95bb0572a3d855683f8d1ba9974c63907683907f0c7256b8d8614c32812449c164baff0a602d7a2a89e1113c808f3c6554b3a3dfb9332bad166e9cf9110aa5361e393f65409da9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1e986aaf8da24bfb7afb31984965cf9c23952abeb6dbcd70e68caf7422ba07d45b39ef71198e002ead8cecc122884dba006e0b9a83260e0b701d4a9a24e874aa1ad95a1a23e1f524a76e2ad825c18af51093f214b23f2e80173e6bccb5e4ec4d4deb33a8ddc78090488597b22b91ed95c333f99ed09dd938c303b2443db0366;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab34af4b8a02aac5ba14db9cd7885c1fdf0eecfb081bb48e5ae5f7242b38e8603e2718396d0b961124ee56eb3dfe68d1723ab924034c3e426ceb7fd795a4ba7668a2d3d58b94841d5323ff06a474fbc4c544f4109fdbdd6d392ed8a812f5952594cc99b238aaeddd671d896f93e0d1660b56d7559bf2499781647a325d3839f8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd72a81afa8f9db197ca70ba2b2ba2190d17625fe58c1f7cefeb3b5e3c7951a4ae8ac43ace751efec2a9a1e5db14836fce723c223cfb3fa129d020bad7f1d658264e2516015a66159b1d463b9b309548c3b726cf7a5458bc173d2a20c6c3a28995eb1b490b2fd55a5fc7799ee43a5bed3cb0eacc942f9d30c2c2626e8a8ddc9e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68e19058160b891a62a71cb095141f6a6248772f4db9587dadb175fd952773c218a639b7970a4ee99a5cdfc4bb54eb4f5316e3581ca54da7f66077142430c39fc31a66cc1707879a6d918d75333620bfbbcf7210e47406eae0f005f7260dbfcd12411979cff8d61341a2a235f4f9b79774371b79f9b70a02f563867861d2bc0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59134660ae09fff9c8d582ba722096aaa51f3e845666b9819b0ce6e1229ddab76c367e7087052087ed42d967835058387441d7be196ba4a8af8065c9ee5a53b94c7b30db2355783e1e33903b4a8acd19d0c97938906b495aeb9db881c4ecd43a54cca22fc50ec8796d66b1734bde6d99cb98056d3ba24d62fce4cff931238a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h918aad6bb34e87591f30d3d504d45ac8b12ea8cc06bf5a2e4e3ee5ee74e1794f020d9ff12d65c7ce90d2365600365dcf07d416a7ae31d2f4859609f83b93e7fc1cff486488ced5a0d03827fc66850d74cf0b95d1ee44d9016cfd53e33928b6b3eafce79b4b805b45239cae0f55d4d375095900d54517866b0aa5ee27d44dfcd9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10c2e2c3615a5994648f6448a76c30b4ca942e484857301f0ddd7de3599e160a9910ab3eacb837d72ae567acea4181b8e527576b157c8ef9552bfb3fdbb87d9515a218ceaac43e85d5f6507bdb22ba6492972eb8597962f6edb0116a9c2224627a6211346e531a541aa30bc076443071c65c85d4e2ef128bcb8dcfdb0479b096;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3438cdc78ea23be3192873736c04f3c41d2bed5a34ac8df3fb66d01c31d5fcde891ea463719c3cd7f8181563044e2461b000cecb72f4de58115082e78696cb13ee0166aa74a07d543c7bd79ca8bc1b967e1053c93fdfcd4a93359b99a9332a62bb4ebcd71f99ffc79c1d654d6626cf2e3d574cc71af90dad96c48fedbf8dbb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd995c8c5ffb490eb067c1e88b33e108b53828f2e05691b24173d4829c9b167d7dc1dd841c536b7210364067595b480dd7d3f265def9147d81be900e3de5f2b2a9d9ce70752b5ba6d02faed99788a26ce3b8abfee90bf1a6ddb2621dff6a02db455d4e5674105b682f86072cdbc281b450f90dea6900ff72fc9dce550e4f3ccc3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5c253de751f14716df47c52ce301e5d57449117ce68bc60e05670072b61b19da42cbaad3cd821bff1ecab334395f234ea1d7cd4616b48d9f2d036edd7f4e52d6bf463dbb93b60cbdb0aea47cc5b36e607cb848815910f65acdc5f33ead46447a58d96f161148fce4c3311db7307dc4b71d7fa067fc7388dc4ebbb99acca5925;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haccad72ca3bb20f0cd22f938cf19fc7ffd59d93780432554f221e8cf58348cfb2bab6245956a30ffa7fbf6c850c22ab9007b20e9a3470633d6f4178389329e24c7a7dab7a2251473f1abf1ef642b6f7afd7ac1fc37df147d8eb5fc562c9573b3c1c0c8633e8dbe4ee5cd5c0a5ddf3c93097cdd5e87ece9e416332730a758894a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h373af7c11a7fedaa446267a1e0b9201ba01bd2fe2f990f1df24918360044f4033ffb9e87706abb4af6fadc05b0bcccaf1b4e76ee5fda03d94c204ff5c743a647b964e0b620b902f4e96a2abc06228ac7bfd4fff2743d7466de359181d5613c65a81b13b170aa4a7a19ab07af1e8a4ac44de6d35d02d7c0f98f1489574b9b4ae8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h766281bf9787e718a766f6ff136a2dee98114b38a379f7163cc2f766b1115a1f8ac1f68ff0d81d7252c7081ccb7ef6505935bc60445e82492a5e49011faaeff05e1e2325381eeaee1491fc4093b8e2858ebd11f85ca2198b4fa48460a94906b9e0fc924ac7a8abfa7b21231809fcdcda0eb6343919837b1de232498fac14bf7b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2926531d697bd71960bff8e58676027b02b5d8772b59e2c429015b357244a3963207a96319313bc1bc016d7e26091c8ffc5411ca918fd24d8dc538bf7e337f64c4429b87bcf6742a750ffb3a50d2cd991e89ead86701cf7a1b546b60ca44dbcbe89ce6059bf16a3edb73ad00de90da47528dcb22c2e9398c1e8cdce74c9a8e8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h970f4c9c62f893cedbc9b25439b46190d51075bb90329f5845e7a1b536c3b5bba2ed103c29e54a4e14176ea2da852e8c258a576f008f6006b318cbfe39b67b79c99028814fa0feddf11aaac114d9cbdc024ea92f5c49cf9b94df939b7928fa5371006c0987a9dad7db39510834b05d24490690692f33ad7c04ef0b03b90dd89c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e98cbf0745b81dc4a166970fb1b0c055d93b0a4c4df1f17d9c4a9adf9b10cf7d414a5c972918ed0cc1d645cc508f5a0ddf5c56b067b6f67cf1d271307ddce8ebbf61aaf9217649c8a2418d15df593e9816e6c975fc393fd17dd68d9a7a7110422dd53348c6c4cb76fd01f95f05cfc90be8fb17c1fa3d5a4431dfa7f2dd39770;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc93a92f47bf13b82b9c1122192d1061cc08a093192203fe42c2578ce1f546d5309626bf2a31fd00f443b8e7ded3960f709c15ac7c6f5aca4f76facb68337fbe2b32fd4c73dc23dbcc3d46b401c79cdbf59af78c216ed7663ce3309d1faad982446efb76eeb4df6eeb867db60c977cfe79578c35e516dfabf66dfa4398e8e56d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb88c890a9084507c1a26021b1a860c78ed5837855528f12dc9d31df2ce803b091b660f108c899ef497974930984525600bb38d36f7b8dc47e265b230d83d11ee18f37aec57469ca689a58dea6166e954ff99b2064904452df5a0bd25f836af5f670e50d827e77c3aac14a5149f1e6f996a2065cf5e6a0b3ca1836ca9af31d59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a3846f490915e2d3989c1f122e1387142eb94075a88d65a8e70e24afbb0458cc8f366ff4cf69a39963e22fd1d445cdf73d1892676872f1cea5fead98f2521dd88c7ae404e6755bd5f53b97f5d7cef3408d44086608794c37cd9147dd7c206803f172a9192b90b67153a6e5bfd4d596e78362a33eaa83b0c76bd9b72bcda9424;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc898b5d5e5779fb4b5880075b84c8b26a9a9b9bc008bdc699ace1cf71bdcdd1360161c60c97b6177af1d3a3645f4042e895e60590e58b573c14d0972dacf1a6f1f07e74876892ba10b827bf173992497d8070dd176b3897c2329de094569c5bee66e23b0fc1b27abf312722d95066e88404125d33c31c1c4f64deee28edc7269;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56c29f8698bdbc62f4ca4b1a5c8ea2435ffcfb71f0b977b76ea91add11fa8fb9a111365caffe1eef754251af48dd3cda4e485072c70a11b1fb44c84bb08ca8c24e2fb01ea0645ea91d9af83e9e03f78e92042fc73f59ba9f7fc832a365eb81bfec8d865df79b7e5d102d7b10a97de05e568ca9301151f259aecde3b60d672d6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58ae0176e8fc55e8a83260cd5c372266543d40f21386e461da4a2cca571aca6bfb066fd11a57cd9f9408d989736bc5a820151c809b41b0b20626b564d62f73758f420d3dc87dcd8e287de7e7e9612856d11204c0c69e4007653a8e07afdd4f62089907f9494bfaacf8d6759c02cbc0b7c8ba8bb00e1f245532783b49732b036c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2af2cbac510af47df61e0eaeb3d81c2c15bdf445bbcf4916ca13e92f14dcaf176a46ab6a22f55ad9aa26299358962001bf88a95ebae68e430f794dc8939342e00d8f836f5480a4154f6bf2a8bb5a868583f47696e96f4d9525e5375bf338b10b3012c5882d06c03cb828cb208ebc207db48c0fd750188737c68221b7f7d3f31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd97e8b757201c128574f7b147dfa010be43be03cbbccff5f01da571c83a14066b52866516a3d5f6fe1c0ae243399ba86f233e02ceaf2122c77a9737ee8ecc292457f160cc30e9a3ac35b1253322499674ba558cc33b1f1876a51a83879455df88ca0977904abd92b9933df7906e78b14b1a3bc7c9e8354e190a4ecc5a77f914e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa13eb775666ace63c0738675d075695e85f525c1ce013f3ccf95b39653542390df2cb7e95d59d5104e05accfee16a291802deeb5dcf36129b12d2250316d61f2ad827d6ccc37ff407247c5c0448b8bcfd7a6b5c7513df23d47d12317c1e451dcbc739894d48256d1f12b7786088fe5496c24dfb242b03bafbf54a2012fe035e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaef239a44c8ca11a5b5c3ed94292bdccd4e1d349355984ac6e1638e7a1402e4663af2119b0f7b772fa5d98ef68227ce24da844fdd76a810e4fe9bb7adc10af65ec1f425e68bf0c2004388c76abfb22425b4c1ab6bd104911c5f1e9c28b7df4c47fd4072cbe16bc4c0a74e84a2762efe7a0317c8b4052bbb8d85eb7474ec11e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0e3adeb9bdace8fa8d659b1d9447cc36557611e082d339fca5c4a779345839bbc949b6e988295f2dc73785b8402d0ccd7fb9a26c82c2431e9534405eced30d12683220a2cbbdab80591c9833e6ea612cce0d35806d37c803fb331054f7643b2838e126fc59fc3525383e1eba75b219fb96f5afa53c146987476fc239cef4823;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcebb1a87df33dce3def60e5af57ceca97ad4eba763fd67404fd435bde2153305073e4f36e9a54d4657de2fbe3422fe3cc1315239f2d27e14ee1091aab7924af36c5504b0769866e077ecf004ea1c61a711ea3157f32328c5dd98b88af007f45cad0d0095a6895445e8db12856b30ab84ddc38547563bd763e6868206eec6cbd0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfddb16b2d705439149f99a54eb85131537aef3bd75236939c64866b87f2c79c5d34e208076b6a9115d435a4c718779df2b2245bf0ff449b7e79049672d7ead94a4420930e40c58177b6a9e28daeb101a292ff956b7d5297f19d49e51cf61c04b3be85590007118ce8f75df35cc9231f8b0fe5f103395e94bc98c1be7c484171;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd23699e0fad227efc5f23a2e8bf6e65e2cce01138e783d1561cdb0acfce752530cd8a87eb3d6ecc6c83c30069355180cbfb3d60814d1c39c99ccf551bc1380dd550bdaf20c5edba4b283c14a84d6e9b9023616382c4e2047c7e6ed4a0bdf2d7dbcffb622d28df974f5bded45d74e88ca47feb9ed39f13e85728b09ee85ae6ce4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7270815507e90b4004bdfd3ce91e6f8fa0aff3f9d9c71430fff21d5a4f8c55e1cd4eda584e8fd7389ce5f7b01c47d577e819dbfa6beb07042e0a3bc438b9e54745dfa28f775712b2a96256c12c637245a213cefe01413545b8fb0eb4f7ba38bb77614fc22329a4ea0603414cae7cae920326cd9680232cc90f302fe653537c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habe3cd65a081a894b8a53ec95136758ead3a5ac62663308e6f6241e9681ef1fb223571b40acf5f6ed9c62ca3c96f3535ed41103e7949ae3dd9ace89866e4abd3cb2e00ed0d5f740f92138c9e5fa7ab813eecd7818ca9740a99bc4a4c747c05dd25481a41d146bfac342b42d46e71fbe1ec2255d209316fdfbe593307cd29e37b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h876c2e7d27da11ff054236aa2ffc73ad3f5567c4bbc100a7dfe9fa56a28d14b51ea353ef6cdd31c70a2e88833108307183475a82a72db6e12b643d13b74b6f6a44922aafbac7b257bbefdb2949684e83529b34190d16b4c7938b0ba885814e0ae1bddc4a8e1ef117964e37c74196aa3282ad7135d00ef565ce29969bb8567258;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55bf1ab58469424d18f01b77e172783ee69a5a868ca9439a8b51b35b9f527a1119decfe81b73690abd73eb0c3e4028f7a6fc664fd45044f62fe5bc652be370c2273c82b2e211ee50cea18b75bd5a9ed3f3a8ad2bc5536061e48b8aec5159a9f7debdddf466ac7854f56134042f3c0cda568a822bd731c6bd4d4cfd7305a38fb8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb5c0eb217a27e5c780ce884d17a8d398a849a77defd5ea32b25da5c9961b601c0a6b88d46d24c5864c91ed6f93a76e7dfca9ca6b4707ff09b9a733593f4f671becfc0b07104e8f78682aeca3cd4ac9baa1793fe4359516862341c127f3f9e29af511c0394a1d89a47c9fc94bc052ed6f6b3fb0effe4e08686aaa6a11fc72215;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc89af6edad094db497617b10ccff0a7e84720ad54d7c11207d1f6625d76407b683769430f67b6a6cda5db2c156debd597606b65c2649da621b94f08e1e20b99e861265cb66ee6565f4131c4a6cefe1992f361b9b3febdf797b0d74414d1ac6ed29f0ac49c9ae9f4f63be4eb1bb7ea257cb85b0e1b5cd73f1d75eb8014a1f26c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce619683267844d9dfbf982e40f3d6606428e0e2d06f5e6879edd4a49baebb590f9ed45d950bb2cf2b06f051260fcf13cb011fc4b2ccae92559fc2463877c70c4c5b4ef64d16888bb2e381c7ad11023a0625a13cb754f5637bdd47918ce8d85ee0e7973c0a80ca9d0c32ec28ba446fb53012519fc882a9c972773963fd5b840a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31bd07283c53206e7360d278a92bff6ce94e7c95d606b0bd6e88749aafaf873934ab3c97fe7539499672390961d8720c3c06e4ea6ed7c965734395f2ae17cb19b2bb20584377886ae0d451de52d87e326929dc9470c8d8d6c8e3ef103dd54728cc44aed765e85d62e26745ae6efb6523825c29bd4be3c17bbef872e6f63ee6f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5eb1a63754e0c17f543ef2535b766a161a70f5921113fb44d3606ca062814db90c1b8b66402882a5062c46691e6abf9f2b602d32ed7f5397399132195aec0546ecfe2dfcbb995654a8111446b470d424713d51a016916a1a4208836084d9206a04c4e32645cc3e49f654b0ad76f57172784414212c0458844ee2827dbd8420d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd4903657b199435605ef06d45fc3334158bff6d768867653888b13f67ec67df3b9499b109125dd7c43322460b1511a3489b1053aa777dcf244a3ec95876bdede74bbb04b3aa79abf6e2aca02ffc38a424c3ee5f80efaff1ed37869c1812555e88496744a8256152a2ee9c3924cdb0fdbb4391d6986a2c74a6506f323236784b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3679e934719ad5a41cd99cfecba09180cad1209eae8e88ff88f85a8e5f8089dde3688350ed106a30646c12f74ab24b6840b48dc22670db1525def20bb954f95ea690c0fe55c031acca0c4c002333f4bffcbd0a390a0a6372312e58d41e75e8a9b6d0a53bc5129a830d3eb8ef40f5fd7b3786877b8bafcb3ca2d9f3a2c0bd56ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7723ea89f5182dd4557b2c5ab2e2e78449d4b52c6887a396d89439ec50bf22784e8ffaa08ccdf2132c81816b5c71658a6e825db74e904b82f5932b076dbd2a0e9c22c1cbf788b709857d7a36cfee219bcb5a7b1a2d31eb4b66f8134aa295a711f7ee6c304850f77a56769bf35d1e142d97a75d0b092afb6b06fae251730812b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4469d84e9a4c8c4108389b05e47844514a97866d5c95d029e27c3fd54d2d8325858486760344545901f742994b80c0ccc838b09f532b35ce83a7571af89ef51c5892791460770f4cb41b3a45a88b85b87b3f3e7528f73bf9b2290e6d7cc233f5392ab3072e89e038cd015b2339bd6db8206a94b856476d8b4bf54def683c7a9d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92129a2b2e66e23eec419f5cf9800e9c6f2b447ac87a02d17984e2d45a089d43a5ea7e519aaef255e990184b3a1ede784c67e63963d735b0d846adb09f684cc7fb46ff9eac13abd1561c859ef15d6600c0a4513ffae738df603fe8e5ddb1f1334a1dba0e89cead8b20be4edc1478d05661b89efa3b063d07630b6a0124c98c9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c964b79f425374ee56074ea72d07c7c8cd9d87422b515384b1a40874772a9043808370ae1af39b0c49a03da9e4b6219906f9ee5f93d76f83c24d509e53b08d3603f59f1bd560b1a2de68046d396062933e971b66ddb262b8c8b98189b3df2cc158e8751bc14890fc410aba8a4d28a64399c781733fb078d7b08ecfb918adee7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8481f83a0988667e77fe12bbb1000075ae017e11a21d4a7959b52091c6d3427bc702b20e5b185e1cf2ce8a72f522078d165ffa951db7ec87e741532b1d534367179be511998370501ae6c6adb3c512fe15955650a55874c1639ca2942e7dee9b9c8e15d5799e1c7da19226875ba70408092ad0cdbd2a4995b499f4bf76d23073;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6713cfa075acda27b4f28ccb508ae468deca53ed381e747438266b3c262d2ba6558e1fd04dd75956aa5d1784b03c3b4f82e74bfe4c25fc914b2c8e65cbac4ff99970801fc0e5d3c51d7c6c079f0fdfc1cb57cdc38945ed4ed0458dcb9011d563de1becf2ad99194f3603667ea277fbc3052f572601a94ec23087b09135c6ce7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86c842434c672dcbc1f15428331a91f4249743e9408932b8786c204e5be48516806d6d4887dc1ea68a4170f0d9095f6ac61ab3332aa9683ee70610e40cacfa694f211e944d38e363920d3333bc794404bdec55cf0f6742975504e96d3d8d943f07ea634a9e827ab460fc4e41f2c3bec8fcf37d9fc0b14c9181d560943db2602a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8960fc2fea50a45d2963b5843cafb78e8ba6c4696d57691ff087382117b0890bfc5f21816bd3a96fd29415cef7f2badda6b372fb6859404e99fd114f4644d85aec00b3c3e84b2ab3009ddb20c45762d9512cea99577e7d6f8c387cf3fc59fc73f6c1dcbf6929105ce2db543dde40fb0eac91078bb24b29ecfec285af0d9c8ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34e49d64a249518ab3319a567f2c3de5055e1d1016632e4bf6b18cdab720e5714151695bf571528e25d3bf792a6225c737e99507c7803cf9900cd5e896f03c83197ab31cf5e6870e9d363de6c831907a37113fdc97660cf194e1f272f7eac0de15d1a2f4b1afe9808c2d28c72eb81b4f172e8adaea70d100a2cd3110ebe15a05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50dc16a4dcfe77d540803024329e6bb9297be02b33229323703fd9e4da872dfebb44ae20bb0e4933eca3071f2e159fca6b20e4dc2d60919a35cf7c61ce6f96f130b5b7d96d5a7346e1b09c9a43d853bad4de4907f733337efd01303aaa7bedd80b75d2011a95a3ef07ecfd56d5cc6040118151f5a42f2c7a027c5c19f57b17c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had573dfa3cbd93f379b42706b4df0e07fd1f4f146780a7089e7e2e790f1115fbf25b925ec4bc131047acc83eb611916295f056cc38f0b5e1f5426049ba8a0f32fc5f106dabac0c6ce9ba7cbeec725bdaeccf91534560e677aa9494d48e8a6f43193c2a1709c497955c3badc9c5bbf39ff0ababe012f303d49cc1cc528dbb02af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ea51503bd9b3251c9b5a6ec460c876f6221f1739f88093cb771e011b8b8edd6985567c26d77745da278054690ca99f613fdc63528a6d832adbcd186af163d5a5d3722f785d5c1d560ae43a7eb63685a5ce0947aa0e98ac34b6b9d09ffe73051044d1a4fcb7bed970d7673709ec966dd2df2c27f239fd295a856342b5e27a193;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haacae9402bd142ec655bc8891d189a31b425cf311e50a8dcf75b6d1a2a79aa5f65b2dc5cd897417021792e463db23ba00d6a02606c12e59167246bb69266184349cab7abe2423bac47e8b1ec29ef18ebae7f87ba50f68e80483b04395c30d45871ef438889b7e3883680b37b6aa519ae3662bf3ea5a755af63f0103bccafaf4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74df7e11a7391831e0e6a1cece4f3b50c7206bd743a9134a020f518f108195da50e14b261a128fe2c9ea50d7b354e8e532308d4bbd0938d7171baaf304a5d3ed623d2e071afc4831dcfa524e94060d3816d1f2103b80a4aa1f23ef79437d7b18ccc15d2b45d2af57b1a81c1637ef3120608dbde838a58d762fb0438ce70109f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e697c43a1dc51863bab2c16fecc74808ea49fe46a1f41333eeb2fe35d3830f46ca12e3b757c222ee4c73659da159c5a82963d31e3e7eaf2b28dd5409b3088e400603f56d78ab8987eafb266caeb9a2dbfddc2d534641c305408a004f1e8dfece642dd7d4d0cb5950f4f582afa113d2e2b59031bf7c4aa3f053b8df53bd45b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7f7a933a91e4ad1384d5e09a83f21a51cb86d80412c352f69159611ffd00f3702122b68951d1200580892fc32c97ae9488679f1abaecc84e39124f35f75de3b1d95c1091ea98debb1c9d73e79db84401d43e1e2dc1bbdf60c5810b620f2e6dedc1449429aace54e97c7230eb869160d8e51b742f8c7ae7f14a667ad087aeae8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b411eba65f937460442750bb134fcd372f6860ff199d729173e751d043570322c24d278c732799ef8bb1396fe0ebdcbe064de4270acca4443acee9c4a6150050c5c9a4651464bf944357d2d88a13169fbee816f802e995bd0170927ad292e7c3133f3c609d5ec3eb8dada1c64e409aa6926f89fe5f96332328a57bbc38aa54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb65a2090946b94888c3aee113ff59fa63bc7cf6671c232921db4b8c21017ca368abc5210a3a4140a3ddc228126e4158444a5487cb390170a7a82e9a0a79e94b15092327e36948f2a186ab90caf85de368208a626cca9061b1f7ab24074ce2ef09e1f14e4337cf3c9db0c45d99c34aacd6cba3ad0700e6676aed43d36572028c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haece151b4a0c9712412732f13df58e2b8b05b956948a5b022db290fee3e0312f6c6348ae4ffcfc98f3865a4ba41ffb7c850763253e60d1850a3fc03d418da3c92db57bbb33a2a283b033516dbc7cf219bae18ef676fb12adbe909fd886d9c6c74d9565f7828447f57e095b1a260c26ae32aa0b6b52516f552b934dae8a51b364;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22c10b589e70b04bfecda611e37717c304624d165f896f81d0047519c9ad4fcef13d4bd21ee0e0a079d228153f4cc77f6c23b995d1a1999ea1861f44552d4dbe1eb6c33e0cd34df3ac3d1e58323d9a15f7d85b60e592832d2bdb4b0889b91db77fbacb44367c2cb6640104d4e1a9b1e2c1ab9343f3867d210b2a732373c362be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f6efa8107fff5a6d50fee336c70e219e69aedf13205fc782a8cc9fd5e811b9e32eee9c360ce3e34296818259afde2071e1d6348a5ba356ff76422815362b2f0f53122bd51358b34e2b0cf5a1f6b5c0506767701334bc4e749f2512d6676c41ea040970301b3d398955f2e6501006a676c76a7a3aa99167f6c2cc490e8e46b73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a197e0b7ad21c7201c4e9437d54972e27b8fee008074276954bcdf6088b57f6706821a304ce5ca97888f5e21f4b00a72983e7465ca6bd711083021c9c3d853f74960d68334637c147108931d1177e115ce8fa626dd679de27604808e82054b6cee56ee3671b80c2a283cc813724058c7eee3be86ac4f6b258f9ece571828d84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb0328ead36958c086b02e96928900ad54c89d4b1443820bd222cd8b761c9ec47ce05efa52b5a14f2a3cf08f69994a382f369d640a6b7a5e799f1c3da3426c52c2c89bcd6a65ce8b79e6e9a97c170fc073d02e388c11dbeb8d45a9576279385a50cca969b5a1850d64ce94035e3fd17125bfec7b873cf176a02260fdbbb86f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39c202342f43d41d9640f1b466f4870792f2b2195d9d6a5660d471f6097c1d19016ce247183faec1a1376705e8ef9979e01b03d20600e513863ce990f566a68b029dd2156dd25e175a6b7efe90b48c2e70e0650e347b9f1d66233d1f32d9e27f8d4f1ec30d21d997258dd90600ac43697778bbcf72c45131a0975163a3ed83a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hade18eb8a66f3c509e5bb6ef5696b05f305358d547a39a55285516b66a9a0939d69a6950040aa38df2bc6d4458eaf77115b2e93837c56c9e1fa49cec3c3300f060722d291e24e7de09c0ddbbaf794962588f8a379d95814b0a7b54e01301bcdbda70ea43a05e10d04dbf752bad4fa8a34280f05b3c3fdb0196a587af3fb69e3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf47742da57c123c72bfa49000f14b2be53a52302f0f989bf642df9dfaa2c33f4b7afb57a146509eb23d3a65961a1985b1cc49b97391bd6e45640e1ec608ddb6d7ca9ca36c1b5426228a7055673c00f418bc0e5a85bdf3356a8aa52e8c22c2b3d0f30e33a3163902817d4f26b1c54787b8aaca367a81be95a0ce577c3aa30434;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1e6da640cc155821a2e3bfb571ca12ef07e9f713eae15d7eee75534b86ab52d259d65d7c693658609cceb76cb91f8ebdc6f67456438e78b34ab46862db10c75d20ed26c6974c5fdf16d173e273a7d011ee07e80fc3e3811c6aad02f1674f2042e3e9c4ca8ef96b2d5cdca8d2ad143dd1070c2708ad1b750792b550e0b031946;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebe44e7e5312492f545b98072f924dce2f474a79a5e5d037d5b4763c85759e2ca716be01675eb69dc75cf009fa6a8fb4d22de738146122b9f20d8dc710b2420f3dbd51f8d1b374156274dc204c18bc5094706f121a17838fe08ffa50d095c13e61ffd4dea89968282834eb9fc40560cdce6a8e17d5cc6b45c1dc9ea2cd96e6b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h413b1bc47c620e9e973f84fe8125e7865a636e5ca0e777ee142a57468d367277fe0bc1f580b809f0164a50ff1417bcf750d1ed43824a51c40b4564d63f95c5d1012dd98defd77d979d3100ceaee485ff2d6e3f76109f6d87c24ce5403f528d6e3b8b3908e8fcfd9c881ea9631e5e8c67552b48460c7ee17b41e526742a039906;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93bcd6f93b73e670503205f21a33c12b8afd7088162c477b127c573f83d41653b6e7876983d7abdb243943e60fe41c576bb1d4d410dd7c9c122f7188c6465eefbb9301acee14d24768c43f9c9615cc0cc301b4167031f824bc3ead9291999c746e3016b6d01da59b5c43c4744475ed7fc2694caf502c5dff52f4ca8a4cf07bf4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h772cd74a52fca1bfefbe8d0521ed7d53a1b7f4826d7866ab373ec1a301b830165c973e6687d262c09f0a4103309557a111f3c5f446be9d455e83786da92bdd901705dbb2274fe40645bd1eb6cc55c435646443564c9ecefebfea9afccd5b6dbc7d9328a90f7cea8587a8433752b086dcc2acdbdd5b24a0d95e16701cd4d57b07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1653d82afbf6798533593dbadd013ce493a7ead98d92bbba72884523749861446741301ce5b8c72ec3d46a57e9f2ff9d24c19e752d2d6daa8425fcf390eb20695510e6bd3777dd18761f0d8761379109ad2fcb55eed857ead8efce6c9278a87e017e672998a33d2508d7b6589395fd7d3dff76bc7824e33369a42c8eb11279fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he00179c3b438caf151d3028c4f72dac9be4c395ba68a44aa38c7bb39b2d9c728c5e24ad742b4a1513c0d4449910a91907704d899e8480a5c9812e23a8f526c00c7808809470ba2067bc121aa55888e59b7f89f46f49624d4a06c68d5c093fa115e327f2e0c936af2091b94ddece2d4fc2fdb3d7ac0282acf1d42e9db938c404d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb822c36eac6b97963a5cd02603ed35336d98a2218a003235cfb2782167427da0cbd44aa67b0c42c982732652d5970c73ac77ca35031397d34f6e1137da091bd25d017466fda2b86bd27ae5673875379c7e84fe8c0f84829a463b2e3a55dda258be1b7a18933d86b5a715b5a66093d8fa4bc3cb306094a78ee47bf2f8406c0db8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91c279e71c2db011b6827f3a34d2afaa56def0835249429865bcbecad48044137992db08c4eca11356642218ff29574f80fb2ba99c1349cdb7af45ee72e4577f2c0b2dd019810842005634d9aab4a9f3810e1f9bb2359f3ec06ab885d635a8c5142ef0c6fafc3356d1ca2164daef698dfcbe1d94a445956b2f33dc937b7b939d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3c0cc7d6a2c31ccd09524222362bbe12d02884487baac884516b8a1ebfb71bd39b83bbfcdcee708ffd9a652f6b9ab6fd08096420c29ebea67495696533de828435d48156526b5fc6edc9447b976ce8cb8b13614dc5c0785a5b20fd2bf8e85764af307636cfbc28b31221dc1bb1cc277f4e9052027f1cca49f5560f30daefd0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f9da5cf34d0e2a2d5ca31db5394e44e8895318875a518a2318de4dd3a77819e942457f56cfcef20aca6658c6321d7c7c0166ac28800ac92681d47ce7837f803f3ae5481c3b8dbad65e41c3bec96c45c79435fc131a3c3919bfb5d2017ebd8c409baf53444d0f4ab8df96783863c32fc7d4f60cb22d4ba3c4a21af68f988823e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdef20305514f54c05ae0d327d5dae1064a2fad4a386337659299f31a66471d7f3547039f0ff0d8903ceaefdb1f67b3515902457ca13f40db46c88b08950278ee4471a7fe9a47ceea53119bdfacfdb6d5d5d913037162c139a382d6fa4a1a0652c865da34ba83124cc7d8c9d7ed209b5de9cfd9889407b4b7f5f3144afccda0c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8885c80da2756fc4129745c0a05c5d7f678adea39ff265ff0a73875b99b9a2ceffbdf3f963f6ca3c76d4d791ad515e70d9b0b83637f31cb0463c023b72b4612c92bd79ce0dba1bfeb6a5fadda232c23171a430b673ef026f7de11249f101e6c4bb7ab0794d5daa0a66b384f4269135a3d9dfb51462508f399747c36b740d291;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8cfd1b9c8ceb3f351b27c5bbcec4eed9fd70fa32838a6fd3ad49e4e49a0c760645c2d7cf6fb1872e4f9cbe28090f11ef848dcec6d53f27024e362376955d3f8e87a6aedc3e6533509c6b7e77a3c74678901f07b383ac0e61d0b10db332e6d7188de861bb6b7f2b60f9208c1c48e4cb9a32932d77995236b3797ebcbd2e49c06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9122e6377dfa457b2fc548f50126d4e18bfc53a87c93e67eb8293f62025047cbd658536ece099b80bbc77dc6131ac2265959759201e44384f2e6e466afa89c99dd2ad52abfdc027ac7704855ff2bc29dbe80fa7741f01f898f6dec87d1abb35b399061cce57a2744d42bbb278d275fa243fd5bd496d8cb7db281d6b01a9c8928;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha642f6d8c7a577b285bf11ac001b02c2f82cbe287830214059229ebe2ee0291bdc9ac674b28c0b293e2befcbe8cf4ffb5eec7885705c41bdd9afc1b40898f5160e72cd226af652e571bb0087c93f45c2fd65ae4fc362e459b0486e95ba77f55de19e401f32a0cda7bec2a356356f8d4c6152d040688af455505d16e5a21b9cc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc0eb8422d5a60eba92b497ec4908f7e6c4d500a3c58abf2ce9606c90a38ccc0be1dec074c41cde173102f907b0fd589dadce7092d47ad74d0ebca50fe867ab936466b475ffa5cc758e1ddaffb2d1984d5ed990130af6a89fef82b1543230270203b20b0da6ced4f0a82d9b9f170ce9244af930fa2728235430136717ec0c363;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h864cccfc199b8b8ebb86542adee7ba01583312375c4442fb1090ec82ead6532ffed9dea87e403bc22ced54fc1346890c294a67d5dbdef28cbeb8482a92421ffa2d628b3c405eb966bf007fca136d5e9e682ed2493170389873b5ba9bf62d9b023d77975d14a07c1424fdb0942f442257f5f5eff33c4947d762fe2a5467791ec2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c68b9a7774bbb9071643fc5d73228db7429f011665c453d083eab75f6a926a635b27e30e403a064c5528f4bf26eed28312d62e009d0845adfaefd0ecdf6808ba9c44ee358c3278e2ac6192732289ae4009365d4af450520da01006be6832f42b584d4e2a6b65d453db6e89de7ec42696496799a512e2968ff2ee989f6ca18ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h910c5b62bee23a99b254a118fea1ccea6fc2bc8e712cb45649fb7a0964da6cf19fffa520310798caa415cebc2b7437add7cd349710776e4532ef311d161befd9ac2a15794bf413560bcc7708e46fc1c04054fd1448acf755f988f6fefe9c139b1ab385bac8299668dfc06a6e0a012f1a3436f766007ed34f1b5cc405e39ea2c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3ff34573e05ebf15ce2d700d57581ef13d08eab3a97700a2056e5c56a0645045744ecc635fc1d045458ba629946b0f5eec67a1ae9a5deced96719e35e454285c7d245725882a0713df05218e315aa2323b9f79c3fea5adb6cb7be3933f1343332abc0a0ef19b979d9e5f6df5c41448bef8d183e71387d263b27010a7926fe1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a1929a8a00294b01e307cd26e7c3131f3133690998622829bee6564f32a1aaa10f6c842aae24517b196776776cba4dabda4d3ee59c9863e03e4a792c2f0bdbdcb10a4feb3c7301e07d8c9955d838f6e658790a402eecbd9f044ccbb6c42677dd4856103579feb0b453332bead56712b04a9dd7853e10692bb9267e3628bd8f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h298fe12a9311b8930e697eb17c2ac37eb06373b7488a1de095088ac019d7b90c67479194e7dd25dab66da8190ce56de2a72003a5a906f6cc69e22a4ff0718f6cd13c918daa9d195b1e8009e93b9d4e9e78aa793818c58b105dd18a15d114ec80ea07d452798ddd40c5b1fd5b06f960b4ba00d22395e823f3699a3300706e37ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97daf6d049943ace1d5a0fe11ab401252f62f9665b9ac33d834fed93249832b5c5b5b5259839eff4e2464719b7f38ec3e52bef3d3a531219abae36b419ff83c28cb306d012ee114a1d65ec80a979d0d857adc7ad94b900dbac78346f94092f9b6812e0609deaea43ccbc97f00197d238697e262a66d5da0323fab9b6a048f074;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66bd68da1a62bba32141ec29eae1b25148070faebb92c54641327260f17227038be8ad2d14dfdeefe5adfbcd1fbb9b8782958c9db867aeba51b87676a95164d44d7a45dd2959666e642a4a0d1ef4284d46e770c7fa89a1c105bc8b8b26e3d0540b531ba9f0f9a7257a237cc6e37b595ee090e97c6fcdbdb70e4fdb8ff0228b2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae7aca976973f5422c87d8e8577b70e0787fa871f4aaf66b4f6834529d8010c728e4cef38f3334cdf6e8b25286be82febcbff087cedda0c8e9ee04e5a6439076ff3ce2d7de5cb726c1f8f0498bcb7de2eab8f89da648e87e411311277a32434569743d91a6a293ecae07eb74be711904eb83143b3621f0305a184decab10ea8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5627e8c5aceb5f237776355ddc3c7eba7e62398360d12e778c7bdc4903e39bfa09799edbd95f2fae83edd6acd0724eba0caa0072e7d55e8e5ce71fe5fe58ad3f727624f1abbbb1307e85666834770bca3835aa4aebf15b5a26520c6faa5198cbbbba4b1a6081da5d3799789acab1b8ac45a285a4d78b1e2b12a8adf3df5f7d9d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd4d5874eda3fb9dd98e0ac52ef80c6baa2c697196223cec1c97eac98a1b56908425a183705327ba34ad14a4ffd504b490488756bb81695dd97bffac7f1657baf2833ffa23bc60e33e2d24450859cc18274a88a269181fce32d5b2e6b2eb1ac46a5b5f0a59bf6c43fe2ae43528728e4d7bd0f1a1813692d828169ccc824d6c1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e28a969d971ca8772c9faa378fb2aba253f920179084eebe318f09c41a56fa44f16adc04c69a11ff36b23e494c5257b0985dc9b137947b98be0264e21ac6eea41d57f4573b7d5b5fd1cd7dbf4b9e1390d1f910b69e559c5180e1bb80a098bbd9a7ce257b3e9a9d5c47369df3b9ee504ed8dcf8e7226f55ba61a5db9129b3770;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c2f83027a64eb37e88f89a7c6d8d7c513ecdf18bb09ec79ad9f0e3a78a95282b57a46f22893fdba8955edbae0c9f30cc7f97935deb33989252eef6578042e54b12dc5c2ec29c6b129cfa3995027703d4dfd621f2eb0d5e97e9aa8decaa6380f9f5437c46b4958ac47e909c0558f7412f98d9f2770ef308384940b0a841bdaa6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40a5eaf0870e3ad602e984d22453d6956843588decd9568d11d70f6ffb84717b997e3e72f86aa50b52fb0e57a119995d09faf1fd58d24b0db122e5048911605608bdd1166616213fcc9d6170fbc5ed0eae35108a15093b215963133ae0f0b7c2c7daa1d9decace849893b1c38468d8fd2cde3252bf32e4f03612aaa284a2e3d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb46ed4e4dde89a860ec011d6a7af79c32143535414ffa7a061befdb5d3de1889c80a17540806076437b6a9f2d64d2caecb1d3a32a8f64c82cc6a80b4c527910d912e99bbf93ef29b8cbcc895fcf6e3b96514fe4146563352255a669d315a0a2f88693050e4636a0c34a2b225285f099f083556acb38aab0f391ab6504046873f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h321b0a7da8aee8b580e7eec760abd0a110a55572e055e265e2ef4ad63893a52391108b0c5db98e4e6380b3c5554af0b5016e85f51d4fe11d2ed19ba999537ad43b7fbf4c5ff263b50387bb39e01c49f86f61659890f9598387b87cd87823998610038eb0c110c6456a85f5d87d7dd23f8dd1e92661c906663437f048f95cf6c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dabcafafdfd302bc6a979e29d7ae9fcb8a51cba25208d9cd532a7640ea6bf9438928f7a52ea39af6fbbac029bd094c6d7f5cd93b745a9694c637c5cd8943fd081e1330a3f1be6dbbe815a536f050a3b7633136cc7ba5fae7b51b656017767ec4fed0646c2bc6132d9eb50f1502bfae16ee148aae66f0ca9d6d415d02e9880f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ced5913c90598993a67926afceabe5704bfcc71cac5f83a90d85be6aa7bd660dbb86da65875326b0dc4c12409cfe25122f686a1d066fe1ecbc72910a87a8f52e359d0c8a756031310f886a9153646e9eae2cd5ff16c33b4660c691aecf24d6fdd67f1f708aef270b1139b3e55da229f5d12bc0c7218f25ba44aeb17c73bdb2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h399a1190dce0ea6f9f8b26eba8198c012f074848ed018a65c73beed53f025ca5b0bc6cb1f145e56ba2cc4ed81db3f6cb495adaaeb1f10968ed9f9ad07fba438fc0551a9bd2703aaebb01b99a1ea2c096ab9bab84f261c7c581a157008150fa6d609bd580be450c97c3d93eb4fd237618050e3d641caa01eec486c4d574a4e354;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac59d4fecd65c5a687d6cb5bf4fd8a1cff187b92799f4cd1ae28765d09efce0070b9e0b83c4fcd8ebf57d927255a95af5971403c1ca9d1ebfd73356180056f2bf0e476365be27096c23d28b11b3d78ef599e05ed191e6f157b802e82e47cc69027981a920c2f1961e284844919702e3dc65068003a2dc8b6db84bf4deb9818c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha647139dddd613b2974d6e3d49676c0b67812774d24c2b78c03b54c023d2a900bcf0a923275f21b6b5d4f7b3dc2d78a694c31fcb5235f5f8d1d70cd5470f037ea928f8f9c480168ca7535037a78c6119527fb23bb58a4a34b1aa981273cda555b7dee5ea2b22e854c71865741d15a56880a25ab7457af3e879c9c2c35a58537d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f06a916eec9a2931166493a532704c2101ac322f9ee4547b47ced29910877f87a9f6df91a342e19be360ae1e80d56fb9866186fb97a65e6e90a5d4117a23b6af33635a1dcb4d64a11229a99f928ff62774f0f9b8705dee80527276aa99426df65f8bc7b32088eb1ea1f5587541534971ac34030019cd8ffe87171b9e649b849;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e69cb11727119f285c5d40ba7f9e13ccf24df3023cdc200d798de261d232966e287f74fd99464605cc875bcac3de9a2abe2446a341993053d395fa52f2c8dfb09eace012de8d12b8c7e7cc6cc3474cedf21858ab40b5f572b23474bf3fa4c9c1cc69c3e264f0280c868efc9d857008394f349d79368eb5814124f1f7912a03a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h143a2fb09cad6122ce07a04fdb22d0ab79a30136a90055d564b50088c474f7c7675a07e478344f08c49ee9ec5639388039379e202b122ffff7cfd9b343f0d75ccfb90dff69f3b82d7f4aa18f631f645fde45239d83e662e1fa27869364e9803cfd368b8c24eb20133605a04423c0e87b604c34e591a63a597d8150fb04aa262e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55e6d6f7158b157359b18fcb0f14512c522685428b5bc966537f26caa2893fc84545614cf96049c98bc4ba6a0a1ed050b76e87bce269f7bedd05983ba417918c923fdbd611011bbee8d9165b8b4cb54b080b15c9df3f9de20035444e27b6e9d2fe23d308f4105f4cc4c36aa14a70765467d82447e77a32ffbba1987cf67962f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7a841df126b48d03921225d23ac810edb3a628d3080dbe48214b492061953dc8e1252f4d5df5da778a1b4fc15cf5803d52bef8b73e1e87ea21b3db7c5267334816bab7f6fa76bb6fa9388ed41d61ab689c9ee79caca792df54284b0bf5d49203f8202d2fadbbe8a2146645a346257ab258a80ba612c7ed601f2bb634e071feb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6229cdf6d051498a6b4c2dbfe30cda25e8315c85ff0a670af11c701132aa586b85871613515aa801e9d52a91b497168e8083720589d4f61d0d28f0b562d39ca11407742aa7d1ffae493519c8c8c8fca869ca1cf12dc14d1f34fae67b97548b6a3ca1e98c284572d4363f21a94eeb2c92d7d7af3709348ef039d734038164d0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd9d0813f13fd4a70bc690e13b6cbf6dd5ebafdeb319da959fa570998e6f9ac3c9c761f59388c5e21608f5c3f19dfaa080bb4ddbbdc250009598ef721b108ba3fe3dd9bb95d9ae6fe8e0e531efb16f1f262f306003c53f409e42de6b0b2cd2f217aeb28963339a3071585d35654837a414c6e450cc7b3bc096028a090125272;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf61e4c9c9b090c56362988c024aec62767c73b0715c63e43560b5784e1924c69bf590f67b702e0b013e61e10db3da129eaac432f2538869efc3affb4d5f657f167d40297c54096b668939bfb6bd93c023f914654e869fd0a01e8dd43bd91b6c1659ebba9312e345717f336dd57d81cc72d674ed04371f3960716f8104664f98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b8122c145f5c7839db17724475a117407360c796781e5817767f26eb402b41adf872fce7f4c08d6fddf9157ba6ccec3bb2422aa979aeca23a45072a26a29bf64abaa5de4fdb6bf962123b4ee4cbb190bcc441079e4353a631571dc889a52ab14ac87c039cf4515f4d0bb8bc98f575e5e1768eea20053dd9cd5b999ce13377c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cbec34bf49f8751696461a3eabd504706cf9e753c46ab13a5a6ed82be4855ba23f00754a90d3b688c57626c455004d33c2bfa862308e0323071679e861c7de72f413240c11c6d764002437c20e230379cfe59e89d1cb2b0f1be51f8528a5371b2ccace6c749caf4093ec0838c94204ef073e69a76bf6c63669cd917b0fa831;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff7de455861b0ee1d63207ec2064587eeef2f7e6824814bcc13848f5cc8014999cfd7e0499d28fa9f66bc004e50862920b1d71fd71586ff19136d39759bb79a956252f4bd1fdc8093b0de98982691698456571337e69563f4515c89190e7ec0cf53700576c7de0d83e16833730dd038bcf65d4b80b4aca3b3a0e697a7a1bc296;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b59f13cc744e5ce64dd9242b9a4ea80c549e700ed619dd448e7cc5b5f96f12f58c86eb69fd17b2c5d97869ccb710bff3e397a03b151de88ecb98635dd1b232574027157ffcbbc9032cbc16aecf56eafb9900d8b9a844dd8a0ac711cebd5637ef1587d3118db70481bf697484768641d0854fea449d22ae515049adf81708e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4b71de800c9c2b7e025ffc2fa81666c4520caf9af77633136563c9d3dfbb8819137e45f56f5fb25efc0394c8083ebd6e61f99f852cda70b1435ded455de541a232ba17516cc3dfd42d85ccdaf13d922966367d22e656331a94e955745d6b62a3311b11705d4e0bed54b1c34046fbe738303756478466e36efff755caeffc032;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d316b2054f869ef2b75ac32a8b6c5f3fbac8bd226ac6b58236d32eb63a1658e8c1e46881170daff47007bcf29e85a25cca045dcd26e7fb46fe92b28eca3b3c0bcfa6903416b096857220bc65d302d8f24d95f8c0842549a6b9e29cb0c9738c93e113e92b56fa717452b49e8714d7d63ea91ece669620a664778fba492301e58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf49994d4e6b161a1835962d1e1f09ff3b159b69c78490b29cdaddba0960ee5b37f2d0ec7f5c52a5ab950b7eaad2397efaeb0fdd5a8ef7ac210ee0e06ecbe1b53d89f98169da936a703dc8d81aceaea43403da377556d6b782fc78cd2de19ff6182270bc1390c9a627a3fb75059ed960a51a42cae7c032a429c5dc64e85d0fdcd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d14a6307f897ab8a3774dc0d4e2cb18e3f87d22387e1a65b1e5539699d456687604adea8d95adf97532965f3d8365db3b276b0c9842a24acd85eecde7164356f5dfa3f9582c4558ac7138d8cb622f1aa2da86b1077d711ff8b6c67ae633f2f2805658c4910e2e396bdfbd345a3201bf0d43859b34691a29c511b05d30316e88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he33dc129aade676ffd0100b431d111088cd30545244573c65630effdfa8d798e262610d385bf844daac8382c5e7882c1547a061fd93ca81538e4afd21428bb34bfd23f920a6a579ef56cfb591a66493b91c52fb716a13a764b31f8e7701753c4e26f51bd50d020be942c425d58f00f0dc200b4a43e45352388a50118a6ece6b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he84979febca86d4d4a53c972623c40db7df369006661f1bffd3d47510ef8ea14cc31f0d2a337f5c2869607a32e291de7fd6da3abc58cd74b40fb87660b86e4d2a4594263a3d90d64ede01c4fbf43b9b630891460e0aad13faaf12411a939d4f2ee874809143f2af56182b0f131f883129a00281fa0fa12331e676a351d3c6454;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca701c1e18f7cf46154ef59eea526063e3dd749d33a646a582d67d43a9fb9fc4701ba1325ecc074050122a0d8155b40f98f70a99ee3e0883a599900d43f03ea6abbc952dc356f3d2f47d968b27aa85f07074106c56796e918b87b6c3938594c9cfcd92acd5c1bc3a30d78620fd183e464ad5b1d6aa3e95cc96e82154ea49ceae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ebb3e610dd40e2633d05075972b28c32bda5302441095583347d105d92adccf97937323e37de0e5f93c1d3eaa364fdcaa9e53ecf8269330798d559b81659280750cafaa2da63efd2c279016cbe4ddcda6c41fc7cde8a7624f59485cd58ec2cb6d7e983aabc729a6b233b421862e82bdf18152ba23a8a41380ab03c3dc1443ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f45b72756a7f80bfc00a9b6f080f54e643f55d724fd285ef1f6b1dd62d12f82bc46b279302cec8dc3473c80a9e0593079e8f291ecb59a99a4264bbd1da2282006cad764fd7e9e883adb1eb99993a9680be341432e5731f9f1759202c32213beda92b6fc46d75335bb4d2d8e20df89971343b4a1768a37b9dd09eb952a3a4665;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5181e98bd6aed67b1d8fbeba5f44f7d53ed22cea62db3ad89cb46bdbaf5450d43fd9d94b3435168189ce9da1f7f08884f626ec177d9a0396588bdea9feb954eb6622852389de778131248e7591aa6168cc70fb1376fe2f6f608bf55c84c900e3a6c30c1645be8e4a709ce952b91d969b43c849035d9ddfeaa2dbc0ce4bfb05f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d573607722709bf666e1cf06d9c1afc7b3f322d04a433ed2115c471157c167c2eab21710eea4236209ed510f57b909175e22802dd4d07ff04b364a47a79ffff60899c400f653c99968dde709e0bdbdf19c1b44bdfc074a3c5de7949294a779c8f74e939625858102f51092392fd6983cde23ff981afc907eec7a19046509c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h896bc5b27c100e1e7e5738db7b1e076642bb48b26e8eebc81f750207ddf5ddeb50d8255cc3a005c73de27667824a588c009ff972cc273ab19224b79840d259152200911e8b53d130e22ed5fdd534fea132f6d61352607cba68150684b51f50f4576b96a93d2426a9e498f15580935fb2e2bfb79e62bec149bf233d17544ec4e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff95b23af62b50da04bb898fe4d2d86b6a1a6340b9b80e9774e6236cee67d9eb0434de1f60d567e3f87e532edc410fc3fc9921d9c7bfed6c6b6eb2d7571ab26755df5ece051f5a050b132b7f835f0093ebcd476514be1ba8921e332d78466db71c42a3ce487767b838cd09e053575e04139f706b8d194b46b6259a2cafb446a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4d2ac0f02b10ae3d3a94ed40a31396f08797d4c94882b566e2028068d894bcb90d899cbf99ee44ba2c8ad730a29a6e97676567196ef07e1b15e0357c685505ada68a04555b2e7f06b77142634ff5550c9788097c4218091e50cb842bff70de630663014b34cd83fcc0d5dfdb94ef02aa097a783e38ab1017e6e97c8517023d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46bb40bd25e3537fde0505f24d720a60c96074377db29412cd5038cc6112af4d0f6a96fa6e26af51ff98b11291b8fc12c70f06d20533431aff6eeb4123ffdef76b74de28c48669cfb38aa16c82454247b7abb222ed3be09a21690b057d3c0ba2059d85ce2b62aa8d50e9b552a7e5c7535862429eeff357002a454cd64c7579de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he525e99753a5f0b305e978334df2432fa40653dff0d2a9ff14a3b860d4b5fab7936484ca680fd05090fee4d321ac93e73f56a50441d1cd3f5ad95ecb1936fec5b52b82785acf4cbe3d26c58ba3da3ac26dadb39570cffac91b266ea5cd1511727f755194dcef898c379c8e4d06bed334df81e12e49cfb15acca0b0d6bf5edc21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ec0595c0254e4a197f984a76399d8fd6d7b60976f527e72d2de031160ca228a3cbd48649cad2ed4a3e176452967c92ba1b5e159bc0e8a003d4a69ea6d3b2552b40bfaf7b60303a4936b23b878c47a07e2a3326afebd89144bb56d54a3b216c6178416a6ac164c6c7ed4e18c35150de636ae4878454b2547897562abb50a6d2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc56f66019bcb971c6e0abe6879a41e428f082341e971f4ce4c5b5f5dd4a027d475137704206d3596572c68cab8bd9f63c28d34f8be5e1dbd2dfa6e52868a5de67b767b64fc76c298a7214f7a61dd30a479aba9437a5c9d1b2712d8553bc19ae481b67da1f04b16b9d3e36bb0c0c356e6f9b1c0d886663d7719e2aa963f0269ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dad117c100c0a11575e533556b41db7a9bf4a9843fb136a6655d607bff49a542d505737031060eee3317220086faecb15e99400380889a9662ee8eaf483a1b2dd68adeaaa7652f348e91454f710e95ac7241eb753c71945a0b37d57c3ced53abed50ac1165ced5165ae9d4a04e0bf0a21eeb1c40ae972ed637cb61f8bbaff4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c9d4d0edbfff2dd7c60abc29d1a75f612222b6d68f4ad26f716a2f1babd1a246f5040767480a4e16cd8cc21a5e977349daa6e3a80e91ecf286826259a2b01e328ca6b87221afee6e36fed6b5acd8f9fe16c4d5deba9ef95785e5a36e91256102ef8714826654fc9775a1f5c786123c182895d837bec13746d094419096e0daf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1aa7c3114e9afeff8c997cb2d667cee11ef332b2bc908bb2cbed862b52667265318545698e13c65fe6730491ff41b3edd54b74da14f1d871944d152efad1d2fc6324b983882a3748a3cfab38b03f3b730c68cd7d69650a501a4d57bd7dffe16d23b1440e08962539e75af0c7e5cac63f9fd44798d3b29787398c7d27dc59ef3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h900f374db8b0c968eef7c5ee7ac5c8cb7069a67f9e7edaadece72d41c748c118266b27090540fc055df022c61cd4bf3d5843aab50438476535fec0ae021be9fa83b2bc43a74530f1b9704abdc2c431e35a56a965ae012deb9bea9ea75f79018cff8780bbc6848b2a618771a434c92fc0414aa6b9c43e1c3f42403d1c236a8b85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67208578b516884c3332bf13d502e30c941d0350f61484194703860f04f9323c777ecf9c3b7c077e13fbc748ea7d509d690a6eb2b5dbae4079f9b6cd7bf85d2a926ed22f61de74f7de36d5dad5c3a6b7e7d5fb6e56decbb9af5e95d53bb51ab454a57c996719db93d61b61f71022d79f2c313163d07096a5843d148708fe7684;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d654d1584477ad9b3e1b178ec631a605b4c0b2107b895e0bd7abae4011c04e3117c8ffff9b9abecc9bd638d392511781f0a7ce56530f8cf30edb9710adbc233cc15efbe3af6ced0312643f41467a85959a81862c3e51f3ccb420706a08c01c398b6d107cdcc9e9c9cf791fd2213b09ee8afd5651244608e2418d17b952873c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49cdd9efcda50bb73dc4aedce40d2eff700d958faad900635b432b8d4af58b22e81615d788665875c64dd6fb1dcefffc374f77f55eda3cd4e5a34b1f98c8163ba7678017646526cbf86692d6bce01af17597b0e22e0ed8dbb29186d6f0c0140e0deaacaf59ce5225ec3c677451967e5b1b4afd88dfabdae5d57c5ece5cfd7afe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7469d29432f59b8f91fd781f7ef573c2c752591a4eab4581050aed4a4bb9bea9ea325559730b09521e2fcd8aaf21cba7090c0b6da0ba1d26cd6dbce0643a1de57d486bcf41d282ab51d25b26a9dcd27b99711b38ef21a4a00abe505d9e65581ba96c8879ccba5b09017d4e0c9bdfac1ced0d199ac212d1c9ec44b052c22e97df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97490a80490e95e2d427b3691a8d6b5466fb2094128c4290d2bd35c0bad80550e58d83878717ca773a975b7188b233d133ef520138552cc60e6c68e1e4ab08848bcefdf2bb48ac65300d6f0dea5a2981b82a197027ed2f59181b2877b244ad6af7ace486b13e0ae2ecffafea6823161954fff58376433a8ee2e4aed886458588;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41d3bb33744875ab2e0fe8d8a328ab9ce2b0a33f246da1f12e9139294e43affe477fe2ea82ad49cde2b903750e8f3561966fda5684d6ed4c4e2ed7c1b58673a944d0bdfba1e99f483d996e4b722026dea907f60fc667c07695e1ecf2b791507e7a018dae9d0ffa1d37195564c7e4b81855e862ea2e0301c6792071de43c950b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd48b95cb50a62edda26ccd2cf5a87fcc04c8bb1a303ad4c56df309d6bcb8fafbceb636d421a66125c072179b036b46908a8a944e21a4df87c20e7c4e01229005992fcba4bcc71242a3444ada283e0ff632f9b807c92236a2f3ff226a4298a85d1a0099cdc86f09a014f35041eeb7a7964c7ea23fe681935bdec74a444e2fc3c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25eeb44f54e439b2ff45301d7e8e559fbf9631f140efc07790891aa04a829863f7883a3beba39338ad7a9408b87a785c0add4c6c324c5169fe0b94cb020f9272073255fde2e2ab06ab77bd6d01b70126cb66a9d7d1852ba60e87f0ee6cff7816fd6780026c1c0d6c971d1b1ccc77393ffb66bb5fc0ae3b243edd6bcbf61382a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79396a2ab8c549a25e5644d238f013852d85bd1877fbc7c060c5a09e7d5a49c7f5e688802c91950f3a14bc7779b7750a626731867ca2a30144471b56ca34107af7207656d251a8265a2ca3221c3233ed7e45f7dcc85c423860a5dbbc197fa55d31cdea5582cd609975e3a47b791da9d555ec3f35cbbf5f959cff4aa030f4811f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b1b0ca494d15b74ee22acdee742ad23a68305eb97005767c1afc06866628f304effdfa8389c96625b33568f26ff6702ec58d84e010940aa863a8fe9b534e24f4ac5574bd464a7b950516329ff2b75fef74d803819d95c3b86c813ed35d9568eb14fb80a4c2ccb583569691d83a794a5453dc1e68996cc14077e26ed28526a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb2287437144aa764bdff69a16b2ca3acb4273ea2c9640aec46649bab92d6b8d31f6a605ac72830064232371e0ceba12279f3b6df82374ac473f94794b69228f0739640a21a60dc4ffb45df93c9ff80b6bf765881641581bac448a2dc68ae5fb708992e647feb81b7d9093ccc0e00292b3b98e5a53262c3596b3982438a6babe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6858e1906805cc8c7799158c64d5e886d6304bd13d84c2fd6b40b3e4f370c6684716c6bc9c3c69c024bd1bd3d0df03a171d0b446841c7c2048a1dee2e15343799d5a8577e341957c10e24b42c263cbc40f5ba1e34869d41983a06e57c6dbcc9e61de759d18c189115374669403553b421259b5e888009dec47c0a33ade786a81;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h768bf05ce9dae75331f9117a1a8d2d2bc80c88914c8d51d2832ff1916c9d941a7bf11c78983727cb08a5fd24d969dd8470343665790b52498d9140d7aa415b021b3cce61560d73b924b0bc5ede1a4c75e2d69eafd0b11cbc1962c4ff5b63b312cef80cb3be2ccff8dd703a30a4506964f968b754061bc3409bc20859fc1fb863;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c6e541161323e3630407670fba9cdbda23ceb03295f35afd3965db4d785308500e9e2be508b06b4707b6718b5ace3b68afd4aa44813c3fa581636659a4792d250613c8b5542366b118cf420ce3a441ad2871b59eb411daa8c5f1cfb1d324a0dda9bff96ece8fae07c49e13be0fb43ccf3757d8fab2da1285fb8257b55ca4686;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bfd6c6d823d4625120476452e4eb41061e769c2103ce5468626a848e6e5c541858e720c2faa519020a8f5b85e01ec8dbb9500fe3b2b6ea0a48d2ab4ec199f40fc9b3d49994f83956e9194939f05210ad90729d886a72428fde718f946fc01be0d975e8e583fb6ab8094ab1add89b4d79d5b9c2a1d39635035067c92d768a23e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2c22ed3ace52e8384ed05043f2e28c42521684f0f548ee1794eb9919f5dcebb8a8b84f562538b77b3f9c40abcd5f8069012351a6b7c19e96bc5af580e85a8b0013be3b651893953db48987939c07dd67016189272c05becf3f210106824d4ee2192094679028806097e6a8310ddff66dada8f9e92bac8d3d753d9785fe076f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11d4910918745b2a1184a4db207e1132147cbd350e012e6e32979f4d20be7ce6b4b9fac93a195765d408912fbd0a8bf59278c81715e204bf05eb0cdf7a25c5252ba6467b717da4aebc64a57578325d70d92b815bf5351581b0ebb3534614137af8e6faaec58944fcaa29cfdca12b4df3ce5d6c1486f914065cc12130eb26f3d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a11bbc8dee3db477b847686b4807110d6a99e31b97c1347318da2b6e3ca4d94084e97769e752ba96e1c7539dcf7ee841dfa6891602d13cac5ab8434dbae76922c63793083b19ab0168ca3a74c32775ce1a7b04b6147a5835fa24d9c47d3dd52b268143b5a7964fbd37ef002041f8222e906866cb3abe14ad43076c98a4669b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28c499a8f1668f676157a0a927f8901fd5f965b83b3f31886f561d9a2cc076d3062836873f0b7ad330b2bc3826d2b9b1ee518206b5bd262ac855dd5ae7668a8d5c5280facfabaafec41acd795baa0bb29a9f6c8920fdda7024ab6611891e572b4e9d83a444d810618091426fd15c9a150c78d90f4c54a13e0b517a3e01cfb1e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h819e4f7437ef8bc71ec231138b90a07c35d52c2497862615532d6d3361babd512602ba45f65175858972abaa076a4a511eac3f38e0f3d4df766316aa67fecebbe77b642b0bda50ec6d4a6d84a423e5dc234e7708c37b09b06ca86537dd895d9b94a3ef3e71715e0eacbfeeede8032e63f9bc8afc1c54c62930c4314df86eb5ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eed6b55865b9da85e9c878596814d44572af883d6c6ec7bc823a5fd96a6fcb3749953943ef8c0f7a19b9914f33f1341710dde5cecdb83f84921d012f180774babb0ab939da035e2fd532fe5278fec6047aebeaed0122bb7094f3a6ead6a07dcba46c4cefe912bfe4bf6bcfcf24cf884b080c9b5ceb091f2f56bb218de5f38a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7571997eb71824756043e3f07aa79014cf162df485f75d998644491ad4287a187eb270ca58e865db728d5452a421eecfe38454ac7d9731ad23ec5fcce36bba81a2e874e05da8aaab2de02a2412c610cb7598f980c0d0bdf5dd95ea2b351cd4974a093fa6adb76935e386efd800469562f4c5b5932b5c7ea519607592b5ce3cad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf15c08280e81e0738e1a585acd5b3659e73eee270adc092cd0c77c2d7e25aa56119d06dbf4bf626d3800099f2f3d5ced96a1046b3f6df7cfdc821912b74d123c4d5b1a9c1752fe5706c2aff83994dab78be09f3a534d35f7c9d7900ecbaa142da46395c7f8c2f6912074dbc652b1b29d66a7a72c84b6e85844c21da724741033;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfffbd91cdaf665bff9555258210c27caa4dd25e63c9bf00b23e28216902da18ddddf4f103c74daafd067c99a43f9b3a1c944d7df5372be05b689c8a1a78ed16d7df3cf76109552a035d41a82ff55bc6faabd79f583f3ce3556e5760b19c92fde7fa9bedc4aa7351e5b6476d99387f08b4a9f7fd7b8478d1df04b93846ca89fb1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d5ddb810a1a453a7b466ae5e3d70e75f9ed2baeb70ff7e342d0cbac4aa3851add921d9593a55056edf5021b8e1616341e40e55409870872698dbaf78fb218652e7c804a00ebf213f4c48ea7673ca33534a266cdbfdd89200a37809805906af6fca64cb01a9f27340fd917d8d000c1661533d7cd384c4c83d5fdc28d5dbb898e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33244c4e60202c20a8e3854e1aac41ea97c25cb3103d5479425181148273e54ad58770385cfa37860ab09e903920f0ad2e4c8b611ba11f67e4de5a61326d82af2c0c35c201e1d9b8a25a045362c1d65df8fb2f0235acf9397872ce198e19b54d1f8f9fd8b32623bddac6933ace8794c9003cf193af37e4e98ba99118c5a3a1a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h509be0f7e53956c5eb75fb0d98d35bc6f921789d23f2975d8e4271e4a39c16c5da427c3430849fb25d081b74c0c755074eb7cef85009469bab27cc2760618044b0a23661a51883e480b2b889bf72295135dd53e4651064bdecf14656534a7c16c92ebc2c2b71227b45c5ae824e7bd6f11f30982a5e815ffe02e770ab3b676536;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb05c68521edab44a233cda3ba0c26c6001da6d32a15890eb96d4444b12cddc6b8d586bc39b2b836b95bcb8e279862d9d22414305e34166782c0eec5f9e1c244473429769a3d982c637b167c02a4a3b2918cdb264abfd611df1b37999cfd89664e613730629119bad183480ccd77c06e9a9b79f4b259aaea394d9e7510aaeab5a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb7dada6f566142630445ebcfb992deaf21a2d78dc5ba16f9689b5f2d6ca80468c53b9715686e260469e9249abcc1f6857aa52e4006757630abe6f442ee336b30969b9c7d4d4df62e32a4fb4da3ee7a8144d032f67f3492bd7d8c9efaa4f2b5ddfaf500e8aec23b37dc2ca5a3c765f02ae4e2efa6981594d9d7c6a3a064cc6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha16cbb3e1fd83709ed4e66fbdf96c2de4af9331c707591ae1764ad7181e64008a753e7bebd52f22c8984bf548c41b363c1e45e659fbf4566ee649e909ea3a447df0ec5bb48950c858ad34c2fafb1a11beeb4e85d90cdac5ca34cbb2283b9715b851167632bcee7965fd0c5a99a48b95258e28c3336175c4f5903e7930936ad0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c2fa6ffb5dd32c6a3c06a2842042db4cfed6990ab56d6007b583bf755a23954b9c1e68c4919ae4629c5176bba4a874957fe53333ed5d664c3a0d97631eb0194eb5f2ac76d4b6481aa29d4e576b86c9adb398ba96e5a66c95cb6d15521307d4ad43d951b866d112ef42ea9727510cb22b4e9b87c66c9d08d270d9f6d9378e403;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacdf3a6cc058e763d64b68cd154f9b617c11619185afe5088d80f9beb24e94644d7aba3864457be2fd3e852b24dd0876881f41b5bc805134e80add1527c8f14de667dad699335fa46874e9da735b110d8cca443bde1eb4f00455f772ea948fd74d698b77f112380f426b47d1b4c474fb77e154a4710835046ca04b96f8cdff99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h522201ed1c5c61e52e189a504c185c8a9ae37305df2ba8d1f8ce83e70e4f6935aa80c2d03498327a47165dcae7d7ebd9373711b29739b6c8ad07bb1803c8499c1e2fc4e4873f3c77911f909f3a6fdb8228b7ffaf05238cbb92b13db14a9372519005ac415ea6708242f8ece43a96c8949e285e3fb04409cd17bb23194a8380a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c3dc7cac283a585300989c8e228931920ec28cf9d59919c76dd6872186e8e2b2cc4c61466b7bd3ad700b3cfdd127ab599178aaf6dc5b6eec53d85369cef43d1c78bef7de784b83df8e6c535a67aa0fddb62707acf4341bdc35eaf997aae91470f6c2035c724f3f65119d5f8fc388ca08c488aa91b6eaa71e3c14607d7229eee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e8e5695cc774eb5ad8866f52d8677c4a4d48b3e50c1aea8426a1aac9370faaee86da6cd0b56bf0d10ac80049afd85ac99ad9780f503ab2842a84bbfde8c7d69e8cebcde2b5c2a0c5eb830e08d26e890999717595930549e7deaa63119a9fcfe470c578c8462509ceca110ad1204732406c36a0b699646c026df75aaeee3c7cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19037196e0facff8adfe1e517510b59b46a10e515c675bfb5ae2a9b4eb141fb7915d5021760de9b94cdee0659b54ec32088a7735a3eafd963f8f70b49c7a70c79736061d3e9dd07aff4ef8c7e42c49799d56d4b016eead07ff43f05c919348420fb7dd1ffa22ae1d3c6cc87f873ac5f5df8ed242c1b9e02c68591b83a8bd50d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6754449940bc5fd54a9945f274e9eb29c453c199633f3cdfb13b1eb9e118c96ef3a3aa6f41576937672595a59010d10c464b57d19d3a89e94552e8de19f98ab6d38d519e77da64160d3a154bb8d437bac4206c1665a63f13a2de92bac4ebdfc99cfa31cad1f780ea323bc076998447927b23f7280943d98805d3909e806ec3b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc180f8948161e49fc09909f630b0396df13115b93b865ffdd6e6829ec85a883f17afb295d3b12c42af04604649849efb12b761967f9df9e7a3858205eb322a23e2a1f5adb40a2d86555daeb0bae90f2c5110aca50e2d84c65de8a65b93d3aa917f6b81fee593f53f0a06d19ba131ee4678f1b251669e207770fe47e3801b50e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90eeec7711f1134b39624949a341e74c18c1a747ccbf1e839ea4f8d42f2831eec59c66ba157077cd8b0f200d9f809595a885dc4fb8c142ce6d475a092cffd0155babfc989cea1137dd7b5dfb46e5636f6cdee725dbeb4c5aff70b932cc0d98082fe50dd2a765ab5c089306351b22c59fe33c7d733ee25aadf25eaaf0fe939225;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99cf79107194cb3692e89be9ef6b98de2f2534a559e2e5412b8ebd0a1d2e55232d7aa44276a882ead23828cf52d8ae488736cc69ef0ff61c92996db1a205ef263028c6f1f6f8e29e9369721f458a4bc7157e538f7d2b1a1dce247d4a2a6158a04ac0f170833b7d0477371e552ec22e88be50433718ba26b6153534dd20971c8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc237e679cd860ea26006ddc9f7af25d22688847d80ba387c9580422731915b72c3ebee42116c0ff26085fa0599da555e2647586a4861a6b9c7a25472222610142f5897228ca5ecae578b30a31c57d1db0b692a3ecd9803e7b24dba75ea72c20ff005bde7e7449c6c928ada7922f64ebb8134de25ec6249441762c5bf9197117f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca5dcdc2a3a084b4a16c44db8e92dc6fc8d35f8af0a2a324f50bf98b5b5923d14d571b89ff4391d98b04b92b2467f4496ef8728c3148478c41d8bfc0c84433e029ae7e26985d39b40a58c9d8ed612fa7e8b63a6c87a2ff5896a5802108d41648e6e1a4170e240d4de4e343c4e50a322b76a454c75e2c79a710fe94a943259b93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95762c5e8d1682bc50ad19cdbcb612ec0ec5c89a7d89aae869ff395862484ae96b692c18a1b72b27f916f0a74eab181b4a051f7e276a910e6dd77c76d64fc22d5b8c436493d77da92b47de17a4c4a6195255131e1c98326030f62d07dc23e1db6404aa4ac54c0cd876610d51ee7b64910ab84073bd740e45daeffe5916a7ad85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3872a38b6c64ae3cd7d8fc2c0990a3097fb8701ab31fe63f3a66e942854b6530ee2e2738d8365e6df10926973e9e889fbec6511064178486eabd369a26b9ac2ddd3d37c1fbdd3b962d048a3266ef88fc31783f6d9b1eb485a0cbad145ac1627a63972ef309ee8a1cd9fcab5a2c4f8b98cd6f01413e1c62e84af860f7ddbae92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9275312f0a524c480df90a69c7487dc840ee665f310241110da9515f9d28aa8776da398444694546db2aef3ca99871ff6f4dbaf53b869155f04d97b507c86815d8e1e317289d9eaf9df41150726da2ff3a0baf4b956319516ba9ae310c6b409dd9771e15907ec1d763322d1b7ee2052b16de8fa9a31777da5ba997a1b54b99a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7691e120f64be6502c2472f2a7118397d286f0514c4370bb7c0001af380621fe6d386bc0dd9b069f1e7a59d50c20abcb90a4d8b93b0b0a256c5f052901762723603ef8427943547e702757f0f91664e2239d9447a8c33f8f30f22a7e3c460f3ce6554750c587ce79b0259e80f8e564a4eb29323884809b3b188b814548ec934;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8786ab657c7075452c4a6a6460184ca7a2ac9483bc86fc460cdd34a1d0f65f6a468b009c201fbebbff3e4c932d3e6765afe2b44e390cd28c30be8c4c8a25294aef2b69a8cb3976f36696aedc7643a27b2e002480615d0327182e195e4137cf6ff1f8f5d14dceb5d5ee68a43eb3f0197a25e27f9771adb0705653ed1b6e4f24a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5af2ad1f4900c1af33b6465aad2f6ddca0c2e7f0f26864102f5bf8ef1146d195b8a0e4c25858e9ea0ae65cc7c9d593d24792a777023ba1f7e14285756efecefa2b44ad09928e2345ca05f42ecdd6a622b6f0a7d8c53eea2f0a7b15c4891464ca359fa26afa43fc749534f4b113b8b6bf58da863ba100e374966c5591fff7687;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e59f0473485875d161b797988f198254ea66d1ba912b11251b0bb1b6ea6b6a50a006e3cbd9a70d2e54226e9f780c3028de11a4f70720ad47c89378ce35e4496f602555db7464a9f15140cd47c6748d9b670485ad5bffdc66fefd3773a989e47a12c68f8293c40bbe7cb17460f0170f9a27b89606477b401aef57998ce6685b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha83a460510753587bd0e54cf0474abb6ee8a11db8099df2181076e052bb2a80aaa2cdc9c15bcf1f973fdb6243c32755559ff0ec1430c4281b811541327d65bab1c09b98dd0aa51a4746d5d594cea4c6b343ae0cd00465a0ae4d96923492495a9076693ec408a23d6a495010eb6fdedb9d68cf2e5db89851e9fd18ddd7390dfab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffb74d3e6e3743b71b933fd9c65cca64e6551e1253a35a20217c7ce1a8ce3dcb62e01f5f29e68dafb3bc4d97de2b4da07db5bab88e4fca41571d9a1c5f55dccbfdb609cfeed1609e2a0e7723f009f9567940cf397ba79b23252a5977b7c565258709ad6b59c3040eeab600d0fe6b14088af5ed4ea7bb48384d72b926d5ddb874;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf25f5b91bdd45942e66f6ccd8be2beeb4aa74070828aa662423e93035a973755503132a2d411c15e5896410192c69c403fccc8ae41899ef3930364885decf548ef1b0c8712cfbe5867a2e207b0bcc6313ebd0c7153328a2c5b76c4afd9276e1d45a562e3bbbaad6431c74da91855695d4bc9ae6de6f82d4fa94c498aa26040af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9352d0ca26f3da0972f2a83979d961a3ef11c023eeb461914444702296998d40b2edcaefd2145b104bbef5663f61435d9687c19e5fd56cce682124f60b666e2c7273f330c59d723f5ccf2029665adcea761f47cb5b3f6b1d673bb5837db55978df7f395dfba9324ac66fad100c8b6284ba87aed8848cfcc06cc6f6fa618ecf49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ebc08fd78520ad1d488b2fbb15f21cfbf51176ca1fc48e46c53c8e482a7ea30c9f58cae4371a77a2bb731b39eec5827b45e9073f0019789a66d9881a2a2076695dc065034b5ab7f4d4fb3a8ea81df50e75d47ac519afd3bed658d591b094fa54fe5330788a70eea96bfec4de65270b06fe56f6f1970e4c8d67469e3acea771b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he39abb8f6cf6af7d07a632cd4e97c00c1d6538d46927539d72cc87c4a484ba6aee057bea45a4bc8e0b277528d5b25b482f9ae8f3db8e336a453cd15d35db29b52411fe4857d46a62421f31c5bbb0da22127632a88352b03d39de55176951241a223fe395f7fff75486a93ed35965a61e925f5386bad74e7b2c9a1dbc87f995eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9fdc5647651a8f0e8373ddcf9e79b2697c1c241e9395eb9af3caa474649b39120e4c41eb09f46a5d22a10b0d9bbadad5253518ac3b3c4cb2c1c43a58dcc672baf5344cb8ea0b264a970e0d10e2eaafe7481ef3f2d349cd2c5577b55faf314b3c45bb87459aec332e6f10504cf8f94d0046cb37005adb765695cc70c81096e37;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ccbfe77d817c16ecb898ba71da20232a452aeee1fa3bffb195277735f3e9e957a74eaf56ac0b325a6938257e22e5847e9cbed0b0ffd2ba78225472fe339e4fc556b7456f03af34d8a2bd7ff827ebfeea87ab1660b4d24712f4b549e4fb56178dfd086883ceea1f9dfb46de279bf645097b18017c71ffce420345ba6cd9c94c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9c78c78df2795c02d44b7fcea91032bd260255504801da33d0571601d42a171d5aa6216c26e11f73173e903e8304d6dcd5f3a5cd4555f2fb548bfdfacabbf362456c90c442d9f4e2ef13bb50ac6331ef06d32e4d226c6368e55638333ada259960a05e71f30b08eb170a82bcf18ac4dbbb1cc0886435bb7340c52cd98e57daf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8241df1f54eedb3c1e069f6026a6f04c566c20f37555062810a37e5722508b528c1de47400423725f24e174713e473d470ee69253948e5c41cd8d53beca6fa76e250a23815f9b7ec3b750ba90b927d2731f01942e0921fd820a29f5f5e9df717b9dd990fa39a3c58c0ca44a4a35d805031c09ad0a8850df8b0efea198a8c7ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46d01fe6fe31dcc22f7460e9e78ecd5630b82b823a7bbb19db7e1c0c035fb78c4530207d0437c7be5090738dc8bd50f973bd74a0a44edce0b77b46bb568fdec0259a079719e44e912156184e31ee9f0bdf09cc9bdd52ec87594730036d8272520589e5b043d268ab4e61810964f4f1081bf82a1fd17284509f925b4bce341eb5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14fe2b5290614869338d846c64ae6f99964f6bf0db3b5416914b08646c3c995da02554c43c83492fbfbec7defcea34a2caa28b48eddcd58d96ebaee00501974f82669c9858ba42ae3618a4a8a7a59d2cb1f9407d187ef9bd6218cc0c07e3b7c6068daa5ba1c719978f566efadc31117d445ad74eed17acfde52344960358efdc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b8783c0fe274e8bc1420a0f0d6636689bd5d7d5973849acbe0484802917044ff9694a82b69dd0e0f1a0d7b1a110ba20311e90924b8781de7bf0e6c5e2fec05921db06cf6ec03147a285f3688d01d13b93e19cb2d9137fa8340524fca51d43593c12574fce4cc0c2d950780b036a731bb585a0fbf51ed9ed96ed3dbd1ba2f4f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31f3b1f06edf8b18bd89b529c4f7276ab6d5c43552a54b8e6ad873e37e173cb39747c38f2cc990213ecacb221d3861f3e2b07f5ec665c77f32484aa24cb707cbb4408014b500f0b1c9ab69c903bf4804f6a7d452988616b8816e095dd2fa379e290afa154f9a42e8296e8bdd7a059b68c9444b01590f2a4c834a3ca0f9d2be0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h109286f59596ee1b840dd35d6f206de316b9d3f95a52984d5f7ab3cb5e6e5b132116023563cf12bef2db1355e2f810e489d041c63e50b9ffb168ca159c1dff83bce1e3713c88850e6cb69d6b1af7c7b329336a23470df2c42f2eb20a07e5d40451926efbe8a519902bb3c54f38aed15f42354a0680fa2f251a61dc82aea7ba85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8562a0d6f8a5bd88edd534ce5acfc687dba95e43ebaae2b298dbad345211928d5b5ec4bf70c5572377dd1464632d569f4b1521ef7cd1ddc1711b7754499bc90c5eaeca2a7b61e1d73cebbd047f0a914eca109d7a34e7808c550092ba3a2e073efbd8e72a92e49dc4d89c7ee2a25d2209096a2c914362f824e99a524da57ab010;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d76235bb6859d8dfd40e76a08299cc5d325a81b0434c18d0087c7d269159735d8f729c9507d810c41db4138f92ade962d2b6352190422a79ca3879e11870fdd9364037011e63dc7bf479b52f0e872456f72dfb186461f6d14a79f5dd5ee366781afe7698ec318e1e30c12665e9e6e0ccc41e97a93bedc0c590c2062df460a52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb316a6fbcba402f6cb3e67147033aaabe200f28e7dde15647b918643913e69b3597f24ad3516c7a3323118ec03f943be7a3b29e779867950ff539f7bbd81ec0b06b392f054bcc483c048da5b7dba569a149bfb8ddf555c2d009f48172ceba233ae3dee3732dc4581a5fec0d63e5d4f57bdfa3204efebba0c51b5e92eabfb49a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h139f85ad2a03b18f0faf7ddd24762897574c8fd684c67f5a766a7e8d0c6638a93fac5489911ef514b9b8ddc9b6f58bbf26b37cb8d23061d949198d2b70926a85524546d83cad1641ba7daaf5cefe353d169290af13d03917f0b976c68914a98c80f53ab836c6d9dc7d5f753ee7a4b7d5fa51c87f72b78bb250d0070247976653;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d2607cb168f647c5d8df63932a9d542b835d491ebd5d011ff618954c60dbc82dcf6948f9739a5738b083ebd47035c3ccbafa50201ebd6fdc854526957eef720cfec0b13972fbf3d958e9fd9501b881a72fdb7f0c1eb1ebb17b6e93490c694992482c25552fc7044049536f2e35502105e9375596ab1926c8b8b474a5dc77d2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcca1d65e5656cf8606f351b7ca75a94658527dee53a2f4b4d14474658f643a106efc7e0fa9e909e1b2eba95a96022feec6faf9b1e9b41f4ea0540f45c3f47451479fa35e595fa6e40e6f25bdce673d6fee91291150644d3ab7cec9d2bd1e488ffc2b010e971db3c4be7dcc90a472fbc5bd93a354dbadb3dfb1ade063fe8e834c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d5d47e846150d50feac2f440fac202e2fb9990d206a133230020aac1a2c501bc8b607b70bad12ca5b3b7470bb3dba128dbfd99c96d11b7e3ac08683e959cdf6482ee2f80b5ca4f20db085ba6737f21de1b9a456d5e2e52f7e0ab7259132e23fcb382e2984af25e171410458fc9c19bef8e2371d6d7f139420f47a15e7663bf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9345ae73a97b30903df074e9cd71485ecf847fac3c2d62d3436d0c454cdd926b104176e08de64cc1faf51df3f44645259025d145d56af0059ae7cd74843de9f9a65ba04486784ed9ffa935e44b088aff7b495f10c73a428eebc1ff230472a9bcd6ad287a235fc689c39a39d56b16d284be4353cc1ddef6017e90c574568567b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h709e172c044ac38ec9012a2ff5b75bec3977e19a06c13012cad441707d15ee5b010ea6425a4746ac4dedffd06a07b005667ebd86e1e94922f11599d6ae2d40747ce587eced0e72e5ec67b8e02e767f74b68b6b0930a4e92b271de93d27418c438a7d90912439c212eb06d852cbb704b5bd6b4d86d8635306d303b9e77fd1ab21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h263634f7e7824accf7c8599b760a945c1a357f75094f97166928c1b859e905ec70c0e78ef5968b28cf8db04ec88b52bf113695aa5199e54e80b3829be823c9b6047d2af98e3334350504ad3289f9b5a23d7404672210e5afb0bfab2f0e298e1c30eeba7c2f1e500a17494741801d7aa7364cddd34475e16029abf209165a5689;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaec19b7adc7ea18f4b7cc06b7b52ad6690bd1e969b2d4d76ef7e7c71a89c6e84d910230d8ab9dcd84086faf91b670e4b914b9d2e6312d04dfa036913ef0473341d4aced074a285b226a642f1e2b162d06613c5c8747cdf4d533cbd5602c0ae8d2eafc2dff4e8d1ba61d5e10702ddaf22cfb40f885e1f1000a57b89b8867303b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47be8cc05f11d78016fdcebd174e8bbb21cac8800830940fed7afb1a85543c7f8b28837cd439b970998907d65cd5a263f76ffb3ced0740124256a0c7c3a58b8a8a6120cb7b22d02a9a1b7c462997493f5a26cc525973f11ed615e82bddc4beeac9e6486d45477b5ac66d01fecedace741b00a87daa838a99246e85a3f794eb67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1adbf028ee8637517dd8ce050ed31a2a2f1f363b132d9083d7f099e1dd6432717fb5d88d3998ea162e9571cc5989d881bb93a0323326708ffc93fe9bb0ee17077f677bf31c3e2f3d65a8060d6bb58b5ffd079ea187131b8208f3e73b17ee1fa40f6dd653305a26bcee0a8be57e3d2e7ca18c43e62892d4bc25b226fb00767e27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54a25ef219c3937516a869ae182c39fdbc0025a7ba84c724ac01f933e339d4c5082297e8f2b6c839a695a1a88e452a8030b521064e59d3ad2c284f54cc3eb8fa882aee0847ed482ccca976fc5cf082672e4d4460d61565f0a9bcaf7923ad304a8029b56c2b415b78e5ad426e31fc881adb58603601e436f298cf86a570553538;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e36fa8b8bb607c8c9d1c3094dcfe5c736c3cdd8e931962d250a0fae7986bef85a0e32b37752db64b3321080709d13eaf7ce97c068cefe479b545ca42e3b7f096d7aad88744d45e8e9bd12444bb78b5c129c092624915ae6a3767287055101bbcdb8e62601fe8c9ae1dde5bd600f3c7de9bf3436e4414d8920eba2f81a5ad60a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19e484848bd5a8e915dece8f87e14c837504d13653e425a47c2036d5038568a8afbb666957234d119a766263d2b5be7c305570ce4865ae0f69e97f1625813191796fb37f4e8d108f228e3e86f131422be941a0c260b90ea702ab1e5e3951b47cb61684ff97e43919582e67614dc55816e13f85057f379f8cde154a8d78bbd93a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e595f8db7120dcc766ee5f78a2b6ee49b45775d095d8ceaaeada72095242815099aeb09b21d6caeca52f20245bc3c432f221d75859a85139f6095faff829543a789d5a07bbf68b285782db5ff5190323bc1b56431a0debf207f61ebcb4a17d6ba38dc208627019f7c48a5f715193f7fe153a304831f2d0b5ae450505fc98764;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ff18024ba549fac7d68c18bac46e6eafcc2c8e2df0f047d9b6a9de9e9e62371d2bcb95146aff7b8a606a17c9d86e63881629108c7d5e3159be7b6b3403ade67e4e935502488900e737f5dee679bda75a867738bc146dafa87fab3050e78e0becaa3872f978624b7f5ff9af8a3e7ee14ca31aa2f678f67e94a35ae4303f2da26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he33734d22fac19f4e03e07a961ae4dad6e47d8716b35f281aff9ed78e2a55b024f44cc6f8240abe6648e0a4fb8f5b252c367c24d2a17445000ff894ef8418f53244a72f10b6a732ee0e4182c81841f42360adb83433c198819b4935af94e927f4174b5056860549a20a9b5890b96fb220c63ac2eed3c02e4d1b1d32eff72821f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7a257cbb36a4da43f06bb951de353e433a3ebb681ddb75942f31290bb62ade89e5d011c7d11f47f35a6520b79f59fb35da1ffee8ac33bc530b6332b16971315ba47e04df7fa8d082ea52693d8cd298159f81897cd69384bc36f0b51256fc9e7abf209f43626e486e500fcc569fa3d2c110478d75a051b9aa8ae52839b225e44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6082371ffe70cad1b5f9bda9875cf782ecb1325a5dc2f3a52c3a7ec8800d78816286b4439fbbfa33f06a0a7cb953b68165cf65ff89a28ae482cfa1a2779dcd4660e3ae71055e20818ed49f4337715835ccffaa5c28310d97168f066c89555635f55fb8d931add1c097ea185f84efc1fd61ae3430bfd56542e3e957fab6a1370e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac289a2c353f6c16054b63235489048af46f164000c1af817b83974d0279b898f3e0dc750c9c7476599b2c5c210ff4954aa7f6dc8ee5e2bf07751a6d22dc0533662429d679d07da90ae83cea6352a174991adc63d096f45c7d172e7f097c1db853f83e40bdea86fb649b8627b1bbcbfa0de0e83330ecd413b2a758fe2208517;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebc5bf392fcf317add9dbf6ef9fc6c71daa9dfdf6e5529c865d3422fd5dbc54f91a56c355a00b647b6e3b768485a73563db78cd00fa68da8f6a36220cc0abeaa6afc798f129f68fdf7d12304f4dac963fe122bf5972ce415d80d13f05f9bcabf28eededdb761f3f00ae28f6f3aa81b074316345c719f8bbbdb4468ba3d64242d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf42d4f4103c0d750c886f5b6af030fde32e3fd0259acc39c999c032e465a4679e1c3296e008e2835c0f481dd59e3919fa6f37f4aa15f2bd584fe663ee2a4d90f4cb0e4ff517f167c5bcd855255ae644aefe891141967d05b8d4deaa2c1f02ae2963076177f38bdcf550295859c556ddc9503cea4b2042286ae76abd919ea13b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd0206435e56dbc40e14af71f9a12c7e9d22efa3bf642da9cffa301f502a54e1a3f48f5c963c8c2c51a8b83ddb20ee2b74ace73cd6f545a5caa620ed1c30c20e477d8da77f0b2d5c3eeb4fd747250eb6a6e157b58413a2c075c190bd0d444d5ff3e303c4856ab6679b48954d64c67e8c97927d1defa267064a32d2027710af0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c73b2eeabe39248a06c6ea1e146dc8ab5bb72062468019f3e5c2e50162ec06b4b402a7eead2d31272f6cb0378690f1a3917e909a44bc46f389f646e3932ed982d98a8aee1e5102fd8fd24f746be94f99c4a566fff7047d27a7a8991d3754e75769d9ec6ca6b300a16b5b74e25756361fb71e887f4e54596c626805e725c61dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef03619d33bb3f0554190830730c048cb6782411328627617ad8bf29643326116f7407571a656b4a671d4721ab1076c9f66cffa7e27c8da1d4c9f584be45841d7e43fa1e5e8dc2e7c1c3c7a1643547bf69197fa6f74f4dc6a6c3208cc20253e2c33f6b8eb990b503d0500ec14a5889e6c5cee12e1b0f0d7e2ce958f746d0832c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23b5d9196d44d458d6dbf5339dc493f2b33dcc2e5095030eb0b84ace55698369a2d4641b7ac806bd154be58d638dd4f67c8c8a4f4143c8ef6abd0d0587274cd985c9ca98611f44675c179f4e6faa0b3cf2125f55878fef9a615bb16d6154875d6e3e927dd8a8f3e3dca2ec954dec2c6055a17a776a9e0d6ffc795c61bb56e6b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c86254790a998eb9497b8ae5630833e7ca9541f92fb70a7e54318b770673305e377233a161b68b7162b65a4767bc914c83e470a8d4fdb49f5090bf0d742cdfbfdc805323385ba90f52e4583ed7c5c7b4e496ce07d0060b699dd6ea96363f02674240fe9e7386867b3fab4d6814fbc6aa0a6bcd9e850d64c5615c5f667b964ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h386f9125a8e0455ae2f58e165f786e6bd85002cf288fff683192c4e3189244f44612eca14c1f4b53c33615b7b27a607e1d523c3714596cec1448d0f2c6a5e09e9ae35c5fd4a1700406395680a7fdf4d9a1be1441abda813960063b3345fbfb52ca5bc63d8d51c2ddc70c195512aef62fcc12e6abd0bc2388df763eda31b86b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h798db777c9c89319519359bd6cb13e92e91875ca374c864e4e3f4193e850ad159c5488b5be96533b72b7e06df7b9da2294a57f6f1883f2aeff8bc37c3fbbe28415ff1280a215b908d8ce7dcfdc2dee96c278d237a5a599d60548f9d756ba7d0cc9c748a51a7242081411243486308fb011d9dbfa5f6099f882c139e7b4f6242d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae52cfeb2dac6dec1ccc5cd81736732ac471070e571498ab2955f7626b8a0269c735f8179743b020d72e3bd82fc2f32638268d5fbe45421dce318d8dad0ec88b0f80c2e1c9504fc14f9a34f31a3790a552948511e3d9060552e3f8cb0f167d34dc3fe98d401a1be00a86a6fb689b2e9e841e38f4b645f36eef7768e1ca368b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce8415a79b6350c078c41aa4ee61051097f8df5fe9ce2916ecae2724f767cccd8cc612a39ae772c4c5a80b9b16584573d3803615c5921ace4566157939d1ce815103903f69c09272e273626605b7135f772f83382b0ea1e7e233d9337b582ce78019db345b6b1664f2b24a1770d6aeffcea03db8dd58aaf7f9e3c894d2e1eea0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c803270fa0ba2131071b75e39b74e5aabf7ed5523ae16c6bedee85d7217c521abb9f34ae1306ed05649313010576ac1d8211e84f75f597b66494e1856d40dbdb2bfd92009ec1171c76a4ac986510f0fe7280e89b6e13e86004f745d0731eda564f679490e45c613b859ef0771be91c6678714da21f4df432bee2f229c68a2d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fdcf331803a4ce60cc7c4f6450ebfdfd4a39eca873ac8760252d321d937e6accafa9d82e4f27ed1a6dcedc984f32fca27c86929cb63d3454810d215fe5b7f616e1efd4948bb99b7f91452657e5409b332f40384a5f283742480fb885a6be6619811c2a1ebe193df2996981aeee98dd3e7afb90edb3a067972a827cde5991309;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he85d180c405fa8594950d35a989de32d166337bfe66d11514e3e40210c29b3adb6fa4eeb5a0e8b075c6d3b9291c77943d00a9d8f264f26538543d7f389b14dd9fffcf417301bdcc31967f13e10284f38a50416bddc8ef07a15d2e76ea0a41014bc5e97bb6a2df6f5f9b2f6590e7b902441aa17631059fe0c275b15323e9b0af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc537a6efdc32b292a3e4a50563f2ea00d1beada851944cba502ea1410dd08d8b2c12a01f127287a2d23c22671572ad44eea4a7ca692d4cb5f5c0b5739ebb77879df597a3cf55c98b653d5b2876ff60f8c70f6840889ebde14890c3c729469a5c377220324d5443540f31962b4742780e408917f61ea45c051ee62d0d0bf5a1d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcb0c51449a16a53fb4d64ae7ef5684c2b5dbf9c1831c44582d5fea058f5c9128f3a348480d576eb2c352af8d8a435ed6473c2bb7636e93e1b2f387a56f459cea0468e992057f01f0e7e55c97dd41933c73d55a0554164c293061df50e1140e93744362475cea6a55e40fc10c6336ec0862b4b5258e1308c871d2787cb7ac421;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd59b4421bec640f37a4719f28be6a6ec20f39ede9191c7952c7504e81c3bd94883c16114c0cfde31e169756e96da917cc1c048dca70cf7d4ca1f322f0b5628a9579eda958b7be2ac0d5eebf26d2b7acdc772da1414022d8a98c9d8f3d69cf5d3c8e3fd9a115709bf7eea6499c8b5557fc11e96eeed36cec0799ffa7ce54f2b3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7eb883ff64599c917e5915e5a08f9c1f79a3f2f6692eb9ec9b62df113877b1da2c31995e97a2eef4b785007ade1e1b2fb602d14029fd8ac297e192815401515a4b65ec83ca9bf6711eec3a55cd8e89c735852afca471353d8b0bfaf47719732dd82e0cbd66a5cbf40511a5bef57604b5136dede6dade7f415afd15843945dcab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3deecbab283a03ff6bc64df7f0425b7b31843741dc34ae0f1d50cfdc082fbceef15e4ccbff263458aa5739d1ef1d3769b4763b3f23daf547651310dab638f935da66e947d74c1bc7af7a87e60cefc4bb914c66d9dc704228b8bebda42f4bd0699a7884b54914eeb45b71f3186befc656327f3f77a6574d5aef77bfcaa437d6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1dcaadd30135a7c4efdc54a7691bf35bb552f280bf56585403f3ade914c0d66fde603cad874310d7b0b7f6fdb5a4f361a011a717a023037ac692039a68ae5b050898b0b7d645fca202f4dc005893c9f802b7cc4ef5c4c961bdb0e3caa804ad8761ccda448bac51675d633855151dbad8f9a6e6012ac02590764d1cab97ec796a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c9ab5660e71a79245b26815e8f9dcfb624cd7365d44e5c16e4e9a51b9ffa7482d1e90d27de1a99d8a6a7c9663039c2eb4c90c2223922651ca935636af80c04e78bb1daab5b9bd1c203776c8a4b053d061126d34b06160a42837616984681f180650b4aa8a80513fc49023cbf958829216454f848979ce5b7a13c4cf434e9872;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he64248e4faca971399b75c89cbf7f9dc524d9cdba65828d384826e12627f428b984754d7b1010ce88278b00302f4b07fd43343049ce92f832a73a52a9271b75489017c85335f035d011423402a3d0a2125c2fbbc9e3a72df75f244a95c562a61bb47b03afd2da7590abd71c9d571f3fffc194dbcbb259437cda1de5a346443e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44b97ad84b16feee6826ff4c21ecd5d3087406ebc1afa4c24dc3df685240fb1047d5038d2f5177df4ca105193cf723f78f32a0b2e9ccb64c91888e2cef1e8c6cd7d2a0bc54403e289d5ac7702f77ba401ffb0ece9aa41d0b91ca16fb1dc58b619ceff8a1f741d5f5091aa4e4b06749ed20660bfe4ac85cbd8da538a2dd4c4bc6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed3c6910769554ce89b1193b77c6c097945f95edfda1292a2bead046e6324e7dcc790b99264f907ff4dcf11e9196726186643cc1dd66330f6825d1212ef2d5af25792c44fd42d317732e2c442c96fca8b83be8c25ebb3736f923c5084a46b90ffa73c80ba5c21568707c9f2152a670cc692a9ddf718702cb4dc3ff6ff0cbb9c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3949b0ec1fc803fe0d0258f0891db37f6dfecc2330e738eacf8c0fad5e28c3be079a6426f6ebcb07159c9ba60a79d8b78343e06025ee21712d5598e30cff227ab72ba8c9935d7cfbe53d1b8c32232896640869c22a60666f924ab1b57984a377685231dae2ada85e35a4e2de42f623003fd5fa71282784b4ec2de96d5a4d81b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c57268dbdc91dd25741eead6ea26ba665748ff3b0871de709af6d5183df59df750319bc70f76b38a9a7583fc034c04425ab72c463efcb5ef26012c45798f56a912a330d9a40a05e3e4c7c5bb8b67824134e85785cbd47a6c4dd0cb2ec8efeae0f79eac3f1c2e147d0eda944f675d1f4434d79d4b491eaacd3366d8048126c64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8166cf1720b2f1f4c9105a6da897e5ba919f050a2748298466f4da735914ce98b6201199e329e0a3e02de16f95b544b993eb9e8df9aa9a09deb36a437cc32f4f4ad3afe83539300a451b82be09f6ca6d5aed128bc5d4d7653104ffd467995fca5ea8997887e1e2a40fac9956c42e33182ab4115a3454a42e8e74bc85a5f50188;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacdaa38f5adc24d33f8fae37f3255efe7861cc06a204d0f19f0a89b0a37078141978a2306facc48909c1e88a728bf360e5650ed9b10401d3ddd27bdbd6ec3a0426c15c14db2faf393762001e8f652fd4abd0f73dad8235b9703723bf801fb7eb5190f1dddb996488387ca71cbea358ab67d3134059b074cef45bce7a687f555a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdefbafa6e48b79ba51d2401ce633644eabd4e6fced8a41b62e96fdc914ec1e022b79efcc079019132fee366227d4cde948e08468465f9ee91592b658dc1783e966c3574656a624394cd08dc3d71ccc161a3d0dfb49e25903c95bf31c72504111e54ad121c31a1eb792c4d2867c6e36be475e827dec324c0327b915c5ba6dbbdf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19a8245156b943bf86590cb1e8d68d622d83a50e0074ff0b5d473f843065f4ed14aa0ad554ee68253a03fd2fc98396af6cbffafd6747d6c3e58bce0005724e360f14b8734f5378e4cb892c8d45483d7abea0a77f6789f01f2d24e3da9989ee0c18f064b4735ca4d0ad13e12ab8ef77965c7a5b9aebdc85a4f085b62b470ea9fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb60231de7d7d2779896fd8e8854dc40c1fc057935eea09f76ef7997eff50b18ba693da56dfd58f350ac116d0ba51f7242c08ae65a4e57a42313d43c7c2ca8702a29ca2c89f51163c61aa3ab81158a3af481d931c4480792cb0131e2992b595bb664eda7ff8ca0018b68120a7ae94b428666cafec0d0e2529700e44acd5f8d321;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he671e1ba6d7893890dbd5de6c0dde25ab7c4285c70c39c6e677e75208c7410d64f5e565ee3749c2b455de36c8f4cbc3d0f509b82c8996c6f56586c50f40a89d0399a23ecee7ae009507c4726749cb3af08e6ce8701eece5dee77a453139cbf403613587aa7c6ebb716f8ce7e37bb0bc2b2b5ff0b5f0f7afe25092c7e89aefa11;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h634e5d00a84379555b97f3ad341963edfb156488b04a890539e4f5800f60c0425ab07495757bb367755917d983f968ad245e287c0f26f2ef3cd53eee38c799daa2f0327596d6557915c19df1f1cb4e5eeeabc4331f67d8d285ad32062d1332d44df9cbcd5e0ab12cc496763cc5eca5ccb6f9fa16d095771792453c4ad2574e6e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d6a9d362442de081216f8581be5957881b0510dc92b467c20e25d5348dcafa2bb554aba34a4e1c5f3d771eccd0805532732d5b32b284682eb28820734514a471c1e2f8cc916fc3cb5e4cfc877c6d78b5999afd2ac35855d95d2562ea67a26027d873fb6f9b7adad01cc7611114551208d388f88e6894ac8451c09c53e9e6156;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc2a66419aebf04bbb5903d1ad753b81f8a01b40f12b8f68c3afa5ea6e5d96e9c10f374c7683a55d2d9e69519bc16ae1be5db9de489e10b11f6d905ce6f87bd2688a33491bd805825b9337e9ee41c03ca7f3a25711bd27dfddf4eee1ef46f3e4806da73bb2cb7497492158b824a9dee21a1e44979fc8c68a1b2a40b0b58db03a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ec96950e02031b02214e43f8b5e78f7b4522278aa631a1ac390493056f97afa6161c40fa7b4fd141b1e1001e2f0755ddb8dc57a233ee513ce6c0a0a4674fec9bd18289a6587ac76a15479b0af8938d07dde86505ea6e2d451a0cb8940b46e657b1cee32acbe817d0910484392f4dc66fd7c666cc2186594afd114ef4eb593dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1eff959893e88a105ba4010c9786667275249a480464103ccfa843e0f6cc1c5c9367285b2fc2a5dfb1e63410c31dc0f48c8aa3a3f89a91b4d4c3478f5efe3e3301a4eb66a81d0deb8acfc0f0dbab7ecf71c81263c9970ca49c9ff43b4a2dcc06e527c91cbf3c152443fab7d965194e6f0deeae6a895b84c25c41dac1a869f821;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd28d3d431e4653e1d9c7467acb7792a07e2820c5e3c7ca9bed82d102e632cec723cd627f5a4005063cddd6f0aed2c477c56689b87e971ee364f56f184898a43126179cacf143f51f02e11ccc0475cf9ff93384d8205c7b63533368a64122b0d6e2ed5de9dac237d4bd372a52165e5f2405a16dbf019b6884df3fe090b1d2648;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3b60d3f9ba36690f0521a2b4b376d74784e4dd748d56386516583d246556a5683243c56d92ec19d2f7adea76984e0001bf3604399aeb30d384bfc8ce1598a5109711b64466866a277f1922477707b4b222cd916ba1f31c01a328c43960db4a35646756e6b050c1903b241d00b9062eac109c14fca7024632ea91578e5391afd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9bb7c85029a899dc99b77501a0b707a1671e549a7a371b37330ce7314e1265fda9474d33b618abad73f05e7e0a609b80dc748677cfebbd0ca69c8ba70b5ab2d0a34e8e3984877617b122e5afb6f1d4b7b07c6e89098b19f0adbc61cd1471c42d1bb190e8ba40d45a5b886dcf8cb1dc2165e833de183c7f214a1870fea21535e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44a9d36af1c10c5444dc82a5048cff827a9008f31a596a7ae2c36c8b69513f1a0966e11a832c369b039a9b5cf861f359b37864f9b0bb97d297e5b27d9753b8948628eac3d79b0d3c45b6592c1e57596120312a912b833df07f2e2cd9833e4516cc0058b3b8e7458111a85378b5c950f678300a6d1ba904d10e078fd7df5d1137;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c064eda410264dc14241d0cea96b65aeadd10ea4db67b056188082673ebfd04ae0aa3085d27d1d17d28802e17cd75e38d4d4b25597a5971d4e9d89a1006360c220a5243438a0fad6c0307b0efcf6730977601bd97a41c38df60b1136c68353b51335282c89063cc24d9075523f158006dfb6b914a29eeed5f735be555e4fae3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h598fda28cf1d5f6218a174bf7be8a2d6bdd02135a382cd0d5a8320d0b809c17b3a09be0641fdc0269be5ad58fae2ecd2c5414fded1284714bb4f8064fcc68f3f347749916b184697bec8b2a88599cb51e4e8400114a5d3915b3ea7c918a88ab948938aed6d51dbb97e781389281f823ad81d948ed33a94b1d857b3fc072e0fc0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6a7dd8433bc4fcfbd6b0e191120c367219863c37bd56839f181f38f87f14eeef9268e1dbcedca92c9f85c6671af80274397343f5fab83d48675270efffa2961916017f65c4a29850c2edfa9ceb187bf20b1124ed8efc92f1784ea5ddd347bd5df11b8417cf1877efd721fbc4e630c233d7350583e408ae033e15a7823cbef1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5957fca28722679c18bed9da3d00e3dab0808928f23bf2ae80df6a80c2a1d95ecbe0ee2cfe9d361ddf041f009273591c99dcdd75eea256ae46de6fee11b075ec5d803f161ce97b5c5bea9a8c2e5d99159fbb6968dd2a17ba6e84c6f01391d575841bf3675f52746ce39a12a336fa18d08c9a7dcbbafbafaa7dd52b451ce24159;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb13a57d76f9c17e6c106bb8b1b0ed1b11d4002e8b6b3cb42e503a9afd42421764cd077ee0ec4d39a5077f4c7452c5ab57b58359597e090581727960303c859db6abf29c9e1427246f54436fc37c0feb7916e8599041af5893dda7568b41fad1fe18d3f8818a343b4505b9122b97bc6c2175bf4e3a570c3dc6308765800f0fbd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7aba531594003675be1675aca5cf5454d2ac9c288f0b3f27bdaf5120c4ffc0038970a8a25f7340fd3ec715f413a17a10222b5712d0595162efcf01d9c556e39cf9c9f58c5ce34e164361f4ad2490715d5ceed128401924111a2138dec38eda36ac15c2865e0ef6f4791e47c90b91bfa0d35b58c870a6bb27c0dd090199348ea3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf317c88791f7f13909ebbd7f54f766ab23bb722ec59754c2866e563a7b04842a38a7a88f87b6301e72ce9a8cd1bb368c842a57f1cf2c2b7057a42276a47f295b44e50b74dac42db384d7280ba61aae3a63d88b1edf1e7a474255a422aa7e47131ebccee03a8371da92a67d29d8d44a358da19005afa9fe88b0731ea788bf120d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8d68a951d0e72c7e342f30f0bda2d5091cb5b8291f9ce45bccc098e55c6b40e8281edcc1caff81406403896ae04793fa9bcdcb2bbc42a959e952c21d970e7a62bd24e1bdb6ac55bf34b8bd8c5d699b539095436bf941f5c612513e7e3aa5a9ed5b40cfd67f3406decf7826a84ff976a3286ee4aba786857ff6972f0485e5985;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10925748e5525b59c95ea68427b242c17400561381c460620678f7d0935a761ec83275f76ea030646acdfc9d923f7dd4e2e83c6b094d21ed9e2317f839c6c3cdaeec95d723efb3fb96f81ed9307091ab04081572bf725597914ca4558533310de6de86f1899201a8a6ad4da5654a2f6e71506eafa453a408d1de83c763eb9791;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fac007e6fab71e017244c5cac5380a23e3d4154f984ae8c88881bc6dffad8681c700202b6ea23fdedd6adfd4ae32255cc922d3bce5fdc586a4e9e059900af1aa4b5e8efdfde974c9654b8395ffaa981879ad5a2a71c634b87b41b51a16eb78f314ed60a08cb362f7f52f2fd3e2d0802dc0255b417834f9c3d6493eb930d7b9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e794be761468e852100def35079538b8bc26c2c872b069e6928c764c70f735a63fc8e13a90b4eed86184a9e9a894caba587eb29b7307b83e8d6069391e89942e8d1c3d63b9f15c84b7fcfdc7ff0db56019091412ad4d6abb3fa7a93b5db7d019271bba24deaa7295c186391c8dd255403dc0f04fcc9960955808f8a2e26cc16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33a89b56ee0e096518321c7b87f52c86bbad520212164f78a6668a37966f40c2e48f9e743fee44a3bbe43634cfecd90a9cc63664a317889509ac870d335a20647f8f97cf6641e2b10b7c78aee398a14a218df49de18cf58b6eb441bf9a01a74ba190a09ab070ce1b9116a208aa1fceeec6675718375cc4c1561b4ebcbe2b85f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4810f12c4f7ccc5968fdbf3c025c4134bf05e6d8dc7fd559b47ec2b86189bbb4b6299bdde0bcb671005149196ce2171cea2700fb64903f591f0564ddacf61c8da436e2183c2cc26af3f366951eaaece9b46f373dd01d4793b27a46230a5498c8eb309b59c7e99dc1cced1a654ea47fe63bc4078675d943ec2b4b80adb846ed01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c0e74a055edd3507b21d718ff89d555ca3469cdb3424df310968da7b6794e1aa88b5214e6fa3fe45e76a237f80f4bbfc9925c55d55b9459d343fd57661d48f58ac20fbcdd2e83a94c60f610f54094437480abb007f4a956cc077b39c24bdc7767a493a3d316ebedd1c552149d73a18122a26c07f905e1791fae0a2bb566f1d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbba1d4915b5f76445327c18a28f639f99e1f06e0dc41e2e2e6591b33d9bff7189c4cc42baed5c6dc8863cae60ef5d841b2fecf1d4ae81a3b2050d944389628862be11d8391774006d87279a5ebebdba242ade58ec53950e22649f8075a482a58777d0d70297c8f6557f2d6fb6e147e3cb6716877ff78ac53548087ead6c34b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c73b020c9a17999b1ef86137255f0a7439c6da0f067f4fd92f08881b84d704dc129580927dd9b20fbd79200d8cb4e484c2826236098d656f771d510049829d1c4d9681b8a26b5b5c31a4a7f3d71053234d1b8749d03a58622d4c72acd96e45ea8599cde7d184b34dc83cbfb4836a9e1e30a66ce622e548b1d2663d7cfa49b65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h777b1bed5aacc610210ae1a2e5c23b311b45fdfc7bc429966b89c90512c2413f8649ee86619a7d49223d5a44775a3f9815843e3b6232bff3f9773c6e9577cc2816340c0947967d5984f3880f934c358694e591ed313df277aaea38c37bb6da3b2e03dd6cfa1a881ac13239c3ee1cde9312b6fadb6f9f77860174398d90a969a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f81f707ce7279fd0217806dee665bae429f7e5a3d1875203a434ca90d3e4cf3e1ad88b5ee4cef799628fd183bd3f0417c55955db762c79ca5406d2b1cbc6ea97dfb95c69525f4c3756ee95725ca00c139557d04e38fce78102a310669c43302e0ed88e22056ede8dd6e80db50cce35e772cb095a0013ef73bfb20339f771769;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83980020c7ef0231298439d8362035e696f731eb029b0ce7c89161be1101e0355968b4911437431101f8f2ee1d3898e90ef6da6982a3bc30bd605c662f42b52849a5d83b029c8876ad92389d43ba30d6918918190d032e7ddfe172cbce26342b244dc19099bb7bd1f391adf7556076179b64174d17c8bd20410ffc34db4f835c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb2254020da4771c5fbd52106eb92bac4bf332f044b3c754b62990d478b14602bb07987444a565c98f51d1e30f6fad9a3c0f5941a04768dd832700a948bf8719060fbe8811fcbd6eab46fc5801c9b0bd9b05bf941af148fd951b259e56513f78f1512483b76a8ea56f4b67cc0ba2854fe3f7e70aae450b57257492d6e090677a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38e044a616550acf4caeb20f0a21be5ec1c59ac20abc9f9d47f886a43903c1068956bf96b39d822e68f140c1988d776e5e870a29835f648de0a8c5df5691c14d75bd6e1a2328fb863716a6704d403214c6a8b7a8c74c56136e887eb89c69390705878cd74f9eb5af64234188aee1979ec9ead5c28a2ffeb70516c18fb39c627f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e09ca27677c42389749bfba3f3df742ea599ac7b5527773d7e33ef00f342f2c4fd13c403ebe71004691ec73593b4096ec48f4f1ad2f9b47d1a0c324090a249abf9a66cf19b11077acddeb740b4fb5c2f9aef2e5b8706216f7de78c11ebd0d07b75548bc44633f2f7172bd9a5f5a538ca7619722abb17abe1069001d01733466;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1333000ae5bd80f2bf8377823efbe76e17c5b721fe1ae7aeea1c37b29e4c1eb5e4e1ccf2b64b1ad93e9720178d7ab2ad5e64b613d01599994a27db14800af8b5ff19816d26f2e92d4a9511518560532a7fa7d16ea4d319ff3adc284b23bf44ca6e72b98aa88091a14a82ba0ae2bf72bbeb347bd057a12b2e0795063fb2b7d12b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h571b54924a41eb0565ede81aeb66f6ac399856206b0d093d6bf34b256dae44e5650b15003260a7343a7cbd452057da1e93490b5e8e9f45844250303817ff1049ceb3a593e876aed7ce916cb004e173715ccacdbd8eaa5ef8e7829dfd25b35ce28003bdf44cdf212d9b0feea61242a8d98db060d8c2e63d73e3a4a0130a6ad271;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdac31bd65ac30da447bd5e5bb4b68f8e2091a090bcb0232ecce8cba892e7f343d47856d8a5a39c2797ff6675a9301cca9c7e09fd11ed3c1bd8a1aa542f7ab21893a9ff99252c46bac09f91ab37cca3a92ca48ee3fadbc3c9484faf960e2f47c715a1b5e7ecc77ab1f681179380e485a77538f16d723f0c0396a782b95838ef3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h776889fe29602636b176e39042aadb932539e57f4e1693685c473f3831fc49aa46fd3122220b674f7107295a313a518d2c271f1ffd18c60f582dfb53f8c967f86102835364ed5200e0373bcf34c55c319f266e2aff8d3708233988b073f8ae8eb152644985c464f8705c613fb83f8980f8c04ed3877e207ce64b597bed4b78ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6461740b92afbdae4b23b8fac3667c40dc6ed4d5afc6738dc4a967cd06f13d7ff3612334231e0390062fa2b0d65cb02989053421b27eb30cb80d2a3e97990406e3c51324fb522a25e9f906a989251da8918a80ff118f8964f80dcd3b4c728d8094eb0041159058f4f436a13ef2914418c6dae6033b08d564ecefc424f13ad728;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha50651e98b0a9f486e7afe433344b32f5082a4c7986517b580e9fc665590c4cae5f71e4c5c4df517375ed152cc9626753d1f3ba35b06ef98f22ec7986629399bb049d6ba109d062699bc183eb7c26d058c47893b3e33c64a8600d0dbf5ea072a616c0f3c71b99eb10216ff1edf90df5a0cee87aa16fecd529c20d4ad1c0da9bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha58a716f5cb99b6a94e0e4644c3fd5e814e1bdade2c3729840dda3971729a2b8b0c216677069933666ae85285d1448ecd900378dd3452debac60381dd884bf3055f4edd98592dd1317d9f738f5c9eea696891fc4dff70baab06add1ee11b934cf4b6da310509cfa5f615b8b0eec6da2a26f7879db4ff338b418d00103c82a00f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6647336716443715c2fad2b877bed40d2f76ac9125d726739930f6ed6a659fdb782b4ca76f5674b0a8ce0e433a28bc5f1983a6f10791d7484a2eb34e3d832f888081625f44a659b36b83cc5af6947e224ddb033546586929006cbc666404e62ece92c0d3b5b4e10cc8d13026c9b3a06a04f7748713b6330f9588df840b7fe304;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd40cf0c68c83df4d7b1fd8f32b18ace6d2b041a0390ef271a49db0d53c6dc01837e8d3e86d0f84859f4567506285bea9798375858ce7ea1a7ebd249f17bf7737cceb00bb5d156b5d9e258f213079068d370bc057558bd39910f7ca9aee6fd71cd9de3e263f15fb9c6b24dcf8c77fe47ac59bbaa781d89a9b58445a2f6446d47a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb8dc0ae90b6411c7130ec97822a70c53ac085ebeb7d0cab15568c871dedb1a50ce57d9055085a42a3c473d988db249da2ee0aa0dd0eabf7fc16b2137786e99a8399e62468f3910644d98431a1e5f341b4a1804302e8c9d4bcd663eec3081ee30a68150687acdabd46c882430ea3c114add85abdd0b5b626310491cfbb2b90c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9d66c75cfde873e35942fb4eca95876071431aad0bc71c82ec14d74ec9b1335a9b8b788ca62ef9c124fb484ef51ba90b430b0f6e0bb4e77602775e5f04e53de6083504aecffbc8454a4174f3dbd9aec56d815a163fe1e02b6edbad035098eb50db5a27f1f977e7ed61c5927e1c0caf96240a33b7d21a3d5fa0025c3a47b4f96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86a29b5ed4ab187daf16b691be006ec5b2c6eca467e350b92a5f3498d6f1954f60cfb5f2f0f4b432b28b6544e271fa436f50f8d52c8e86d60a5ae4d89fdabc8a8a59195f7815259e821523626d6fd89c290dcd3fe907ae78134683e0135296ba66b855a04a25289f2cae3d1ca65043f42241b1ce687d81c2b666e1d7671b0d6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h333709ca02048ceb11658c97589b38fa76ff4feb7689972e89abf25ca8cbbe587f946e3970b7a81c608aa5c8d98dca6ea6df4b8991eadc351d7bd84be09ee7cb8391cb25b89e509223de7c52b5d123b8dc327f7b1d3ef4fdde6c1e95447e6cefcb19ef44d524a6d7fe1e71c8d87abcc1065ad2f7fe0e92b7c456b3f182478bc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h638b9ad638c7b12407200df4c1f9c9f58a9d53a7ed39e0cb3df7b19e0c411d262ac41f47e4983f9515a0f43d1bddae32a93a23cd6b3a89c9572ee5212e5c2f697aa13400ef9b597ecbe9f169a7fda3bbeadb38369716592546f038491f8d0f09d6918de18631cb68eb787da8558671469b451829c7978c422f6abdc17170f7e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cde70aca8782ecfb83ed4749fcd2a023a7e315face16413ee2f09e99bc6ad64095ab244e690144bd18584f96d4255bc57cd11ad1242ef4005542047900ee8ab7133a2ecfc7fa6be3da398b710c834989b2a52ecea5d22ab0855cdeef6fe164f9000148b05c3224a72f908ebff560c5da61b15bb705220776c887048a656c9b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dbca0a190352f87d50a84697252957fa959b18e4e28b7521bebe61428a52d7020932e240470230cccee3670fc7779a6c6a86bf1b60ee42917f1c0fae4aa80c578f2d0d3a025a42b27c24b1ff30db1d5d1860f0a81c4ae62ba332afa80afcafdb71c238e38d515ccf5b34f3af22a06edc027423d5df9d6c8bf4aa4598814a258;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c4dce4e5aae5bc794f980133b2b7ea319104432fc009a8f9bea1c982d13ffb5c4fd3e59b47471b61a3ede4566a881c68cd79d323ad21d2603df24b6e08ccc8a22f6a5b46277453b0389a5ed10b44ffd5ad3aab2bdbb00f93858fefdab24a31a2c013256103b77fff997c04f3ce069d54d2dcbbf017a3892b42d88a4c3ba54a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11121ed75bc2916dd753c004eda7feb230ced2a724c1b88453d2fc0a4ab8274d6c741cf725a081019fd1e25cdb0500835bb6d47d93f8d3b291c0a1d06336c33ae658e332fde3adb00681a339622a1f74430dab5263ed396887de0725edb06a067d05d241537f20a9b81f90c7131e9718c4c0185d8f86f895e7c4184adb1cf1d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b90d695a23aadc21ce8e52657069515084cb58b3cd8ce2cb7f09ac82e5e73860df1436289bc9b167236c8605b83e5fcf49d49d5d684f33c4a8ea7c337a9710f789b03bab0cb2d6d39e37a41bc7c77deaba801f62cd60acf2645b5f12d45b3b77c644bd8c2927cb54ec2c09d17fa0721a59906d28be0aa9ab919ac90060df8e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e4387f2e6edebb3239feeb9bc6ebd9443db2ceb20833eff7f409d8175f2667b69ddb5d4449a5757e11b571247421bab3607f3b0e504079f77b39c14bcba27bcbc374f32e14e4c550ce1ea506e57ea2c2cf26e07ec06fc3c2b193761414ed760c02bea66535d3421bafb9546b509ed2aa66769525b883cae414b9a4372699512;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdae218b6152eef9d5c5261ea32ee7480b8c38b9691248a4e55427e9ea6b5dd6fc3d637c95cecb31d29895b8e3cb0e22d9610ac42e3ead4dfee983e1ff252851e1357ab12288dd742bb9cbd4813c6e0e6c3f85053d984678339ea7346a74d076930600ea0751301c68047ff2285f32d513399c77ec3f10ecf98823b98a8d261e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc59a0a476c0e7429c8573218fc1ec3a40a3f65409c77b4617b41df66ca8718eee4e61ff1ef13cfcbdaf56e60a879fa790564869e826ccab7146b710d1963fad7af016df8ac770a0a73f7d8ccb4d1dd38ef60722c936002811704c729b48d87c5985d213a7e2855cb205e1278c87984e88735b3a62e206fad3601227445cee99c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dda06274f0303d5df7213c3883232ba30ace6db1c5022ffc0ed087c5acaaf1a232e4f3f47c98482e77b2dd223ccc1dfa86f0d8247e480514c2df50c0fff30eac4d9f8cfb77d841ccc8292a86069b9a8d902ffd65b5613bcb3051ae3353d6429205e260f86e80013cc746e5ae4aa0f5af18b2e0f139faa8ecaa0def0eba9f540;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cbf01c9c615f1b7ecc918db77cf0864bfc91353aae2eb230eda4b99a199449d51a586178a0a561bd7562c0212120574595df824bc561910bdc939f817420fb4b42fb43c24a0b748ce29d6a42abe5eedbcf1852137855b3d70a5bc892382dc2d9039edcac410119fbe1ba273460d79ef7068212890889c644318d3c1cad65f09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cabc4a4e107aac86468e570f0de2e03727458de1f67bee26dea6695af3d204f2f3c2ebf0358a9d387e95938cd0f8aeca784e05933dbe1805aeb48321f666fd7283bb93fd103bef3a15086cb647fc886129d994b9df83a8eb835c711a88b70bce9ca7152a0f2e8f8c81849b489b2424c42e0a82dd691912b37d7d05f6a9f1738;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ae53181779bb268fc8c5907422d7a836911df4daf57f9b79dacddfe1ef8d01e80ccdf231f8ec81b8937ce8c45b0054484c59f968ed0046b86935dd96a7db5f095dfd9acb51a4a2b5e8b07b6b60aac80015b35443f6f1398ced79d3d26718fced4c7448226c591790c5799974ecc27b9b4ce4b4fcd815d65144228b2e34f22ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6050bad7067d5c70199a15c3cae7afa61609d4d95dd09fc86590604425c0b1f2893a2a300e4d3ca1e2cc9ca101620363d834b6b1fb4e4c4964197e17913b94ec4446c9fb5bf958535a66476996da2375604ba03487ca05cc096a6f6898137e4d165c388e1384d89cea248fb85831162fe3178062d06655a0a1d1dd1c7aff4ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe31c963b938d6e6011494edfcc7c3e07708e97f43504b1ea4a0867e6897879ff09e73cdd704725f43f1776cc9440cc8fc9de600dbeab37422b4de3b8d8dcfb917fd1676d793c608e86c4ae8413aecfa729bc3a1948d816d5905e85ae46801e37a74fb602a158acb03620a537d3d5c721535c206e7159420e6a8c2d5ce4cb856;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65d2e34c23c04dc05b241173ed477703fa49bf59c5ed726c555f6f8ea0b058663dd75c6c77653effa49d0b2c32d5a4e1667b32319137d5b94e73a676ce9a8e3f949a85310b621f455907c1f9fe5f8ccaaf37764d9cf7d229c4e69a3a3e8db4003b8b1ef7561742e1170a86537c21e27c77d8f9a71ba98aaf924af0e3c6467de4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4c368e1c01a75f4a21d8576461e36364a5645a016bc98d61ebd855a46a4955e60f8343df6eff7d5d5b99b4d1063285da8ede0c67223d3cb16b11f676740b9c169269c8f616d700a60a033fcdd67c9ff66484ecc3dbaa982d0558728ed4527d976a9b29c424f649aca340cd1f6e40958193cf56d2ee9dc1eaead3952d0b3bac5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc06c4b0466d3f85325acdac7b304b1b832ddd18e34c81a9f82290c06da2b74aad8bb706a3a1603d7feb72181853bb42a62c4f366ba863c197c681f489f84b813554da96ade10a9c826b93cbf66658f7c5ee24f5d7afa71c69e1008ccbfb250e4cca82a5de80c6ab8279f480857822c37e4a2ed8f8276385e5903d2b5ee64da9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb39e24e7f2f34afc9b49dd01723cfb142a012af180e1ef411fe26f433ba3fbee4c8d7e49e84a08f15b9fb9455b23549bb0d5a0146a7dff78864792daf77f50cdf7239f576970fd5c917b2179c53a2bb8f974f157f2bdecc58ad8a5e2b1ddb39c256e5d03f55daa2fd5552c6ff27ceb95161a37dab53653775a291a76613d00b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82ba59155ab5fb5472bda516947746387d77c10d884172bcc4a464835130674dd79755484d56336e4ed1dc4b00bfb961ba914fa0871d71a775881daaa7fea9dd47932df454d23cabaa44878bfafbc3ea71ae42fd8107f2cb709b09b61abfccc3a41b643ad60ee01091371868f6a20764ebe6e572b216548793c203ffc9f80806;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93c75ba5b18e40389c05de184561297b5a6ad63f306aa7172b3982712ddfa6b6bfe414e9e0d344f06e8b9bfb0f095b8b02caeb4184a3a4010fbfc41da36535914f7c67f29529dbc71830bc5689e8acc780e674a31d5183b3b48a320bc96b90adaf61a7786e9d757318aa64522efa4c8b0678687620bc3912912edd80534e358a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h413c110d4ea3955d7a05570fe8c3b26339ef1d0e37cac028f62d5159adc0983ca3e74beff5300b1b5ceb12fddab3fc274864e2c02d6860e0c2607caf08eb41148f1715d60bf6715841744497b75b83401d8217e25020515e27462b540400e2303a801e7214c1bb53437e50b82389549c56e0aedd7dea79e50b4bb1884051787e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a63fa3fa43924ef349a101fe3ade7cbcae1b5bee86241e12fc91b9bf11dbf5e581a15a26467c51be1efa5204553b2b93ae0984f065b8190b78a86ccf7811dc234e8e4189fffc601086007f6472c5e0b514895b51178f8efb6d219a6136392eb270b795805083e29191a34011c2ef0a66d23f1caa2a176a6b643beb56037bc14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e402710ae69e81b54821d7918ec2216505b1c593c20113c04aa0cdacede777b32c938de6ba3fff46c2c6a3bdad2a1d0a8194d86846061aaba105cbaf58f7812f4c2c25ccf6acac0eb69cd804fba4bb05de7cc01250c87c8523a853c103a8c443a091dc6d27b4a83f70cdd7ae1fc6ea62f67613d9749ffe79bcf0f4bc72fb63f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1368edd5634384f6fa201cb224a899f725d91bf9087589527c27ba05be3e22d5e0a08ed6cc5fbdb9ae2f7b798aa6cb73a032386b5ae7eaede242bdfd1a360d5ba10f0082e8e40d2211543129960bb1fb95195051fc8f4533acb87e571786997ad596b6ff761af72da794ec58a0d3964fb16fc4e9b1fbfb733187cdcffa0904f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e41dee359b37d347001ca1ade6fc9aa5bd767d3312a80b34414bd21b530ae79657625fba07ebbf4bfe26f6ab097f9b4b3856b996a6824951ef6e2feac1aabdcad358a960bd644e8c2c8bf8201b758d8d4c2a8f6c502fb109d3ef6f66cc45313bd4db70792da4f86af6773ca0413d7b8bbd305525592e306b17f2492bfc124eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78f671c2c015e2b6d987ab5ea24ac2d6b8317d1bb40714a1c9df481a542de26cd702a5cd69045a5defe73fb90b55ba8ddab9c6e75f4b3419accca09512b52c8b6528847d287b048bd9acbbcccec3c89cf127e5458564eb49b5ba4dbf77899ec97e386f58fa6a6c51c2533f2e8f1f75a1ef48ffa2c552e430dcb6a6bfc16ce2c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba22e524959b1bf2dad4e988d395b1081fe59ec7cbe4a7bc2398b31ce9ed37460fb65287f043806447e1f3198561a7650e8a7c1ef164eba7692b9135a5ef1df0de7764ed7afcea6144bbd20f3ca571d101945626b30735af3cb570463c176ecd43f72ba5638406f48a7362bc47e1dea703599b5dc2ad712f8f7d6b818e5a2040;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4f99fdccdc107031e267e375924504226866da81864e645b468dabf5614b7a4a30e6dd98faf3f7ba3003a8a83b384a6566c1147c505388f6a601935629262cce707098dab8f26a27ead5b262faa3345ec0834d6f35880a2d6832b5d92a7b7ab27db49d3676c08777d2dd8df4c5225421a9df4464260deae1ca23ba2846a0303;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecdc249dc1474adb8b3b28e9259009d3709a5c92f9f30898a442deef76a41d3e986abfa67aa6e1e2a606cec49c4fca612619ead3e30000800db73736426f806cd423e3b95ff293b9f6a9dbffce7a0743ecc67fb9151bd443c19894fd04cb669242b9748261528ac6429fbc7bec607cb3b9f328550ba72cb26c21e1c1e6866f8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h465c32d0d8a2fd2aa0c021e3eadb22bcc61eafde50be960aa9bcf98f019f55b6153d8de333e2d3e2874c5cc38f23550cc6b450fbf3a02a82404a2a3500bb14a07454747595b7bdc6d01dcaed19719a7982d8877e546a251035ed414764758ca5ae3e93f705fb9fa79833c84a7184d90395f1273994be37d4ad0cf183883708c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5238d913a0f78a9084fcdba0489ec44e2675a7e275762ff3a607026e95bb9eab0722a9a41ea62425f54d86e0cbfbf60c38f3f635dc2b923929695c7e8bb05a5e83253eba88d3892d4d67f71677dc256ea17ed7b1df43dbb76edf57acaf8c502ad91737dbec755b5097d2168dbfe51bc04fe0334fe04fca9efc125a3b20d72dde;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h279d371084f76eae29c9d3add71f0d81e30a7749ba938a149352ebb47490383315f0b132a447d8d1df3a42d82dfad6069cd39fcafafc3a56980dc72c0f53de6aeca06118354db9075757ff1c99548bfce0eb840b5d2f36d5487beeae629f0bf8ca688b9a0356a6fbe10d59933eff5587391a83ca04d7a11faee19e97db6c1786;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81ca0480ce2f7d513612031ebc7a72afadc92f7c60a0e2a12f83ebe4b6b33a5d86f312d129e77f68c23213375df0411a8bf11569d0ead714c9276655a2807ae3ada62d2b315ab7aa2d6438aa9e3432e3e5d2b39f4fc410b1aedc50ae1d264dab83970205def252b695be7392c43825c8880cfc8a5900a7e99f9b3074e6396a45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdb46341a07835df0f3fa503bb39a8dafcde81cdc27ad85345ff165862d0696b8af0a2abe91a3b302cad407dddd8ed1ca13899f460ec4fe5bc68d79397a5970c60c051cd9e3c7083074ca30fa312fdebc044dd2f7668b35c0ab02a41fe63fd71060b8373e732e41ea9bf88165ad4eb99fe08880a47135d33a1d911847e367033;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e7eb6a3ab06dad877fe0c10d6fa29227a78a6d0a57aa2e8b911c7843829d2f625c8eb0ce14939ecdf70836629d5728cbbfc49ce4c6d4b483e308747568d29b93d6b8cca230169fe700be507ec3324fe3d7b13c26db079b8cb3194f2ef327771dcf4fb6b0af1c434ba51694d93fc272a0f35226fd2c185cd9f506419c4975df3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71d7d5db024f2b3438c057fcd306e7a857470b98027b6416d880e705590c51c18d08c11c9fa8fa570b9bd9a9189663407f54b0b1ecee043b858916cb62c47f15d2510fccbdb7c4b83f274b9bef6f6abe3fba2a08fbd8eb85b25f91e8b2f6e01da532350dceb7f3cc0dc58b09fbc70b7599eced3ce8e2a763e30617584fe0611;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb863950a7ece6c69f4c1d35ec280fcce99d342ce3bb74e2d67d2d05d27fac6bec8807abbcbb70709503ead6322389030e3015aafc00de5a657b88b77909f724f7b930082b210d8ce0053b0f8873373e1ec572738abee2c6a1e2b513c64f2b13329013e804e4d40d5bbb0609f6a4ba2ba91423d82609d4105300e0ce29dc8f66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h379ca7ebc0c1f0c2ccc5104038b17cbe2eb8ee9b8eb27a6cb9f50f82aa0063f6de852db3b73a9b0d0f213987e8a443672a53b098ad3e5f285843c80c28d4c816f8fb1052be040d908bcad5cc1a540f5adbca17dd4a24d7673ee6cb89291c83418591628e340e48a2c380265a82a3cb7836103f7aa858251ae212956ad0a1a7c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h161d032a6a190cd888cfbb122135368b4bcd4442087dc6cdf62e52dae9c1a397799601804e1c34529d1280274c862791185ba65693558fd401f81ee1abef8c1301645ff6ebf278481e6f2d9ebb203b05c5816fd0cedb5da4b02a5036e05efc319bdff34198da7a5ee039f33b9106658d382deeaa9371a83bdb04d7267a34cf4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14cc17a351c56fd1230447829fd40371db57b56b2454f90750ef1679f9a00c303f176db8ad3abbc139919df19fbe091299cb98e41fa31cd0e2d1b764ab48e4cf859b4af2ae843d777879a4ca9d91a6b323abacf386c866cf987e9b8a509e80aedb83cc13a0984807f50929542a905612d1ad395a9fa20fa59b8ee796e4d9cc22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h498b1760e2d573d66ccdf15b7a95f7492b85351f736230de3e7952f80679819894e6c63aec081f41d896e66b69ea12739cf7f81d24276264733e88042474791bf0eb0230139c359c29a829a4e0421c5c95abfc0e472a5072b9394b75e311cb68702f5dcc4eda7024d6c2e66431b91e25897d49eafaeb3c2d34d6bb3b16df63d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ac8695b185a2dd522ea555c43b3fd3e350a9dd63975ecf69d67a47b7b5e1da98df41cb52aa8607c56b062a22641b329b5e1519a5f8d8403af3d5e0531bdc0634f351f20385582913b97ffafbf4c3ce95fa22ee08d3245072b9f9e3d9510aeffd96f26ec5aa15cb6b97a7d52fbddf8cb517d80aede180a0eba6203699e31977c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71d471d16ccd94ac6b5f7f63663a11fb4c86c6f4516dd63d47447fc7edc82c9946d263edf89fef3347f3c87a126257e0fbe0640d3bd9c7eaf872988f6e36b3b8ee05bb79b2c80a7f4efb0699bee3107a4ac289723f41c3b46c0ea50fa9adfd5ef33e9bac4d4883c955c4aed52ea80651542227645eaab77c4a41e3a1eff5a855;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cebf501b4b129eeb2b451f4a2249dcf4de142c5b237f77135f9573ee877e6b983467e5da8606919a1e351cc1a2e9091ce40ef5bc7387b19fa20344c73c7d1fe399ef8fc60b086a443840c5e78c028125e5cbc45f82c8d9a835cf475e373fa2be2c83f6c68713438a0d34e889e1004ee1c8a19311bf9fd9c4dc5113ace325c7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88ff494f7b07581794a15d96234531408fdedf73df01673ee657742d986ef814d5e7ec750902992c4c24bbc8b23ad22633c32e8ee1b18c9a2daa277e068a43a172ad0023424fca2234d47e6e9927025577d8a2c71d0ff8daa25de88ee43ef5f01c918ea214fb803df48b7fbd15aef5d4e4d4a53aff1a05b286cc6e8ed8e28935;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b592b3e045c550f6bced293750b8ebaca52ea3e65528d63f232079e23c696f2100548f5da90b4a754b53f92fb1ca07214a39dfc445e186471f8609feec8e58d9c4ca15a9945b0e32c7c6110aefdaa3701331e9a52e25a456b256b7daa5194fe28f45cdc4254e1acdfa6806e52c4749436f435083a94c1f43b4831ddbbf98a0d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1dbefe84f12de4323048d63a6a6490a79d51e32f99729bef0b5af7ea9f9e848b834c199f030f71ed4f5e5de0ea24a6177cc55498fc94515cdfbaeb0926562f34c8e178d15dc2813198e55e986f2c69aa01e10606c8d9d883f5d8acb1508d6b5e1c576e123181bfa8dda8dc35a08030a3a74e2974ee19b16f21f300a8dfbfc11;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h412d2bebe7b5e8c6d4f72d119a8e9fd03da7077bcf02c64cb19db28f76efb83332999694b5c9ff62ff5db650c022a38b2d62306693a0abf7c2ae3e22bcf7f630854921200b1738c78d3c965f56f1c88ab46517fbf641178579fef4f3e5023190790be674008911e8c090bbd3cc209b7f841dd12df1881e33def85c006e13a374;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81232cb09150de9f7bec2718ca161a34d64b13646c3d5509688ba8d3545ddc52029e85c397a8375625a1eb625c8be9a1716e6c869ca9795e30171640e3da8da3272fe375458cd94b06d43c1f1434070aae7bc96b5ece08773bad32c50d1dfa99c2ece7c86ff3861ce790e1cc31ec2ba2470478cfd914f162566ecdd6003f392;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e64617e999e8ec1bc50344660cf3c15a4bccf529f029143f8ab6cea6cfda96f52f52c78799e7b15e67b1a562cc8bca1da0677bcc5f1a2ac6a9c97b30bd9def81418409d03d46a08e285024a5e689c99d35a4b29ad557e1381064387484e09fdc18afea0f15b0bcb6f10b399b2f10d9ea11aa61f2bba8536095c17fe6460f85a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6300be7c238038620337b5c57d09b3d2b3677df22960ddcef864bf4b69054e43ebd5e8ec746b5a4c4787a531b564b0157488c81f2ab50d2777e94b3fec8776afe36d290f0b9fd177b7c96d4d5c8778a0c07136b2512e187474353c356a31fc59d86c7c809eaecaf1e84758fa7793827e1122a41703ec560dcd0136c4fe222f05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc4d7aef2b7bef87401b79fe8c15a0ef328ae6d9822330ab6ce4e31b43fc90994b727990ab4c2f8ef32aa75afa39b11ec58d5f6fa83bcf90a11ddc686c23ca9df986b3ceeb4dddd33b1a17f5181bdf81b20f43165908d552012712f182ac019ed631eb20ee5fb07484f03d62e850cc808ddd4d63c4223843ea0f267290ad3e43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6888c2979d18ad73758de113b4bb7ed03182b04a4459ff7b12cf4e44727278aaedfbaf89e9db6219dfef3f7f684c872955416634f618305d55fa6e3093fa3fa067045edb118139b791a7616cddb014ea567f7865a6aeaad79608534283bfa9fb300ed804664740b1e1afcce7c3961159fa7385f9ab9135cace17d62e2683debb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77237b9d987e64fdb7d58b794a275b611c2f50d4be973ccac21fa22dc56ea610433546abfb1405891fac27f5fedd50a3ed8117f0e76575aeb52720078533659fcfb15bc202a73daf422bb23371f3d9e4d35fac9734ce6994cd869537cda54ac45d3cc1b9f27786aad2cdb5508a90544a031d002ea7e0e45518fc8f1a6ace7768;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he98638e082b0f675112d06ebc5a42f8f67a84d1025d5710aa9c02918ec185069943928c74076215dfd761d8a1e6c5a7fdfe6b1c41c22ab27125a29eaf93802994756bf259b1254e5254318302e077e232b25b34d6b6c68bec71fe8ce4aafde7744a3592100a048c1c71415c22166b5766855981312ce190d6cc5b5a72135967c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h523900fd6caa4265d01ed08c277ad81fd52f893b471357ddb131555f1016d431e0f059f66d89d803e5a4704497d75012e09691ddbebc769fe9e7cd4c428717de58966b8383bc5a11f0629e820994620a03b9016f4b3554f910c390e103401a19918498b866ecd792151463236874ba164c6c76fd9a77d7d292704056c3cdffc1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ea0e0e16977bd479ab17381b1b5db7425cc2ba798417ba3af7af85555ea65af0294fb76f35924137898582877fd4e0324b65dd76ce3d38683bfc06a931768c87b757efe0c8df583d4d74b40841ba8e49f4d5a04d3e8aace754ed683f67d22bbb697b2d4fbec216457c188e503f4ced475019d54a91471c5ac799e9427b2df94;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf66204fd637f64c885e08f55de73ed815b36835a25855910955fc5aa7697e5be6d08c3f854210583e5cc07e6104f3e8816ae6cbfc2c60490326de3fa95a35652d6955f3e232ef558a949a9949a874da173994e05f08915b9feeab630a2c5b79849699cd602d9bd5fdc47be217f93c5214b29c0d82d1b73946289980cb23f4381;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h445f797bf4681f4dcb6d11cb3e4528cd921e2b442cf6ded6fc74e212d33e47ddeb2919103c77bcce4fc1244cd023b17cdb385c4b03a6edd2ff3e18209b7504b4331d99845fc38b6e7ad40b0eef9143b561ab477c0853a918ed93ee066d856e947a5a11cd4f2f3cf4c0cec7dc5af34f6764d7de2d8365b88124d84cea926d841e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd31a4df7d7881aa8725e180612e897a6e5126b4b22260dcae8562280c662f0606d8321f3b35ef7ee4d4252a61a4333cea46d79443253d8a986c5fe013636c94110688d4bf784fc059df7292aab8d7be540cc173d7181086fcb95fe027b529c2b74922387efdf4de740164ae6a565583a2d3d82dc58baf46043bd22521e96ccf7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h371fda61e3d5be4543f7f5d258ed8d811ba6d4f367c823efa4f9f2f0474048aa09a3f943faf89670eddd43fb3ef5f990bc4ecad0734b5960992bf824b85515ecd7cff33f23d8e7307043bda9a417fb16407a7abc84eb9b023cd9d4a1e1ce4d0fc7f2ba21a67b83ed6ef7e231e1739c7513c77275a1a20d1f16299b1a4bfd15b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6d620f5b3311ebb45210f7ca049b17208387ba34c9109fac88a3c8ef122c48d94fa9fd5f6407c091c0cdd401d706699e845a55895e6f2dbc43ce8d86360c391ff287925ce84acdd702973461ec6654e132593ae52f91a79ea465902d692d639c10d64c021eed30276be93827525911cde01d24233e52aaeb31accb05c19491;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bc4101823eaa34ae5fc37816ed546ce78fdfe29c92028a2271d9576fa00736f489bf372de16e9dd69775eee44169668e92473539121647662eb1f0f56aa79d38c75b7e679f0ffa5be8f2c90e3f91d63e0537f61a7594e82f4d661bcfcffba7156a68d252c9424c16c8770171b030bf7d8b82ddf55140fef825fedfe70505316;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60c4c5d3658d0e9f7df7973fa53248e6f73f380146b8ce4edbc15e5359fe4a8fbee0a6adcc9b3ecd4d6b4e65ee4a2f7c3f742cb5333832818f38e151c44bf994c7a22db23f3ab973356e91544ec9aabeb87a2ea29dcc62a8b77fb72161b7a7ce0a0f7b992a7894cb128064eba0dbb48af8779fd0812cc083bfdc008ef07a1d52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37ad9e8ad4838c32dd51d34797446569caa36108b310f435127db6153902d5af215c298d17d74fde1e4c87b56140db6861c1dcd0198448e4a095338af2238603735d5a5c2e09304940774a98f18d5a36d7f1f845acc5f16eb5ec5d9d8db974f7119556b6b9ab416f5fc7b1a7b88ec8e942e2e9cf1568510c65cfb2ee8c992c6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67b44e8739337960f8350633bf8d095893ba264a55a54f2996856ac71fbe4390b02db4e07e5b503ec95662f6b4a45fbf985ff9dcab1776655411b176855a11305f5942ded889ce89671d6e8035370bcf9f52f0e91c515a1c60e7cf000df8a1ef12cea54515a0039e20d6416da6eb12a7bf4341fd8add551d3eb0c5fd4f1833c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf02818440c8a3f6aa655f0914c165f840f71dd5ad875b90230f82aaa0f9adf6a9cdc560b291b055781828518664183966ab40c605c7c8c3b63bffeeb46fbe0a246e5a68ad244960f9fdeb36e7669c84b488c942737a0a8b1234c621b3cdf16c916a0572041019fbd8d6b367f222a2295df38ee1a9bac018d612ee0c6e1c68623;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha886681c5a8b1a6c62e28eeb69bbd45af6a8199e2885a41d82d485b983bc0ca29f4984f2647932bc1090417b16dcbca4840f43f3cff1c394b3430736ce1052a35382c0d3c143d37e03a7ef8b67a066a053f03ea356d783e47252e0c3978e0e8cbae2f8fce14ccfb3e0faabbc7aff75ab4c986e8254ee9805ad6c9d720ff471d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1249ab1455f988c1b3b008a713375c7b1eb60e01a2084a9ed6fb0a90283fd55be2577774cae60b368610a3919a04df3903b7750d8e411fbb086b179b6e7e1b002082fc1d38656b8977e3ab2533905a87920ba62822eb782e432907ac52c3410e081eb827715d5e3978c05c897494d368abfb905ec95f6b87be4df4a74748ff01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8622525c7480734c8ee6a1d516b33102972828137bbe5b07e9b643e48fe60264dab3f35f890b0452ad09d100f30dccb72482f63e8a11e1a567d0538d1912bd577a1ecf847f2cafe568850e1f37fe625f5638440944083209e98d9636f1c3e7c92e972096746d50391cb80b206e64f0e8ede0b84f28ccaa4b719de4c544953f74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ffabeb2a01aa1a55b8b233eb60140a476f96eea7874cd0de9477802bfa9177f5256a79e0b1160dc605877ac86648d2864e7fd50e8ab8595d4d8d841b11a6416fdd4ded0973570b00b46c72b39f73edd738b79b78a7c532bb4e4f0754b11df950bcc4c6fad735f19ca7ff05c123aaf879bd664d3bf5d9c9abb04736b0923d203;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2af50aeec57ab9c9e32ae5e7b961eb0fd325db2eb5c09035d21c72a32eef3c49037a37410ca6d98c8c2ebc97d1b8c84eea2eb969bdf211919ec8bbf3e2de5df696a3b50e080b2756c605039b1b436907d0d478e9240b485022c56daa282947613bc438b35d37653539b30a41e2693ba83dade16740304b2e787629209788521;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b8d0597e1e220411201736ac838d074980b9e5093801ec260ca99e0d4aad6c5855d0678460053c1fdf2210a087431c1296f25ccd5d8cbe14327037bfc959e6a7abb73039cf0587b4d231641fa0c59264f19ff2c7962a0b4bd794fe0e3c7fb6dd0851f86fbd3e87b708a8d8e7bc50bf9cffa735859b714b27d9b370f0dee64bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90cd1166e7fa7fe9b5be97d1bbaab8c838fd5223b3e8525e5c42af4ff9da6dfd9b244b3d93a1e745c1f2d69639e324976a6d55c014be7803c8e6e6c90637df93bb90f8ed3c380f06355a95a6610923559a2ddfdd01f47bd4a37c966c04fd0fd555dae9095401135923d4d48bca4a52af698ccd9fc376fbf9e54b894f80acfcbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f05d92623f902e5a0f4bf42d56244cc0267659dd1f64f2f86026269f9b34308ec8e0aa443bb5a30ebcf79bb6126d371d470b209559e48eaf3ccc159f8e5ac0786ad88213c1cc3eb3c223a01704ccb8874cc2951eff6caf2bc85817a6c9c6883258ecd08e9b80bf5eb25f0ec1ec840a62e1223e1613f21aff04da1b95955ead5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a5ad43fb19e515fc19fc32d47d90953f92d317b4d57714a97f8e8fa7e348045dec9a857610343fd12afffb3d96b03936dfc9dfa65d26a43c70e1de214bb5f6e9b5f49cc0efe8201f3807f9dd4de0b99d94128977c09b48b5030400740407c6515015b533e7a710f50f3c5b152e5282ef90e545c9de1b7eda8667ef70d53bae0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ef248a86204492552cc2f6cea30b0c6a18d435fb7f6a5903d75e87b5de4d4089c75dd0ea80bfa8b100bebd6cee727bdc76679890afa9da1cd11aa4048e70f0ac283500b382ef63519691eb70816b6f551a2ab4f0d5d4cfe9e63f5b0aa248d22b10444ea777b7c83f56133ec836c6ca413ee2a43fd772ad2ac29f69ff8bcd982;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h317f456e2410f8bb6e088805e34d55600fa69f0746b5b899bdf266979bbb8001def99cd8213632907cb67faa1613f3703435862d06f3b06c7a49d53625632377e3101392f52e14b5ff8221b6fd8e94272fa9df5074a1842152e5a10a69d4da0d48f94edbfb472b44214d76cee1b6ee7d3b57ae01ea15f51d715676649a8f8f8d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2903ecc116fa87c30f4642b45e58141d13edad16694a935646e3716b1a1ef6c8fe87377399ef6927d7bca011e98c28e4671fd7f08d2334915465e752832afb2eca9ca20bf073020d69cef810b1a86e92b3de076a9b023ce4bcc1015e8b5333f792862c5f2026644c375871be3610b97f51bc505da7d8759338ee3c4b79a90f18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b07445cfa69e3521b3b897a6321b878ab852c06a7753acf112abae772e090df38d8eb40690ced1340014f22c2b5b6cd8b8d8adb77b30b4e93d86aa6bdaee04cc12f02619645bc3bee138aeac1f9b98094d07416ed2a434660349d60ccc35944244ce0ff32b085c9085f3aaf97d78967b165c60c0471e8e359f7b27b0bd0fa4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h818a471c0dbe2f0bfb699a58da126d5296cdc362380f274c22e40064b7d64cbfc9f74e0df357aaf491035257c31e9bc6f84638037475ad649bd50fe66dbffb9a58da6da2957789fa79097f9cc3158e998a97fac9e78572e2a338867fca57d315934648485c407d8536709b74efa094bee710dab5c89857487e0588cf72c07e68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5a2497ace0e692ce96a20f7dd4b45648621751f7f4837358aef8b9bb9c16918e8509f19e52c68be469dcda521d7e2d98922b06bbfa2a0394c63fd8b1d27aba504e6406d34f6fbbbcdd526e31aefc9f5987ce192fe2614c002ed009028c511259876e0044cb2dfff63a492fc73724e4c62af93492b7f9428a13572388619c252;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96714ab76a71c7d933929fd4ac7f080b4475ba1e856801275f60b898d82ff4b07975cdb63a2c936686caa53365505280b427a14bedfee3b1c3875d6c088810e09e3ea6b7b4db585283e561b615dee1cbf0a7bc946cc55ea4c9ab552c48e41a711c9e96e6dbd64fdc5b68b188722c6f98f7cdcc2f093ad896466ea24be0f98a54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha34f76df1e385fa50d07f1f58e8dbeac3ad16da4a99525ea5fe823e0b357d14b9c480809c23ea8239cd67bd2f1e643399d18a8700e752513993c328b08fbe165bff9432d4a67a3b3119a4faba61b283f80d0f6a201bc140e253fe3e91a21468d3df51c2ce48dc5e2f049245064b39a1c1f3063e5fb19074b82bfdf7e54f7f186;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ad199bd082fadbd6ab1691fb9c845397b6993085193c28b8c2d801ac98c529831de64f0dc0db8643d8c9399864afddb9a70a8bbc6dd08e252d612c9d27ebe031d659aeaa8377de85a7957fcf7bb6a8e968747dc0f62191af93d42eec2b8efcc34c4e8acc7fe5ae93c0159399f1e88646b238ed8e76e48625e1240be9f3a8fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdf4c222acc27052bbd389f8666b15759c53f662f1b746fda3a512fcccb89528247abccca90e9ef1b7afa529d82fcb54fd1a7a1fd28d9c990ebcebeb92d2708d7b4705d8b5d2a1e12c9a58fb65d063df80c0a70c15715d6779b7d6950ad50597936c3ac5d65c30cfc86c8ad1d35ce2acc3502adc1b5d44f6fa1fe51ad739dd56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1491544aa527743184f6581621b58416e1e075d1b24cf5f5c359827673a6d0329927a1153b445ceea24b0be0581e3c62101d03c71b7ed145964f0b29d25cb1d8a5a8d12d8be1026d382f5acdab7dd00f15badc8e1083c456d1468670cbf81a2a0891b25eba312d33e93124a62ae63bc5972652f3071b52c828c5460bf778ccc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd86624e6d7e82d768a055f142aa21999184a3575d54598cbd12e67167b11c062823dbacbe981ca963c18c69b968467ef030761cf81f7419084210061f2c75e0ba45f513fce12c7deaa0a7900241e029f4a59968b3dbfcc5887523817e2760b70e241e73e7d543671f361281e1372d5c483e402c2b657e4c466c2ab2affcc432c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbeb4ed895c386506fe1cc8149a431a884403142169dfe19395e60e41f4447dbc89bee94570f34d811cc18d34f48c199bd90a7cf9f2633909747af5522b77902a3b0872f99b80759dd39d051b2bd2afc3dd86f7d8e3e30cf90d3678b929885eff01675dead8948b4d573aa9542e6a1719fc0bf6696ae6d6cbd859bd7bb89e8fd5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf499ed88f5404dedb10715dc7436b5c1654128cb1e7cdbc6db72b9d762f406340a11d2dab23d07264c774e2fac26985b75a9dfdf120db7e38b4a10702fbb76fe82961670372b137c8b2f13c1b07b2e951ce707cf15795e414557752ba0c05d3f48a2b7b715667df20ee037145f73c2875b793f54e3ac0d87c267f56b0779d9ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98e0d5770695a681cb8ba0a704c6f144ef2e9e40fc8647ad3cc66c808435c16e8e56d3545e9d70a61c63db3150495cbea45ea5671761ab90d6d1cd0f94e369d4a48bceb337f273f392bede9077fb0f3eabbe18f7f2992f373d3847d12912ad608bb5b691331dbe75966b50c9fd4dffab9996a7fd0ba36d3226761a52cb4582c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb97bec40847b93932c4c4e5d386712829bb89660a3a62dadd319e6315cd55d4e9764376c8967ce6e8b61579c1c911ae88ee80e9b62a94afde2389bef68644145363c935dd34236bdcdbae1d0110786ad0a8239caf8fd4a262c361e57b79a28c33dea1d7613555b762a0f00798111e1945600fd751017c4fac6e06d5fd58e4aa0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf74f88085b7aa71fd699cb21627f6ea398b1da8146539242c802c18542a44d63836e8a711718f391e8338da4f9235018c0a7c8c5af500fd3d16a859641733dfba7fcd7dcecabf85a0d9d18a2f27f491ea871f6c41e3a0e309402fbb7095e11475d3e2039bd6a7ebf9810f5258dedbf6c4ff809014b8c086b24dfd5e747770016;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4489f1d131d334a38ee8ae88bf36c955fe97675c17f5d960496122aabee291d515d2605228d75cba26dd411ec662d3bffb2361c85b22fa60ab702beaeb31da99b24502a539150886b52ba0b61dcd95eb10e013b1dbd60623de90d847329a9b307d0cd4177707788570f10711f4ca8b6e81cfbbc6d6b1fbb9f1987bada371dab6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc074553d7da4f6984722e4b98592ab450a8b895b58ec989636499ba7f1eef3abb0c8c3f9e8937e8c1cb6f376a7e85e8bb4485fddde224c3d94766835e525a6944171b82c07faaa5133d081ab2dc379d8c2523c08ba31ee7a9c5b0613fed958184e908802a7f57534aef022e7a725caabe9bcc769a0cd111e31185f9167bf6d2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1c0ebc2dfd954215d2175418da117a7c7d8154ed41671f7b1fba8558ed3f9da16a94a8088ae6c591ab648908cb586627fc9972f4664dd428ddd8ec784cfcf91722ab582d11841e74218b74285d05d00d964b17e6d4cfbcc309488bbf470ea62994db2d811392345b2f706602d2bf94bf3728bf3e7c1623de843f1f73ad91465;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d4ba97c870fbab95fced7180f1f55dcb663fadb1fa2a5421d174373e6fd6f211b74b875f142566eb60139227b6144dad764995ea9641ea1148edd865cade5bbf75fe01d41f4d8732151099d9c681bb61e89a242ac0d02f4afb0ecd982be14244b67b5b1a5eef8ddbb046d747b346e6f27a64cbf2bee2cc2374aace35147d1c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e1f50c291971e6944eb331c7f87cd7924240c168fce3ea82eb2575eee7c4cc80e7a7c8e50102807535590f0de2355f5197980da32c32b800899f8c4f35d2c8e9eaba0c13fa70fe3958f711812559e4e9deb1b6dc859fb2079d252b663dd2a22d8a4f439f4ce493c530ee6f0939f6df263c19afce6bd70cdc3bd63ad87a3a631;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfd8260ee4af1e4b96f5251f8be63bde821ecd1b8e686e7c5037def0c4e8481524d431bea7806c3550ac9c93d2d7d85b65335203db13c3db67d8a5be5d927e2c06b5dd080795e099448aa07f65dcff7e02e31601e4737cd58cdbd2647757bad8df3afb902db76e2f2bc53d6ebe27a647a3f5e926dabad00feb0a98439100c5e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bdf767b4fad3df1cf2e6ca1b3c12a6ba386d99cfb59d7f11106d9d507d72f3ebe7214c7f8422ffcc276016caf29d7b7696eba230ecef01dcc53ca88c4a75ecd172ff2c33155ee80726e258e693f5430853e612773082076f1f08e959d117da665cbf381dacdb0907435bfeb0aa55edaed42529a45a935692a470b196a0c678e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4d78765bcb5d81fab8518a386d2a2f3583db2d9e8f42bc35080cf920cc839827077f7972787e048dec4282309250b4a0762e778a0817c3a1c3a0792b0f36bea091a818e52ff53f50fe9736fc4a2332898cc3a57f507f843fcaa2e7d8e7a30fa7243f7426d9c8283b018512295dcd7267564d5e12754088e5d31a5f435b717ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23e41fb2b93f2d7bfa3c08dbefe7f9399b9f03b7301b12a9f8db25139c4d60dff0b01e9e69d8870a07b0204783329b36c35424a7f213751652e85c8dc5384f316452775e9a7e8b6f4048742b5aafb2f8b219adab4fa0bfc0a9a0546a2adf40e4d3e81dcbab76acc2c3d867cc09cae0f333527b2db4a5baffef5cc94fac4e9ff6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3162068c1b42cbeb4169771a520cc839bdd078219645ad3926888b7c8fbc16eae8a4267df1afff799a29703124dfb4f4685ce40175c155a5896e954f8d8f6353aec664d8308c46adf7850b54ab88eb6a26f2e9f5d1a083790577bed6ab859760b3334fc0c708277fd1bd4e5d01cb79c5e8cd6cd83af4cd96cc3427e47d239f16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf7078e89005ff48f681f3f62b30017230c115af0cc4bec385160cccca206ed54f41ec49bf887f420d7f61736f0d7f54cef0b65e0d514008e4a8a28fd04780e02db21a1b8481131b92ee686e77d73e827c6c7436e83010fed03ad58c16915acd59b81ddb2b138285eca73ebdcd778ec250cd0f5357f2502e823cd9799e857213;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58df9b548cbae1a267c019f4e920b8675172f231064c4503757370057d8441de73ba2ece48a0718e444437363ee98980b60b9f8c8daa9fb6587decb0cd0fd6535cc0d3ef92d23235520c3bc514ad55382fe3de8bb566f476538799aaa77a051a773d634b7db68597b7fa680d3e8a4921cf1db528c91ac759e749727f5694f775;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0ad82b56000fcf6da521d62e9e2d17cfec5db5c70563aad9d2b3aadea435c7eb19d790d61b9eb8a4e0fd85034c697cda177f0e172f61300ad5fd2df18f52552bf3257c07368fa558d09d673614de3455824cf462bb724c1cfe6990af8968c06e165a57343f232bca48e3963d494b01b0fab2c0c23db3e93bb168e756d950fcb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6154003f87b96ac03b868777aecb0ddad7ca2c34630a1ae2c4b36948a6261f34f6541ea044ae8c63c49ac7276df9e1dd093885222406d109ed65ca0e8526a15a917db0dafad46c8c78c8f6f36aa66b3fb49a985aeacb936d151e9fe24aa73d91bde2754b383ec7fe113b8e97d9978ddcd5a1f508e78fb98a6d94b4c0c31a4372;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62a12523c896f55b772636217328025ace7c5914efeb8182376d1db2efd3feacccf7574d207262bbf592f38fc846bb8ea3445fdc5b76e91fcb396d4246d51e9014fd218fc1f56faa04c083d17e9d42319de0a24ab9aa4bb03b95b36da1c4e7eacb285289a24991eb8a28a8b6d2bd570af465a2503485f29264e1617e97bf5c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h282a407c5936a6d8bdd4cbd1f28327feebbbcc152f51b4b78f415b873b72c9e89a0a96c07c598dac93f85c5e7aa584774a059aa55b24a16af3319bbf8e21f930906d21e06460f7ceb9364c76b136d8a74331483a233265f640aba61e1bb202b84b0f5ef4d1e950a62ec0cf6d4f4b20e24cb24dae2c85b2a832b5ccde54392a2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82bb27e2b0f048e9726a98e2158d409c89f6e5b65caa021641f73c7f19c260bf8fcccb0994fd4a621d54fb8e0279bed4b5cb8f91aaed067d33efae92766f167478d2ee4ff01af1080cb415617cff8656ed7dd78d4727e1edfeeaa804d5b7cb2912736ffebb107a49c3883bce498fb0b8cf60769bd85681110a02674755ab7452;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f3faf1fc8785da7f7304e5f4dbc7be1c53a89531d470a78bb9fc01213d206a197bb5da3cd024c6e9256aa8b662de1953f5a44dc8d8e09e9740ea554c7e6aa86c01c4311a1904661fd9d74ad84b2570d3ada6023b0e3e8c0f0f712177d75afe779c674e1c2ce998ced5f97ea8679a1ab78f9abcab684a149342bcacc36e8963d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefc166c79bc714c6e10ad07f99bcd2e2dc4be338996740ed1e853383f37835ec1369353ea14ee8c7b1a73f125622c955b2ac09c741ef0ff3f6335403d8ed32079f2842c0ddf0d3f7d534566533a5a553ed4598e23bbfc18e9abd43e8196e19b3807bd93a3282d85339b3332a10751657707510b09506c0afb28cd022490172de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha18cec5ac309ee8e91c1e747b1c3a9e10401ed537d5962054b6e52035bb1dfe6c660baf60f8a5444d1eb3ec593e199dd068822854720c9b412a23ea94ba1c87bbea6a63583b5fe495bd7a5ad18c15a0419428451bed7af8d809b5d29458a50a630ed42b54b79d01d0a144d03c94a8a3f8a04eba9bdb6f0e124088054358649fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb65f611733af5454bfe26b886318288e448dbecac2660cfe87ab7a04a194772e7a90d372971e2ce8f6b73cac99a9efcf6662638117991e270b8147ccb807be47485806042399f6deb92824dfc2a07ef7b09505bb573de4367e4cc5017288ec2e43db1b841a5d84dd55105b1687182af7371ee5eef4d2a6fbc11161f9d77ba9d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65b6953fe907a13ac5e3b54963f92bf547d551ed4231dfb984321790d147c6cd83eabb451c319eef0f4f460793b090061af4b9a7f7a5f3d5adf8062e6422f61f26aee59b4efe4b77c4700cc50c74e5b991ccab55a97cca41378b2cdeacfeae9d5cb6e1aaf75f0610f6f828999903075192d35705aa1cd37733d9a388edce5be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd13054672723de9cf9cb5892c5d0482be6f3b6ce2f716eeb89f9226bcbdaca98bc6b6212fac8d2b6b0c05df5b9b8e9bdfe1164515957e0aba513ba68074b83695b3a7cc79ccf66dcca4f6b1d0945385005c1daa7ab8639c1a04da172a4dd27703a52268288dfa2f75c5280bc1c5f5e1637954979ed141cc9a3ad2f261279bd60;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65516debcaa165ec955a8f419fe396c7ee353259257baff503300ce540e07bb5c8994d1aec8633c412a07d2b4bc435feda81bed2c8fac6296f2d6dd68641fd581bb7aa186c417c4cbbd5cc054ca2eb4ca3b0ca7293c42d44301074271c9df989012426d34de434c73ba3bdce62a59de52ee24825ea7fd843d522898c800842ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h270ddbc1ffb067e156757e425a9208d04c4cd5fd939e453a85d3b612d0dee20d317b23d075ee3cfde05c217ba92ffc2724736431ddf72a8dfb61ccf9635b042b6ec94afcd84ae3ba49d5e4e1102603816ab8e4edb565866b1ba5fcd815f4814a87c998472c2550bceffb7344228c53f64837de65f383e4569395e8d8db5d54b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a54798189d96eef1f7908afe084ec8c18fd55235aa2857879a2c35189512976c4b8857f913c9738b8fc21a363718d1105e46db875926784d1b7c25d3729d92072ef2ab14d31c6e4cd05b8a0d1851f1f06cb5f143c74fb1bb8a8d0002e23b2923f991173c4c0a089a20ad7cc27cdfcc6d44da09966a76db9f6eb94c8e883c0df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h193dfef59c21dff9b9ddd0b855356dd9eeffc89a40ccb38102d714b2ce8794a30510eb42d258b3fe711360d03893e424f284275ca40ed8f1f8d0b1914ea1cf1b22872554a0ead186c560b6c1e3b0009b41e0b0b8ca449b99ac9df9b01e57dfdd0ea528b910eef7364b8c931f69619d8f3da68b4627dfcbe643119198b5189df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he412a30e275fae0c4f1116c2f39c6aef94f0215108e535de36ed2787ae28d95eb38053ee9f04238f4960645b4ebfb11b3b57e21bcf50f740c6896c7d36ddeaf4f97cec89b03cf563edf95f9da02c914e9a8eec108b22612dece23b27b65c1cdd2667648810a659543b8dad2f07df0ef4312382504c5e6e4baee813310b92eb03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2780db54053312f45a9bade8b86c217ec15d8f2b57d322f18895505d4d31d22674d73767d90c9e0edc65d5535e2528c15fee2eccf1f92c57a230659fb187956a3c9306e0e8af750ead47b48a15ba34b2edb4716c44f2d2d6dca169ac71c3f11742197c2a7d893518df1956791acd4b742743d344e4cf449c1b2a229a76cc05dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67e8d9d68dfa834d62d660eacb6996c92fa3c2718bfc9dabf1bf9eddc1943cea0da5ef87311a7027562ff25ae61a03ef5bd4f5a7680fdf3feb89151fde98a761f27726947592f8f676f031089406669d86e40d634731099b7cdc76dafab7817711676a0529d1ff14da49d991d87fe926fb64edfa0293bd2d653dd33a5a7b7e0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cf476462d5dd6428a43f1f958d1b30a3eccd952189e80649dad6e9215eb46e97672a41f04c6e789d69a7de11cd6c44ed2872f18d4360df47f2ed24647ef9d9fc0d58be9dd6d0cfc190f7ba57d4060470532308bf2c17b8244dc893b6dcf9647347bf624eabf27eac338fec6a12152bb17d40964575271366d1e539856e0e804;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9809266e7f2bbbf8d03274291aa65b9fd700fcc341e0c37562e3f6cf47104fe8f92360d8c792f4b99fd3d9bf45a0bcd9218764047550744de93479c759efcc14ba770e568329ecb73050ba5d613f26aff58b34740751feeddad587155b3bbd647db3249000a8e773ff15a35a7c8ea266784caa3b397f57ce30cc491fa74d4f08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h575b89ce62872b8013ed5bed5427f21ebb0fd14d38c6411bef152300141d04a34663f8cc927e5388d821de6e508565359fc10ae89a4a693cb7f90a1a663c0ff5c6578e1d885df9d37f2941686a9bd1719bac73dfa31cc9901b790cbda762f5ba4f4868c29203c2e877e27886233c56da72991e965f09d09a90fc77e437a8bc8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a183fcef1c073b87778af018aff6d0bb0ca9c509e7ace84f75e231b0860b82288786c88b23915578b177ee9d57a80b2961b28030b7362eac4d07a36c7967cea055735925b61593ab13c2a5b1632b7aadf582061470d6d0165a14bcbd8c7b7964dbed8e86d3f913f9deb6d2f34ce3683626896b2370659e42a29fb2687b6ff8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f189db324b38883c0fb8e5337efc57213aa14ea458e0c02e0c037037c892ae16405b32e033f985fde63dc0c749f26d6e8423aafdfa821f87affdc5bd7a031e8452065dd830cedb820158a1f2f3e09be4ee48ca4675a6710a88ae0c6feec6098c22dec04d302695cf0989ccb1b0883997c3afa22333bc54f074b8059eaf0b032;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf75dc9fdcbaec4c707eb75553494cf7625d4d6907b8d8dc7b04f4a85ca60bbb0b5d7e6feca0709fe8a311ce8295fe69608eddb0822f249219546285cf3606be6edc0346a0f97e94849c6852774359afe55c6c87f604c2f506042c81482623920db4e5cda2e3d20cf33b29fdf8a94bd15d63e0b394379b7142e0f135ab79847a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41704cde3f47ef44ea66515ce6763b516ac63c1e167f12c96dd21d037fe6013bae879f4b4b8deef19713b53a925a72eca26d28cbfee8a6d1c65a92fad44297c5bfc310ceec785e841fceafe9763f694f9fecee67ce4092cc72135756b1bb824a320f37edcff55cda79a8e993c2d90dbe6eff784e0d89b35c7f534549e32d3696;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27264acbece9cdebfd74b3f227079be8617999e915f5fe9b901a5fb691599592a120aecccaa355692da800c1af9f4675e22142303b387eb1c1b3e40cf9fc76a9fea8df95f1edb29b9e1a55e32017009a77fd87cc4d5ee7e17c5dcc536cd93eec1f9214321af24483a95241107935863951c23ae48aaeb8c0b6dee1e9dde4a5f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cc5265d6efc1116850450ce061cd8edbb1b987cf1e1bd79fdeae0d8b170f6af04cd5a9d7325d2f9d5b8132e9a6cf90baf8513fac78cbcd857bb1846bbaf041c409648b1be1930fce5acc7bfc3c6249207c737a9a4ca4aa881231d4582f9ebc228e1250797ab43d95f0c415faabd5565983154f4fea866bbff07c0af93d63c61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e3353fc32548454429dd55f0afc953821c0d85245924da1c76d6ca6fbcef00e8885ce3b0842d4f6721e107f84ad062d038e7d4aae2d95284a29bcb71dd802c4f920fc7998f914e1cb9f887dde0fcd6cde40161b293df60b927a6db85bf3746bd5423dec55e2bd279d865829ccec3535c87312ea9f2c4a5f67cad8e0a4cd77c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46c8704a3a74f7f6eeb7b53ec81956ff17564a3f74b567b9f05370dc8762b23231330f841f9a4eb78d20f9bb849b7358d4df6e232ef8113ce37abf55e329b677894a1cf5ceb1fd91e910f9eedd0f1ff56938e8ffb58979211260a254b55f9cce263ecf0d213322df66abde691f9913d439db9d91fff17ee1a7ed3d08a1be0104;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb1ced79b2be53e360844a830dba2d6eb1c61c2f50c1b8fb8cccbb647df09cafcebcf305068020af81a88d12f0d0611ee61056da94d5ed46aed0b21f6eec2bb09069eadf8ddb8521965509e3f7bda5b5e40bb5f769acd12797be144aac08782381c5f595a7e7a27778cf76c0e92ae7bf97fc52083e87c5671d1b3ea792cc0b6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bb40ab0b938ba102f71e4a354597c580e73b8c30b2d8fb86f8c6c1309eae4c8eeaee67e03c301f072250bc6cfea0ac955730486d01817f1ffcbf1afd8e8459380a0a6edf5b0d0d4f4614afbaa2278c2560444953e3ca79af6b44489cd996045f5ca1fe89c43927be929bc808667e8429e3425f7c9b3b765642b7ca982a78735;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4acd47576561b12086d9ffdf6951cc5968813a817cc04250accf474469162272895d20749c73844f8c4dd5c75e219a435fc1db21b4b387c18374f76f4db0ec18cdd864887b590c7aad75cfa36080a30d38dc9d8a6190124ddf948693c9b1df8b692f3a8f5ec1a958bbc37bbf858ce99cf9801945cc4f4a074cb2b4c1283e18a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb91dcc3f51d34de2693836c485285c58680de4e1e33a13390c45fdbe8502328242e4aad4a4ba0975614b6b06cff472bb051ae174b607e264441f37e766866c1df1916f015482d0fccf1ba05bcddf84046c10b6f3a1af7617a177694ad83cf98b408a2b276f7de31d4ecce6e81d894e3c7c7f8dafc9ff4b241d17e4c68d1c0318;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h347f612d1b9cff67ad1ee90b6224503d8d89654605128a390824ea4477a0f9b13da776316a5ae0907199c66554708a629a0a804fd94e9f7df7acb46382ae94f54e501d9072a3b6eda6dd1cb3c7530c3f4dec6ed1fc7ed87d8a812a685e59a019a028f5bc30ff331dde672d1e6c4f1f1ffe84392e6eb821d4a3191f152cc53cdb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5e2ef8cd2e4bf19e9a7b80a640450afd72fce7d5314cd278503cfa415669b21f1c13e12f8bcb19e603fc4c85bc0cf37c167439405df4b453ccaf65e54f42c84efcb3f039a1c134f1968ce41caf0544089604be320d05ad1159644456ecf3934c2a92ce0b44db4cd9c619dff4ffd2541e8cc3d3b12f64d274d82976e31f54650;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd49e9e7ec02475092140117993baf4ee39f77321e3c796ce1280a448b9f5732e2215eb884f03cf89ce2715a1e15f770710b86ef0c62ad32aae04a49274c3f64aae45ab17265efad6c7aa0d8786ee96b05e0e19d0ffc3f871d77a97065759135a071b6442c55ece999f3c33001e81b2eef869b5a254ffac8b9c1bc56e8e45ee39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b649cfef1a3d5ee5d26efe17f8938aa3cd121b840a2a91a49ecdc6f076fc01e84e2e8d5b04b7d7b9640a86017f02656307d1fd9af432d95418f54bf04de64eef6893da5bf3020fc350977bc1745e58e839963b0e60b4c6de060ba48e3316cfba7d89c14d906e8b33fb8c2f17d8af96602ae9109e624ae69888e871cc6c0cf1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf2f1f475e32dd3e94540d536da8b0cde7c75361fded24f8b384d0acbdc746b93a587410451212e79e7dc9bfda94b7be3d1eafd14baac663db43b1a222ad9361944b5dd35b7ea520aa83a262bc438e90f2d4adc2af5ff3e615e66a55befd821b8f4c6a672dbf0b9b974ef9007ed93001ccdd589e3f4907f0e9917bab69ba5ff3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h474b5f77bb7a9f81cd7af7bfade4e9b3d7e61d2acc6942471fe1fb269a604f765576a72b11cfd955d10264af13e4ad5127d1eeee959482c88218115306aee6a546d60645b739f4f76c61987f8d83806fc76cbf38c966674d35e60e00b66481fda5c9b676da250f57a19016da606e2126f2afe6ed210879b87dd76b1f194ccf17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9dcd52eaed0128e29ac2b32b659c3a180b6c172e2691cffba124afa4ec608a4f09d1dba6e35ed1d82145633777b6284c7755b41d7773720f802fc85df6961b33afee301d02632ac61609eaf52c3140fe3841eca9849c7709217083351bc7f8b6e69d9166317f0707f4aaef5e4a0c5a0a997345f65dc6b567b9ca26583494c2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75f5f0a68d96dfbcae4ae41e242520f7cc2576859b1cb766938741bb5fb305af30867741c713d29ec0ec347910ac0adb6d47bb61779a6543d2a9020c84282727290c2e306c5e44d99c02b29e8b9efe05945af63994f2e460dd34f52ad589121a36d75bb8154f14738937aed29f2fd58a516dace0abfb57f2da6acc91cb31bd20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4dad18296a65691bc4eae9bc68eab3e453703928e856a6788ceca6a3c8d80be54b6ada54da976469ee315148b7d180dcd41cdde21080bb5d3514ed1055795de8b4cf82651ad1a5fbac63ad203fab76c05085dc334986bb2de24216a39dea306ffa2c916bba89e8588bd49c6b47dc4b17640c978d1cb618a6aebe0b78bedad19;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b2872271b6b178ff29bf42f0b5afc10804d5b7db2009fbcdb1b11baebb1657cb19dfb1018ab44c1199f9caf7f328f69c92c7303ac9fcb188c60bfb0ec5b6f975dd685d906d0d5a171b4b5775be1c363998e8a5d7df36abe84e35862daf562678b32f9e61f001693efe74d640e9762ffd2b5b3afb642869ac01725febf9191b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfac737e3dd71495a1555b68bb4e08020e05292f256280f285f1a9638f1376571167ee92d1ddba3fa10cb1d718596fc10b292e05be0f647e1d5a4fd4dbd199f521d066b5f55d5e843299dee4f9a026b213ea545a51f7c5d0ca0b1aabeb6e58ddc753bd7a5f05f1c08af413576bf0955a650cd1579516f6ec0e6442c5e272b5527;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha25cccad031daffb972b3992dbbe1fb89e53c144c8111caccd87b445aeb43c5aa67728d5dbb239fdb67a6f0efcecf2752fd8a03183e702b59170cc3d9b5718851f35bbcb23540ecada158015b51bca515f105bd6c42d454950d5f7d7822f4f54d35a605d225b677f6f64f39eac723518bfff7554c023019cf4741c68f9b501dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c58ab19158ba43585746ac791138af15fc56e85f70529d0cc725e960d34819bacd6ea63abe2359ba1837005fdcba33379fb79b81782a3ab28e5f10517025fa905042cf22ae48fe778f63e40664447a236ebd38f0be63f66ce6a6390ebe47313dbcb243de71924598d62650467f070588c3b8212fe29776c2604bcff19fd44f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had4505c3fc0e991247f60af0028de50fb781f263daa4bf6cb1ecc288aeca5f5feec4c495b91989d69141237e25d550678fddecf32564454d94b87a9e5b5243e009dcc9a194f8bf4960c2d4ff4231424c58721d1560844a2cee1932cc32c988cc0c1fe9819efcadc1a5cef7596f9311a9e9a99ec181f5c538f389de0b8a1ad3b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2091c60bb922db59902a17ac1cbf132825fb7773daeba298c5da9d5acf303b21486e3a26b12e6d64eee8262aec1603eac7f819b612c73f271512f20fc4db1f6be4f7d1ab66d4808f678822469db7a411592484659dc08fc1a2f7f6870c96d0fdd36d38f60d17906e5458d86cb98dc3320551dbcaa384340233f34c7ae9052e33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf81bca13961db9afd9886d6bbff90aa73e46198cffc3b3c801cee490dfa1c8b836d8746b723cc570e9524978c8f828d66f174b6145f6a90dc0fb59ece5b44cb1fbf03b7e2341b40d5fcca1652aa462c7cdd3693f855e24d5b4bfb521b3e317c51d1786c1345f8a4b6c0536f722f50e65f80ca24ebf7cdb2f83d55476d0c7f902;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h947579086ba1cb5754320df4164092e60e12f9b31528f34689a388c06c51f12a3ba0014d7f893d55f938ff0287a9e8842aaf20017d90b2f5e5b9fdd2b8be9c100dd789763ced0a58a82815b83be6c8b9d5fb30be6f428bb5e2a07f9510220e1e9d77c2c8f64f12e6ffe58d68fe3cf7036c2231c8d97790706492f65d97c971fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he68ca00bb4f349bdf926edbd9259ed08ef3da5ac5ff20335cff275e2ab8cbe3371f324ff2f259ee699b1c5ff4954139b28ccefff97d4d806216ff053c1389136d3c763c87e65f558d742596b3407215bf55bd1e7d0e5685ae0eaa86c28ac8cc73da7a14449eaf1692cba4d3849b1706cc1e9babe885caca6de94b0a2e95f192a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbeb21ac4bcc681f7a0b479871c87dd09537f27781d31fca4a886cc23183c375f59bef1ea55643097bb144270e16c12e37cfb5f29b034a4961260aea40dee0453cfecea16984a46056ee113833dec98bb009876d51e1c442f0f3ed8b75273b54a185ef15d4632d16031ce8f9ccca8043ecf3f0a7a4756857d13ee940c340ccbce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h817b610eea609d6afc685c434fc31af14482afccb6977b35dd0c71644e0f5dfee026053f455a5543aeed067074f5310e6d532c0d6af515eadf424bc71330b3e92d394db4ff230e5856acb4d2a216411435cf8e2747818daeb42fe60840ea9534c6e00e3f814299b75c03b635b61304c9ed30f3d074b70a53705e698e3289155a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbabc9d877a7d27dbb3b1678635acf610c16e425da7dac042653f6282b5a6957704388bbc94ea7c613e987e600e77ab0ac719345f69f138152f92c89eb5a74b21ad6b7070ab17ce8e1ccf27ea5f407dc0e2414d28b307cf4f9b77a2bac1856746b4fa8c3c69a8dceb86cdaa0c232dcc479b9c34d5906517fbb3f639f63f1f4101;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1529f9b94027390ee642bbc1a384b51ed87895d8891a77d5721ce9fcb133f0ad673559270deb51c3a354fe7ca73edfe09c74b0ba24b58b686d263328b98252342957048fad86ecd90c41e224bcc45963a5f2bcffa075c14103eab699d59b71ec4cb005635342d00407ae11653c8db416831069ab04ac946e3cc259cfa31f49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf61c26d4ca4d2c33764cab7ebc9f0b4e070ebb95556d7a5ca7ce174155a8d3e78a0d0dab35631f0327228e64b7b6ca802dbbc9944b46fb29803005191f6753297f50f952c3f3c193691083740d2acb323987ea79eb7059f88b53feafb1bd68b6abb916d8bc54b1c4f8182fe8e9e38da6a7eaeee58eb4a00f967795d7cf063150;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f18fe180c7362918f8701265efd1654bc9752daa4dfdbf23fc2e18044b594dca58f106aa6d0d7d89f71030776826dc1c10756e40223c5cd944deb54d7084dab76ef1c0632f203d7a864374fbdca3e1d3b48517a6b13fe92143851057936e8e34efa2610b0e997ac4dfa748491ddbbf5b6c8f6af7544afcc469fa025cbcd7497;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60666d8e17c7241a47e8581811fe6ae698c31568d778f256afeb92df3aec526c4bed7a437f8951f6ea72292684b65815be13bcdd7b63b95f7949ce65fe0d2898d095094f66b1888234a21d325d1d6a7e3e46864d1776b3ead751d69c2a8ad7f4ee54f0bd90b3718dfd8997ac0a52a11b8b1756a89724f6ef5847c20dd326f79b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59d92d10a065322cf2a575634a052c1773f7812bb5d6a8f6c7a7c069b764bc7afab6bc9cf63898084c80e11a3745dc2d5ed82c0cc4b8636b14206695ade9e320beea91b846c4e436ebc09fca0f9ee1545c3c3cc55a0e7d98c92c90a5f8c7c16c4d6257b6b4779d12cc904caa5dcf7330113d1287006e3378f8baebd9a5f15d33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha992e444e29ed89c37b951b99797d6672eb483d62ef20f4602945342cca812ff2801b076bf4e5a801d2b201576e74b44eb1679c3277c22dc8c60539cf66af8dc956093f4919faea9f672dd098321c1735d47d0aa4c49b196253341f355161d3e13f20b5780d1ce772843b6c01927cd0313b380f87b1f7be7e5cb50c9ca5f7a83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f1c4532eef0ea6c3cbfad8757631e6b2a48f6b809cea1715a7b246a0b49fa73873f02955d8e3fc05d935f4334cdc85adf4f999acbaca2035d31c3c349dfbb4f3684fdd5bfa04f7bf0d261fdb3c58037dff55ba79c4f96aab8ffd2c3e5eb95cff4cb7c95842116d392fe6d0e57b1585921fc4c313938fcf9bf40330619148adc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9c24b8803b43a5aa10226f6cb9d324c60e33723aa16c5b055c30aa24320cfb709492e53453083f13368bd4391ed462250a98f7d7a48bb99884c76487d6f3f1a40424425de6966df1627170f1ee70ff3fd4c87be521c3d733994410267f0548d88a2e7a8ab125556b2f07648a5350b92ba970fbeed552103ca16a43619586123;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafbcdc55bf6dee6d5de44309210c763254c9bbdfe3221ed7d2c9e7818ed5737567de15c754ca35f3394149c0a6f2b362de0139303df61d3a65a3e7dee9531ffc831fd849d8c2465cc749e1b20cc0d2f63d894a838454d475e13646795b1264935cbce2c865746fac0a855763845c39b05e617b62bd1ba3608523b16fce161af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha59cf63292fa61ebc363733fd1c2553d8c89612d39ee6657f515e3f0ea4d7b380c0803360bbc8466e2212f98dea1c40d682592e5355d153cd21f3922e0a8366979562d5b2a02857084bae0303dfe515d590bfa83c2d4444502f170572d22448e1e4bda54bf38e90eb8fc8b652c2542786b6618e5225be3b1b17af7eeccebf916;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97be1faadc1f9bf30b3f50935edc12772b42bc036befefe4ae9d09ac6ee21d776963d004f4afa342802479c5d01f521e386ad1848add6c22afd03037e19b2836747d09444883c463e3e3efddb059815a11c9ecd1e69cf308dca731cb92f1f90d0ae4fc7efb3b68dcdd34143dab2e01e0fc4f0de3cd9569bc87e72735059236d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48a7f1bebc0b908a40ba75fcbee6fb2f8492b515283b0ce38f46688184291f867662be6e7e95ab1b75e8e00c02e9b00f7047b402476fed4336ade3244c84bcb7a96879827d90c7b551ceafdb090f176b62aab68e4f44c88d459f9338198aea244d0edccf54d684f3cdb8604b75daea470e17a1dc17ac3cb14b55dee2ed56e33e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h528a59bcd9459c7ecc886ad77569becf878daa005faef802de77a9ea735709b18f243b11137c0392fea1c9984143f4002c710f5a151996d320724ce397ec4d41be8398a8f22b944e6ba5254877bea2723c54421f063479a358617a93f7081da7724ec2ac61731ec68275127b6b8102c0871615e13aa2c4023e510cc525e5aab3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3014f0768ee7ab91a2fb44c82a34fcb96d4f8052fb324a5f6052538e45c16440ea037b1fb053be200e2b0d3b2f57feac193d089497994d5b297c658197cab5caf7ab05f9a9f2e919ba7e8935746d1901218d5e5907f97903d71fcb03fe34bdeb6bb67c7794087f0164dedcf09ac1d8848f4d63cc6b2bb3e60c2a0307b8676dba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff55974c958ce5f9e9b6ad260bfcf1e4066a792be5ec33208dd7ac276e58b98c07be42ce0baaaeed72ade262f03ef28618f797b72979fe8c934d5c6089c67d295e26da8bf0ec4a44f7eb666ad647cf764df419b3d5a7efaf6599724be4ea694e8b3e1a1cac07a76baf8f5d2fc11685e0b8e4fdfbde096a93dfd92b2fc23719dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h271813444368ef9ed5fb3b6f4dac267bccf8bf2c74660d6469a2947ead07740d9f63b03dd3c5cf11fb45f3893507e1c12ba2b315944795349d6427e8c2f1f4e1be562d4131ecd9d757959deebd5a0f3bc8b83434414c5329b3b233c107ef38b502d56ea833e202c1815b50d24fe34f7ab606ec38d2317c8b8bb3e0e7e45e8c76;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea6384a91611e87704fe35b01d9a422af49ce6e73030bc4eb6a296fbc030ae23bb909cf0614b75983b46cbc37e723b1566099634df41240e2b0b5421b7f5819fb952dcdf22215be717b247edf5ff0f20277f1bce34654e336aedbb8865ead1c76c8ef5fb3095dee14bfbab1156173212109f823151258b944c9dd613f134b4d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40c1ffc25614a4d9b83ce3eb767012262110ba035e6d0a37edd51e604565cf5eb1b8c79809b9418d832f924113394d312ef275cbd3def8c5d8f708f087cb091d07a71b87c170743a2b26e36bd551e18837b9b2390475827be02788a0ae91bd79cc0e36964e194a19dcee28ceac6a94e7a6312e70f5e2ad0c319fae0e8d3e8e77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64fee082f2cdbd0bf574ca177ee22186757c947d2bdaa0c9f5dd5c95c852edb307db83d1a03c3023f6a58ca744e62bf72d5a4b0c463a3a00d7676ead8f58073e0ca7efeda1c9b2e0d9f1a9ce1adc1d771f588bbf0db2cdd1b884e848ac37ddedda9a50af8106017b3f1e6afbd200986009f133e60a28c39d74589f6dbd0e321;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76ca409b2f6c4a5a69d59ca76af068cf7c9c23b0ad8a22ab40810fcd10d38a50bfe9bf60d5b909e04c09b6f3d04d77f7826111103dab87ce599c89d8e48c8e1fa615ece9b2e647cf3da864fe8e871329b7066cfd645683fe0de94810b2ed79247f3286a472446c6f003368d492ed0b635888c7b03773239b6be0f7224c7dad0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1da6a40d336eefa0ada59c576971a8207265f4b025587a837b715284530ff78d3d68d28d908cf8e047dfcc5e5922279cb8b37d6c169287dc5041b2b27e8c79512d6a77cf57c58b6789764d30bf43531016b675cd4c7a2ee4dafe33f2264376445d5765d946980fb06761ea228aa716df3694d69f2135f45401a09b435a69d12f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65958337ce355dce81f6fc0847e1da5b8d15408a7da26b5ac0212eb982645caa7f62c57172b121b41b4058389e278196c19305ae4369d7ed9b4a219b37adf3c3c36dad25276bc65ad3e61fdd32f9fe1e033857a56bbbe1d8141705d9c2e4aa11293c404284614123f4528c3045161534e93ee471237aef9483aad2e328955c46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66806b3077d59387edbbc34945c8a65547622212f3d3dedb314a9b4976014249cfc1a03f136e596e4b28359d11f8a59b92574cef1656e20ca94deab9262028dc39725ee37c4c9d3d17378cd0f285da9772c025e981984c2a46c18a8a144a728dcd335ee70598786090ea3af3ef7b925ef02bda0f8daea14cd9433411c4db512f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb8d1156476d4b6133e93cfbc445e984ebe619fc3926209738f57eff8bc10c00947c92bbdf591c97a01f7b5007ad13689d77c00f3c317e99576fc9128071f952e41107e115cceda9af2abb36ec95914d304ab4fc0db794580eef193704e1069d3c8bbbccbacb0a5fb71f0227104a557925517cf9ba91bce62f06ad35ba488ffa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedfa795a0041f89d35e0a6b486acc60fcce04633d488d33f74c619d0984c7fcf1e1b30e542c9f2058f21014a90df8ab46b3f0604fd300797f97571680a3e29118db268d090b794af0780f12dc32302ec8811983eb4cf595e8ac63f261da1b6200e0b2c99c3b5a9d333efef3312d92b85e2ead49db04304429163ed8fa8a9f79f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbca499fa28e5a4067e151b12d0feb19695396f103a20f14f614a2a0bac7bfdf0d39e6730e895aab3fc2cb29392b3d85bf7aa7bda789754fed99352e15f35039f2f389641c19139ba4a9aa5765ed09230e21b56305b50dfab25223eed8d013553562ea34e0bab253f9ed8fbbc42936a7f80dab7db271f62005dabf961d81421e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22acc56bcc309ed72f160a135675dced0cd1da8538280e178715c4a5f2f2ccd6170943f9423573e613908efa69c9e43da38b4a52482784466ee262c04d9bbae02162b1b20bb9fc8ee5bf1a5239db265329f5b7152a13b5d0a2f9ea3acad17fe4c46819e24f3f7d9dd9b5a029cabb7bd63eed8ba9c044e5877f892243ff3dc61d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habd2c4e436144e876f4be04ae12d205f36905925e31cc9c5ddb20185f49cf9a6552e3b61adab81e44be5ac8b56622c869e2ce84eabbe64764fe0c7ef19fe60d71604c7a0548b0ed4c9a5907b6fb8f40b049cfd54ae8aacb2f6f160a89aa76c7032eb98ab476541c9cccb145134201389bef2017b2c4c7f3e53dc8f09bf9d506c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h280e55a14e0b1756350bd161bd09ffd9d343c2a181fa30665df15f60b065329cdaefed2ca273cce1b3bd1ed91df53dcb5dee03e45473b6849ae01ce02bf7608d55df419f454d02ccadd3c7c537d842ea64b0843c96dcfe3931cec27a35ba569552d31c8a31cf642059d14d3a2dd2278a0ba88817fd328ed56b3f25714907961c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h283a2a05171a468e74a7792320234a59824b3c860f6ef6f841f5a4432775506da48ee182e21aec043931fd67060a43d4e58006786a65011f68f9143049a3909dc51efa3e122956c856a5d4ba8d308565fd35350f44c14f483cd9e3aab08ec169da1dd3dff70304d76255d51697e44a9f9da14ff97859bb6eb13f9d3da0630595;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d562c2112003525f17cece52045c474065d0449578822593ebc32cb0de3c1e0b756ab42fbabd3f59a0e3d1cb5471bc2ee576f9abfcbe86cff9a08bfeda044006a6c74a0d93a99c99a4ae045dfb13c50c0f4bfd46f02d9c34b2ca06fc701259ad1b0a139564299138f2afc95e0bbd80a36da6a43a6e505a5b2d1f41ef7e5b08c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec46ef4e9c26b8d9eef920cce05dbe7c3a217929969f0e9565250b8e51d3d3146f729dca10f354b6fb1d2ddc2776ef8b541bf122f0b1f777a1a0b69791c4d3a07ea83594030ee5ed0e88c75f97ec17caa0f358e3f4fb9afc7464074ea0a5a9f4eb4fa347ceee977f25ffab40715f53af519cb40bb927ce553d463bd6370645a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b54975306e068725c040e3830a4cc1b5fca210c0bce81b4683256fcf90db47d6ad898b881b8e6a9eb2c78d96b5e490b1ee2734c1313ea3130abb48add86920d1808a3eb86e91734a3446fd602c12735ccea7da890dee6b73a6b779767eeba3c7be384793145ec2d4812248b9e822044024ebaa2ef1bc4e483e2232a11cd6a96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0c60ac23335bc36b8962a1ffb07f2521806d37eb3c81dc292a3aad9af95871da8cbcf929d38a5880574033ee2ad2c9939879c35c3ce45886cd753a87207d5e2d88915c4380e4699593f58d9393ac61cbba004030f8b0633fa0927766e44dd282aa0e3054d50112733ff84a07169042f31b163f18cc5fc5a2824cf738139c1ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70f6f378d13435d1006ee4c00de7febe1cf4b5f9364dea8fb9dafacbc1ea1a226d9bacb12550ee8adc03277724ce66259f2338f4146e8a07cd6be50d336302bc3df0c7acce3dfed298a10f76637c095e55fc9b92551d607d1c35ea0f26255e1363c355750b80f4cf5f20c6dae283af5edd74bcc3be43bc48c4ad55da9c79dc7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf79ca947ea75e400d706e2a7a3aa348bfedecfabf171c938e24247ad1b2473e76dd45278140d29c7b4409ab10a6a27140c0dbd7b37bda7ce58fba4f4a75360b3a26e73fc62d2dac59d6a6b96e3ac98592a7e058f52bccc4048c3e522e73ec9d5a2954461e953dce2c270e33a3ea38e651ccdc5e2335e8b5411b5f71589789447;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf65344675d33839ca28996b55d7110564089e642c21b5a64eedaaa0b7a855606eb48dcb285879561888e0627f132006cc87ebbbec75e1e61a1cd153a54e6121bb141220476ed080254cd14f8090300b16fc516a2e900f5301916ef4bd2060d62d3ac3681aef9bd87916a70a6d984a09a5764ee97c9b89ba6fe9f7577bde34e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heba8dcddc6a28e38c2130d2e16f08820b05866a32b95e4509221fd99152e901341d5c900bd7afd43a7332f918586bd57dfde9190ed8620ca6671c80c31b8bd141afa2eacec5543d506c5e6c7f37acde2c01750aee351edf4dcca0d17f4e5fc004997ce717a0b2b53ac01a79383fcb1bd38d4d2319b7b6ff3cc97ebedffeb5aaf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbad86ff4c58a4f36bc9824ac25d3b85296ba9c0802a3e90bfa3c193fb88be435d1a0f9d5bd873d6083fa22c24c71f27f69ebb5124d67d5fa7ea41114d188e8a15cd87934b377f932b33e3fdaa0adeec4b38428d17cc830a51cfa9dfdc07418658af584396683b0249bc5d03614af8b13b93c67b1cdbcb29e8a8cbddc56e27508;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fdcebda39deeebf64e335dc03b59a106abc580c11afe3ace891af2e752277eb53d0b6cec264c3a67c806ba29e4bb0f550619d8ab5bf237cf6b8772dfbb6346d7c3dab7ee2d5a87f57bd3a28dfa606c6de796ef3fdbb5c172248431736208bb3411f961a1c67f2bcba9d95f5e42d1ed3acc525e19dec7febf87023d957421861;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5eb17f613917df097b60b793678e6cdf51a41ea0e521497026ed5fe53dedb29d4e562a5bda1ac3cb3dd2d91fdae1097105d90ff82e0273d6036454b2ff1e647abb7abf27fdb88978eb546a054f3fc191a0d9f91a5b716220fe0047de1043bb8cddb3f969b96be85ca4c1c235f30f98357af9f59799de29131a5071870b22fb05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ab57d3f003c22683bd73890f1a126b3a250984748b243b5a0e78a682713746c766b5a12fe5e817fdf10b12bcd01275062acc26421a4a4e5a7227bdb94ad525cd7603e075ec36ac7a59253621ad21c9ba20b64bb6d3067a5dd3b16b8804237b7da1ef349eefdcb8533922eb4126d195c33f8d1c95d3a9d325297c1d91ee3f353;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58d9892324196291a260bc55e9847aa7782a59c91b1b1381c9d48d72b44ab946eeee29725c27f4f2bf3cbd845a114c3f8f5a3b38ae7effed28bac338e4e444369be277c5e00d729d5cfe3a459d22a0d6af60ba03a16c9318f9363ce7a871226c14b7f96e3b38391872cfcbd8ae2742890cfa5abe13d3ef6b48af86fb03d80c0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a6c100909366dba856c8b00de00c56fbcc6bc927fc9954fb7770899be3588f80b5153e17e07d0e44af319be2c08c40de160534f986b5e0afb99a07aad9386f4669f59fa9b971799213f012f130f9b96dee4ab5a93678d6129c3c99cbfc785fb978106e26651fdcd7ee8e964536decbb3cef9a815d1b8455e9fb9be6f7ef972f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he44baf3d07e34ecd4460d9616c66b32a725c803bebcf95d9baefb4ebe8464d17345b88e34064848f493b5631b69e538f820ba89b367d4bcea2d6830f6a0bc6a09a3ce24b6b5588da496e7a43a305c9bff94052573dec4528b48e8292a2d60acb9a4d6fb41e0d6a68f905cd1135d0bf51d56321c401c40a5e0858f1dbb11b2175;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36978076336a049439b0ade833028c9f117c1e47c9deffc6c31f8cd22f111841ec4db7f3f9ea9e7fda35106d67cf682bf4606ef4d4a50c07b418d4636b0c052564613bdcc57e2c47aa7c1d1d1922db599d1863c0cd26410368de2c3126bcb5d5eacfaaf6bd3519567af315c9d83442bb19342a85c50dd843ebc1216351a20848;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e5dba5b06fa22d719207fc908100e79637a6e380eb019d737fca0abf0b631cb6617cb951f29a4cd9508da4584a96eb832e74d03c63964830ded4fda5ad10aa0b58902796aacd32791f00738ee0a76fb8d7bfe5c74a1bb45f5a7a54a0ffb1f571ba5ebb79c91c50c67613c188afb1181d362bc59e7a2268fd1e794a70d53f4c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38513e1b01d154950e780b7590d77ea28eb872e9d04d3d6cc89400650ce894a6c1957f3a7b956c421eadc385e9683e60b5e688aa28c4b2a117c9be702abb934fb892ec8b7984cb2a40cebb40ffa6b3f728b9f9d4117ae2b0030970bd80098fdfa300c9539c61cbdb56d145361ea83cb8042b700f37f092d1315d6dad1efa1b6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f27d804db13cd5e7aaf62a7e49f197cb6fcb0733922d09b555acea5d23974174c89fc248f555522b03b64324f95c8d7ee822a745d03067a61c9bdc26625d813f475d549cff011b7f02fa82adb5d39f1f05643219c95f89b2675c313c9278eae0af855e078944b355758b5c711a48f9ae6f412cddd0cf4bf782c3ee36baef6f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0ce1f11b00966d96fb6e90f3130a22d60f883114df8e2dd52f2087ae66536de4d3838681571e9292045a4f9f20eec694d859c2dda44937ef424d644f97a85e73542df8d445b1d8bd7155b598343f6783a679e44d1b43dbe15dc150f4bf2e2c3c2072d38d27206e7a2fec71031dfaded2dc1289c25eec4cbc199eccb73a4082b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddbc704c3cb384c7889bfb86d95fc6dfd99d79eb003d71ac2ed68d31d7ebabc7985d04714b8635b46c9ac26c32ff114040d59307f15ae3cc73dc7475fc814fcec22f75e64c980846ccf47cfdcd1520aa12e683c8cced66bf197fe711b87d51072cd231aacb292c0c57f5991ec93705a8bfb9009c8d1774a4c156f3a2cfb62936;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d6634b9226c0f6d5249fb393f9c802ea7fa309b74dc1119a1a2efd1c66e1a650023b4752324854a31c1401a1926285ba4dde23923ac25235f9d1d8c1c285ce31bff25b52e6f792206b257c3fbe4d1be8678b7f3e0aac896435be2df938f7b133684950da7a9689c0e0317669554469c8ce4a0300c56c61f79393cba9d1479d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eb2eb32728923e5c0462fe973de603029d5d2ada6282f238440f7ceb96356f3e8af86d0f785b439418063c3c0b85734931d30600d9e3b6e88d9da563bceb354834e421d13d015601f6fa6f66ea97d85dc51ee8caeb7f1faaad4e8b1b6598f62eed0312a4ea4175b1ec1a1d326ba52d3e005e28e31de5bd481ba46a66a9014eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he03996718af41ca5b0eddcb9bce9c9556da2285b64629ff5ce3582499dce9862e656ad9b203ac1462501319bde6bbed378dd101522b1c553c3b26aed6a83b5d495ae2c247d798a503fcdb146020ff5fe113e45385bc3eb8ed8aaac978e9cf78367f3879026525ad18adc49485b6abe98201a0adeee93a23f1d83310876e3d767;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8342099ba07957c45110adfdef0ef9b322e3ade58b5cb2392a2131e7723e938e3ae7adcbd516c0a92b376d947168d049ae808bda0abf3702a32805a9204c02f7f183ba365e89de5ac972d52ecc8d5a6b0bb00b0b35b72eed7861573b311877dbdf029d23b44b15a4fe9ac320b189f2fc25db72aa1951dd305889b11d71a984d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd075e8b8726b6a9f02ad6514111b488791c4593e50817a22cb7474bf338bb855c4a62abff9da03a54e7bd78d00c654bc669440d0b85ec69e462643a0fe1cd2dc8d4224030b2e318c8d59872de047e8f2ad6dfb5c3c32787340d4d3b17267a922a53f1123675cd654f972288412d0dd5076bef365f2d184d61983f0662df49ceb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f4a8d96608043d19409c50ce68ae5d35e2088b221fbdfa43d5ef83ea3b596f9cae8f489d5e82a694cacf63786ebb9883428b7c7d1e0968507f3b27ae4835d5315ffb9d6b920bec76e6a862516d2d84fc9d54bda9f04ac7d4000b119844abc662a8e60660dfbd9a321aa08f84341985d4dfca2df9de158534c7cbf0be4353954;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cee9b0068414c2ce75aa0cca2ee5cba16c683b33b9ece410da3c90116c6fa2ffccbc351e32d65c145b6fdc125e3289ad69a82d8d59845f2c0db6b3cfd3563e3e8bdba77d336823aedc0556f7329aebb7fc60598d2c02050c5eff6f4ae600a3dbd23fd941c2e80ddaf9c8c5d145fc516c981bfb62fd25388121efa67d8f51e02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd38ea9432ddd50697e0ffdde5ecf9c7fa76cc65cdc70dd7181b7e78f60c3810564c57fde18eafad98c2e69e03ec0a5129c41fc6191565534bc1787df85830a319de6c72f4a9494b08d591386fe824150f4cf4a01bf571335563adc4ab073cf9c1a64091c3be7c85e2c0e6184494f1eee581038fbcbceb7b09c11ca95f209ec9d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a0680e5024fbd2256dcd9d843061d6a5853fad683d316470762468d85ec1442c3f797606ddd63ff6ada4c2cdb042ecb5c3d3c1c7bd32a26f27abc8c2c9ab4993d7cf9d8eced2d96503ea6158e78e3b6871a0b40600eec420e5fd4dde8d6754687c546baec84e7b70e776405c8e5aafc8416e74327984e16079c386c74eb8472;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadcb0d534ce70dbc1464967464de6c6776f234e11730a971d6903b41df78d0d0257d6c1a8d42933af219349bf7ee607bfdedcf9193f0f7931932466b7d53e3c71784c5192770668a5350c7b5e1c27a0de052b451555637981f2362b2bf8d08bb6191859850b4a493088a98845684681cc9a69597ce8f659dde643fca5001980a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf96f564d58a73d33d751ebe788eed89669efacca625a72db451bfa089b6924008e7abc1c88071f3c717d4a63bcdcea8021193a78a7e254ed4961f5f07ee902b601c9e734c1c37153a60e16c1721ce37324035be81735b1b74ee14ef1d938c47db649c93c12741f33eb5d38d27189642ba168264a2717b918ef8834291a48e9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546f1fa93a3169477a365b06c9d55824abaf50595c61d644d52c2809a367c07c765a683f97f5ad5851c23d6a25cb47dc3269023e03e1b6326bf796df168d514e9504afca16e300dd311b70818feb0ac6a193bf5b54452e2e1c89d90fe9ee61736710a735ec1c94d1c751f8d2dd139790b5ef72813a1bef205d0b42a987bbede8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c89445b0123532b8153847c3bf1ce3ac66279d58bbbce494c78439f613123cd5927314e3c1c753232069811f0e0f0583d1833cb5f1eb678c427b54c30ca362a14bd2712a9c8a440034545502ab048ef853be6838906cbfac5ed9f7b724eb42004ef16b168e33ab53a80be5afa244d1686cd389fca726874c88761b44b33cdc8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97dc9dc6cc30abd26fa33fc50498568cd1af174dff5527fb5dbfac15d3e14b47893456daee5208252f7eb82c4b771d8afdceac63341d5d53f7920eda3bf2c4cfa6492e58f9a287f2a66be89a9bc922784f32142cf7d58bda0bee14042aed1d21ff9c67a403e5cf5efe42a5c5ec815350896e9dedd93f2b0908bca2acbbe47884;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha38fc2f12d83a83ff1a1c4bf074665bc57e7a13c3a7f2c0b55369f7ee05f5b8ae433852dc8c163f6aeab11adfd351a8d84e41f189dcc4d88b45c9eaabc5be46450fe3496a16214883c6aa17feeb6f2b12c704d6e219a52b6a3e4fd66143368256608b0d3a696367d7e42b1d767ec1c082454152689fc961699f587c99d4574e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6346d11425e46717c02fac1f2b0d3def2ff79034515c81db89749dbefd639972d7826bcd1a7f2420045416308ca3236b32271859916b7edc5817a518a9c07a37e5e4f0aebc7490c487e1575524d8b6be7b6504658556e9d5d607fe43d8f31fb414a2c090e15255af7c78868edee1a475ccd70f86dd2607bcb8ed565d550c3911;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4098add09520a7a58c0840da8f83b9489d22fb8f3cf606f05ea0ae85a6e83bc0eb7c5f46dd99e26e47dab9ac6fa4185f3887b62bad24cb868c97ce7fc060a2c8ffc809a64c1f47bfa07108aad04f1b105a410e9bf514db0ddcf8718f008b78811803be45ca8c20070a54db1bdf48fbe702b26abe5ef5e37a3775e640c31d9a3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e48806548873bee7933d4953ac58f7df81e095afe284e82e88088ef6348c304588f635b16c4dd5241aab02486cd5f459fd37a13801470ba06e1d9215cb1f29ee4e1686fe2d6fe20a7c667a176b7a32176bad1795692e507d87b2e2a0677e70e9befe8785f7c5e0be8e01d3b9bb4e16edb3586f9e4cc505bd69bd635df4384c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbc5425e9994eaaf45c02a3e8cf1a753d84c9664a3fa77352c2c3ba8f8e505ef9367971fbc1a30e3d7c938b3c2b3dd989d833b25a7df7f2feadb89ebbec86333214d04faf31d6f44cd8aa549ce5d86610397eaa93312528962804a455e88de83abed9efc3db2bff9735e61920a5be44ef3b733b9b8eb2e971bb217874d3e9bbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd346d4b8570a9f4734d7cb8fa892ea541c0a41094a413f679cade2af3f7c5ff0ed3bcc3c4cb148fe64135682966df684675a4ba4d0cdfc8a77aa06a535870da723eb9f52155e48f713d4fa479a52da2a9e351fcd655c945b6dcb62eb01307a68dbbe489e05501ca364afd61f719ea26db9680b9cd83b3b95d863a0afcedb883a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ce937fb67842801f5316cb669be769cb2ac3d7603ca04bfc8ec272bd8901ff41c5caf699e861e490a3da365122a8c9f1a0b64805afda95a27c85f9eb5f6555f3e0b0e1905db1563661a89410a7563a3bc6211ee272f14ca2222873a89e090d88bd5f74323a04db074dcd83745c9a431feb9164e2f6e2cf1746ffd1134a05571;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62daeb31abd61c53045408d0924344fa82821d997aa4c1116da01d5f0512aec8189d703b8e486af9806a2013708cabb0843409517fd9bb0a20b579fa17b57ec6a4f10d403bb59f1c406a8c294973be12f9e62cd4298af01c4a46980108f7f190cb4eef7e4bd9b82297be1c71792739a21be44119bc1afb87e4c28b6bc3db2e8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8d5084efee8cee7fc3e4d285b7b643edb472ed0e8277acfb6214090689c7da2244106a6934094d7268175692e9503b223ff56d10087e0aa94b338052717b6793efc8fa4036596816b748d660025c112244bc5d4aa43c1a453033f3c300e99fa9899f220fc443b78791a6bb2fd7353285de7e227c95d0ce3e4914f8ea3c416c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5808ecdd3bf6f74d82b38fbe484eace2e132abd298bd9e8719bf5196885d35bf80f619fcf2c1f1267014ddbdf41588b7c39d0c2c7832827d47b46d3dd68a98e99270ccca9d39b7d56a1734301f76a7d887ebb8714955a4cf5433779de79ed05e54d2f463f8a3d97d06f765a904c3a5f1f29f1e4be1d09b3c88c04d550a9dcba9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8e7b85e372f3b91b943b4b4249c4ab727ddb6a72516f0e713ef1ab0f4cf1e3611505f80cb76daf0992a5685988bfe641fc1580bc9a7d09248a8fe01297ea92c017df9ba206e350af3b199295f9c10a5e0b0abf7c6eaf096742be76c76892da4bd02c173c9f69cd90d56669ad9f7262aa1ea8231b22426d4de05859865dbc75e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61daa5038a90cb39d2b1194429c44ae59e377c99631214a38b98618c401500ca8bd476702c363c110968a25bc57164e800c5985149ea0ba8ebce46d7e97b3f0192135cb77cb6cfd954201b883453ee116c294e92bb6d6bec5d8111a7114344465d4e238a35090d88d1137d23b41f2296da35fea6690076929c71f7026206e6ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1542d0cbb8b706c1c270223e6f8c03ff5d31e58510000f35e7031c6d549701c8045268d5f400f00463b0aee47b2edb0b556c558a15b25a70a82623b9f937990ca0bf9365f2c3509c5f7fd97e2a06d41a5c94386d944f8d18cc9437ee39aef3a930ebe701c3e1e48df3b763eeffafd0eac758250ae9ecf14961516eda2b507a26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5244b2072b5b35bd8564016b34a2946cc4780adc67dd597ceb6c37dd3fe2a775f22bb866cfbad182b30476ce0e87085c629cbf2d0ca331857286ef1c7997c07a2a56d1711f0bb9b73c59cd60f172c77f43f319bb8efbc56b84ca24241bea0de50bdf75b82b45c089d68f5334078e0be6081ef3ba1c9fde33a15ea83dfcc72f79;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fad24ca282781d6aa2968f9f2a275525d6d61576f5d7dd6bb6c4c0e6ce20ee8e9e898e3843d131c4a1aa7e20f42c2aafbaaf8b337cd32d55d44361933001abea3c30b478e783cb33a72d47cde22201c601b067d8a1d03d6958e104b9df720b98af1390eba741101e46deb6658ea271cd2689897017e2eefe893141ca194d480;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38e0ecb69229d1582458ef1144fbf45de3e4faea35b6aa7cf3e469c0ac6114b0c48f58ffa1511acd842769c9a938089c5739e923844810564ac0a43cb5d0797dda278982b6d72752dbaea6a794dbe2eff71867f7e0f49eb55e8a34f7b6e5ac6dd337fe7f836fe671f8703cf61195d5380453ec5fe439c491732906d656458f0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdde5268bd8dbee38850cc4a6e8515926203db84dee07f02c08ab57c730d60c4b2ac2ab7aa5045d8674a2169feda09ef9258764b6d168b1683e7d747a56ef6ff161def5927cc34f4f2788de35b3c4b0c922bf41a51e6b6f041a5b2a3bd48b5149567f56eff9406e79e01878577f7526329c2f5ed604a1b3bb4d23c002e873bbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e8a9dba43b6579fa2fa98060f832b33b85149b01f1fb82afe552909233b00bd228e477ddaec63612eb130548b6ae17450974b87676328c72ec4f2c02eddeb6f27f3ba3b3870dc6694b9fb72f00a20a2b4a3baf1d47ded24179cf8b40492d39f2e390f2d115cc9b3e9e5410d00bf8dfc5006e5097b0e1e3b4af78216e45c2895;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36de94d514e431f3f923ae7ea31af116f3b3b9c35703fd577af3fdbe0306f46377225794319814e8e24b338bbe0de265308c358b6abf5c6d0998a1a00e76d27144b9aa83de5494f82c7a30f761c79e51dc1a7a2a61968d6060cd513cb7b34d268b839c741450c23062d2a769c720ec2753455d78ac52ba979bf999d3e28da2df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc459e50393032fd06cf67af1048967b60cb7fdccd1ce9897161f66b49246286973356e4e579772db82b98ded6f191a58fa89bef046a0fefe276743ac8858d1dcbbad84c8ea5af3b0a25ace3ef31e769ab57e305e4aa754b906d6284fd592935d362693dfbe662f638f9dab2990690e8778c3bb7af83b6b88f5488b69923a5d83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e3df6cfa9211899b8f9f92f60721d0e0821e839bc8d7a6772e07e09979aae4272e1603dbed8e856d9ce5fa773b38cfd08b72a03dfba462dce60bfe0e87986ee5edfc7d3118dabc7c2ac74b6cf72b2a7607ae3c27e4eb8613164006b54e087780c552b5d8a9de9c937793695241661a110bebf691025617be0e95abfcff75508;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h891552860325f33460200b03ee0b5a4f94a1ca81090404b7184a5ff46c7f0a240e623e9f0c029e5bbd068b40907485b9a9394e2d87f45145e88a3dfcfe76ff8cc105efe5754fcb87de46a0c9a35a33f553866ef7d46e740c06bc13b40a0344b8beaf42ad88e1845e28f2d171b00ef9cfaea55f5a8ac414b90460084e4674e830;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95a9553c99c4711316872d60436ad25241839ad56fc38301af8353aab14788549d3d4374ade2662fecf04ecf81b4db3467ceb4dfd28cd25fed3781d76124d5e5c8461fbc43d1f444b0cd26fea57698dbb56361df618ce45e4e7210929d649c9cc1c1395a842c52229a20013858113566c856dec120ddac0c9405fd4ff599c0ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5760cae5df442b5b512285a4694d0fd80a17a28a78605140baa69b171366aa128d9969d5b90ca693bb405b4e365719f2abb250670fe3a2bea28d51ea9f4298ade031f9459e52fff7f5562772f2da53dd109614ae44a714878aa5434a74093711957cc78260a23b97bb711642972feb28450bfcd1a5826b46ced72cf596955a07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a04502a25c6ccd8ac645c17a09b09ddf3fc09309b22aa0c38c9696540bb2403b2a819d18b9f77eea35ddf7f7234b54f76c272d81f18c4f0186843e76000b1f3e1989b544d989e91e359eab979141a388ea2a1669c9c510770baa4118ced1e483053e9ae01a954e93b1416b7cb961140f9dbd9e106d36d69fe17047272088e2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7d132bda9a8c42efa65e57933df9a55d2a980c756b8fe4b63b9fe6dd239e8c8d5ad92122fe60d40850d5797538ae4c1e9f148f392d9fcbc9dd45d0f4325e39b66ffb5bb8d44cdf1ea6616f88a024cda033206241ea342c1401ac42691aa1d0352007b113bada191aae0f3d8e57d8c583e7d8df13e3b3bac9e68a169de4aa3cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6ca3c399698cf1f601a8fd6cd3525d512c4e0a294041dc86f7799d243e92f2f162867b6e8207ee316dd83b79aefab5e7d1366120b4dc63fcf34885d34c206fdd0cb9a17a136efc7af919554d9c692b9177903fe0544de73a796cbc6a0b4e4380b715f0c466fd574f40e3eef4b992bd3a23c5f34f6e432327b43a6c89957b6f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbe7058e88773932d2e07c2f5f31925f46e3cbd0d44efd17883ab74bba1bbf5a39bf8c96a1d72849f6281da1ed47b70046bb43045f0cab56f5f6f245026ec003d2b352b2c40e87d951caccb0f91bbf23668ba937eabfef2b66760377c1a78f43644debeb0dbcb2bd0a1546b49a8755a302aa9dfe718e73d2b8cea6ac0df366ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h703f575dcd51e731768451ddb4cba6e11f520e128ae90bdd477ec9288429e3e1c05029a173604fee53ac6e21f5474ae39117a831e2bb5d332c0f30bfb83b88f3168e692fcabc967e0cf7acc8ddade40611f7b34d49529e345815740a3425711a6f3581c34e08d0086e098614406c41b5f8b0d13eb7c4f887a45b887326ca2362;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8e92b7a6aff0cf21b747bc7e6ac81188046625519d20bc1c03a5f777c4db9543a4b4d320106538d52714bd07ff87f3f4deaa66a3158a61183227b39ac9c9b675e2b9c638b46d2bdee1b610ed2018d76181cd977de8d7a4d91a9299b2a4737f74220fac3a1ff3f7d2eadd57a2d3e29d79ea64d63f38e27b41fdc90aa350a2934;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1c6a95574d3b26cf97c4e940ebc14950a96bc7f673f738efe089a5fbf4199d67bae2325908462bc91574d60a13360f0b2248e5cd3d2255625885e2cca24ee688a88fff8d30646d16086a3a032e20b483ee878bc1749d9dced22930c0f5b28eb3d3aea1808d8ff95264a0f1ac567bbf77214da78e809d37c163f80cc9b84a81e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd77dec2cc02d69747fbd8c570d31e7c801bd48b0a88ce818edcbddfe11d20f8aac058fa19f0357d675da60e409383942a6dd6c9f3c33e95b5b067c3b74c6b8ac0da8073b8cfb538abe13e567c2c21bcef213ab865ca1a7fa3835265ac9a14a2f5d30ea039837352e2831e36a7ed856cfb73db5c73af8b05a60aa9ad9f87208e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2bd9285f39902cc48d63a20067f22bc372eeb4bc806c64a35ddbf85525f4fc00802eaa75d25fc9a98ba0c31b1cf9cf6e9a749c14add87d36c34a962806c460b28aece32b2c438b1ad6464e13dea8f02c80835386431c0ba727fcad4179cffc21700a392110d95bbe4ec524168dc56026fd9c8cf48fab48e313c383acd8c4fe1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa9993ddf19f384148f72759e8d8616d7709807d8b19fbd8784cff2ab07e256e65bb7fad5fed7660db4b42207aada7bc13023e81fe74f9823c63db156337a277eb69175519e2ac69f4897ac746d805a2e87f8e6bf6a3d610c0adeac7739829db262857bbb79d8055894d4c03c2ec54daa799a5659c171e15df3142ab220b41b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he13c8ce522fbf408d773030459c4a6c7740dcd0952ee0ef1c5075734d772fba9e31352275a82ade1b2f574beb04e52b36c57da6b1228280608fb2e33c9d385a5f39e8f018a3a0cf07c2eff53089d990eda729bc01bdb538fd124f010b224f8098f368713f49c0d3a97212e92a02520bd90368984bd2ff8f8cfd8d0903987fa64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8323608c642f1c2682fa0e9da43cded929a083f253be9d4988c8d7e396dc9f634f6d4869405440f5b7ba93a4bd5b9b1253dcda2caa16776674dc7dcb66dc8f59914c50d3fb88dbed6698a12eca86a1fe17a8b7bef15ff8af7aa0a4718e382bfbb95ab9f2a06faf10004a63861897d827b5722c369b4ab69b98f448abad93f487;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h932c795f5a6a37e1982b584cf5e65313426123bac96568c20d57d332ef88a39a729f039a1490ba2c1423fd83c50246cfe76b843215eba001d8e22f3549caa195a3c36c3a37f36abb78baf7bd20a7effabaaf029394925e1279a3812543db5f42e2cdd9b6e9e5d965316cf4ffca2115163e8264bda46044aa458a8d0c917340ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15c17c129278867705922328d63bded159c5e62e4911834ffb7b53b27ea64ae0812fdf03e0b78d5520f82186d70363bbc225ab2f8c276ddc2920af9d9be38a244955331ba2e434ebbd67f8555e5693e349acd2aab2f21e2f44938c339012505eded3150f3d20da5840548677c9af242c76a0a2634e1d8944d01f5a90a686a79f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had4a317a8f4a6aad5de82bbfa75589167f1a4f17a98ce7cbed742c0e401026bb5bce33cd3a7a71d69334ac13cf7d950d6540ae8fa07bcb08fe268a1666c44030f275a97f5936b48253be137e9860d585c11a352f407e84c577967415e636ce1f37b27dbab1922796557231b9058297bcad144ae77f89d6df3db05f27d6bec41a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8b6baa151a4ff51df27b379349556cfde55ab714dc9ac39e61e6da9f1bb4e689a8d4a52baf0ec80de5b89bbbb8376d722e09adad0e9e97534914dc8ea007badf51a385cdb5eda9ee064fc1431bad2a03844326c84057071553f2083d4d90712190752e4737a075133c5b9d9afd0e4b24820c0493bcf97b0e79574102823340f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7117146192f701a34f20a10115831654b6448df16a5a77e0e728036d2f41dcad6f46d72a870f5e7c756e61c94d6b2873eb37ff65ee78ebfce90c7bcd13cca9ead74d29f58f2d316b3774ff7de5d2709666eb23507ec5bb40ce422639562bd73b71daeb55b4d8262f4063227047e633c48a5d40752d3c1b9a1f9f39e51d60a75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5568a33fdea495d17812f170a1b49a5e5d1975806d939f2beb8e7762734172c328ec75a7becb75d3d736d749b8edffab00ef65a8a2804d210802d38294980471a265a74eb6adffd71efcc5cc5a6e4f87fb4dc0cf961ae66131279795337a05faf5373d1f6d9925828398ad96785d8c694edd4d080c68d9d4c62435fcf2f80fa3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h393fbc2c52cdb489042d6f64bca83ed79d6ca5d979e15cde8891ca2d40c70743d21bc2d89334abd8569e50a996f55aa8488af72776a4403c344fd2331636c8385c4cdcc8b85fcbe77ea929f8837dd1befccb5232ee95c5ab5d9c5254a89d34926768fce390d142267c2d54e18e55cbfd80b490b95d5699080c208a54c26e5401;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f8209c3acd0a16e4cf0398bdf120733c7f97c733e0aba12114a53880728623b4ebc6a3ff9b8bdf25af998eefcb471da8c61e598632ba9fc09a956864333bd39a42a6658c1e70822c9205ea15cd9b2c86f49c713fca0d3b6b1d7d43e50b9536f4450ce129049d90c4e52d5441cfbc13aa658b309b47a5513a6d101abb490d604;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cae414cbf05f512e315f332ccfe6bb60fb8c7a87b2a4f826009195f57b40d7e67672160db571025d16c177c2e54ef243cd5cdfd18f2444897664d9f49f4378bda33c8c58f4f8b837bf5ab929dbbff0092228d8af8915dc719847a0462584a7045e05bb5cfe090025d74123caba5697bfc6e57bdf7e68b3dbec1c96f17f59cf5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0bee57d9ec633bd4e9ff28f756180379b6f09f191c440f0606684cf113177e5e633b31996eef7dbf006c78d55567eef3d9149a9e582e568e4042ae24f5ac8d85189dabaee466bcc36fb08054192100e4f214db16865c42c61d5f6db7ca3a2b468b8cea3987e37b647b994792913fba3d0eb08ff78a9489c24051319e65942c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf78f01fb4d77b38a09520fdb9eb72ca5ec923cb084495068f5b7fa5bec015958ee076907c3779d313c1079d5199043b49b8f5a4e585d5ab490707962e209fbe88b842c43d52ba87cacfb867a163e8ce257131a452bb350ad4ab924e7ce293a7739034069d5dc86e466b8322cf111fd571ca1a665d9217f71c5fdd444acc5ae58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54b512aeb72f693b04ac502bceb6ed8187ed61a0c03283b686486d8a6c4f82e82a9a31abd3cd8040c9721ffe113877008547282344aeff6325e425357413ef7ca6eb0d0cc27b88f9bd3b0c08d4e7a4bd415b916d2ef88e2bb304a0abf0791113797c96f1e4f6e633a9ea1207df821cb144bff6a7a1694d498dd4d0539a1e3ba9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h686cc5f79fabefc68c3704c6e523d50586554f2706d33fd24536129f1af6c8412554604973980ba72b077a07674ede7db38043fa3c1e4e9c97d1c9216af84537d1145addc405b20021d8600994e66b45d668ebf0b5b952a8e0007124dbb4a86c45c111cd55873940304b72f546b8f2e41f0619bcc4928492a024f092df5a63d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c42618b49fc6259e051e20c1f4bfb262d6e287a547e2319e785c907ffdeb20b5216f2f813232fac41df32bd37b0adfc968062687d8d80c41e6d07a3a4524c7e0f5245e4a27a20c4bc980b5ff16a8533817a981adbd50d884be6e4d049ad94e2638047d58587b63a3d354d8768aa0d978cd2caeb56befa52c6297336513661fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb94a0cff172124d0e40c85b602de309c48cf905e2fc6b32c8170df11a75dd9277e57974ad8e1fff95e092778032253348f943bd6bc50f927907d44ac27e7d9cc3bf937a5b058fe8bd3751f243ed258b1951606b213721edd88df15b99e8df046cc6fc7fe347cc40c3d1154d53e40c652fac97d33982940b35175c408f8930982;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc36cd1d221a9094f77ba14ddb81b094053e977ae3c68007bc786642c03a653661e57c5e4450b97a126ef492312a193a06e6a0a943300f6db9ca48a7cfce24adaf954ba9403c88431f034233f74ea06eb1b7763181bfab4a70a9baea179428799c489f5dbe6aca9e648bceda1d3169280b2612ce9afb2d5a7062c1a88596e1494;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfce6a4b1acba391a70536afc00c1874a6c307efd58591fda338da2102b8f745f959f30968595b471afaad43be43ee674fb548a5f39b5fae791ff8cd67e4ae01446533ba63dd693bd79baef2a20954a7f5d9ea1fac1107c1d392970f51e4fff99b3ca57c7cd2c8eed92001004584f768c88233e0f8501583c3d9ff8eb815e0af0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h900350ad07a8c64fce5443c50ebc39911097673c592ddc7564272ff7608a5d6cc848e15623f7e9e048f8ae9079ea5226178b316da057992c46d8d7036abac3cd3770ce26b61ad5ea233a446745cc0dca654a2e10452ba62b7c68f7656053c188324fef8af79092b93f3c26defab6237fa1fbd2f91cca4d513be0ff7995a8503f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd12f5d27204007443144a6f84c5653a7cde2a1a4039240510249926476616403ce2b30495f29d5ac4436e88ddcfb886217ec8eabf6cf28c0590361d4be18bc2b615527cfbee268dcdc5ef1d032170385a508121b52dd867e614b47c1a4c0256056ef1a630dba8092c4e27461da28849ec2adb268416430843686f4f1bddac47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h444222096d827e990af696cab7bfbc045b30e83973150e8ab9f2d999b5fae3f2cf3046203775feea9606c10f44ca240cbbcbc5c5a193f2b44b7fc6eb6edc65d9af3263f02e1bdf1f1d55543fd7ad5b183de9e118e50dbf1e00edaf9b7fb30a02dce90f389079ec20f64740c436dc6b80136b97c4703c6d4f764ef83b40ebfb74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20a8282b094ac0356d70e28dde3ce4a33568624aa0b46bb4db4458a2b9a5aca8f9f7bc0a4357f29804c4f0af8e27308d18ef4b02f6cb59219ff80b0768842aa8296c7d91a0c549a02095e6b390c38545970fa991326cedf72587035869a4f74c33284477f50f22d51cbf603c3284f202f6996890ab7f2c762fad68072e1c5c53;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h994105613e43fcde9885b4d6e2dcc88fef7c57aa2cb360268926034899061e6dbc7ebc98dad4fbde294770a8a09f52d1281aee78498c2da84d3605dc82d15aa26412fcfbad99639b96f2d72c7c2c0b2025b9a3b754c543cd57f4afa6dfc0a976627a682b648e30012ba561b88531932932062b0fe48d21af7c5773bfce1445a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67a5be79ddc886b2b0337d350391c8feeaed3b297e68f716b8ac97e3e01932571225c64e238a2c6de10a31da1396fc680e0b880f49adb90aa1b69fd1f05df09128a2cfdd3df21243febaa206022558f86c4b04a817d74d12ea7722be1fad404e9ddd66cb41791dad43e2ac7259abe92939e9baaacfb307988ccc8892cae6bd48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h790eecf258df3ee5436c98b58432cd7c72d2f2dadedf10750c1317a0f963feb5d3a2a0ebbed70d91112afee41fa4fbbd4c9a510ecbbe4b2429a00125f03cc74ea986eec6d1c04c62e4e346795687aaed312fd490dc3fc6b51e6e3cb701c45e985adff055f07992ebbf6a6fc63f9723d16d435d9ee449c530ae847c3199cc553e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0d5eb0ce0a9bb7356bfd61e17ecf0267aa654b292e736385a6f506f0facb1e91509dff73bde12c1aec47afc5922e06dd77f4f59665dec37bedf61dfae1f532466e1e5b246796bd36806287daec05bc7860e0478d4756db7c79a35d3910f14714cf016813f7f176aefa6119575d0d2873a0766bf5eed3f76d53f2dd16c277bd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ff1c132406bd6f732cf17ff37264a5858889f7c6764a5a8292bbbaa36bfdbd1c22662fd67d74dd5cec4c70f0ad1a697bc8969b05752495a714b415d31031c353dc421fa41574c0ee1d6e5393ae92adeaebc2a5dfddbdcb2fa2b0bed11f7ea54fe6677f1d1f14d48ed41f47f1506ec59785d2fdd1fa28df2ba4b44da94a65866;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h354369994de2a852dbcfc5645d20e5be08cc559e67bbed54631f493b1e59dff62ee267926e929ed6238fa2a81d65cb22109dc2fbdd8770218fe62f9661ce24dbe1750b9011c60d0a6c8ab0f8e75b9134d918b2e05e573853539bbeada36312bba20fc3e0f80355471d9f3d5a2691bd2cf686292e3014da49b80cdf1fb968d2f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9207465771599d7cfec110d3da09e22bbe2d12976d82d7e515507bcb64388f1855fc85177f608a6c32ea1119078e876c106d7685a50cb9fa50acc4fdd7aea2a7f9ff75d5e352ba12777a025f5ad78ffb034ddd5bed082a6768d622d014e10b04bf72988939cfa8fdf83ac3db2fb756cd5efc5c2f8e4bf342242c4dca818878de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13e34495569817ec6aa1de50dccbda44d7b8878668d076a620cbb74d84050f971ad5c8d911afe24a21b278181fcf8d1b195b98db63aad734ddee6aa6762db3584a96dd9813e2e06a7427e6a53a7392b018cc7743edb3257641d0f387b37e66f5f6dc6a541f154339dca81550fd357c3fd0501e8d78f62e969af8f2e92866da7f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d1af68319a8bd4be13cba5c6f7c35e64b68b02ff3d4d1104c31a74636fb68562abef7c75ba369c74c98a22939452f5c6d2757430b018aad5791c227381d7a749fea106ebb1a020e2042742b1e2a599e1b780683d6e8a1fbf0632a1879f710fa1d80cd2a54596e9bd5615bf42db01d607fc686cdf53ccc654a9d2678a5fbf856;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fae1a7b085cd5ff0bf2def8a5dd0c6c8782021e2590468cfafa0804b6c0d62c710c8d16bfb3def4315daffcaedecde6b4a60fb6a86af798aeb33d63eca751912f6084c817b5a0f3b4991f9767308d79e4f7cde6bdea580255c6e53e40230bc68620da387fd1ca39b02266ba2ffd5f329fe8eb44b468b82c169c5521679ef335;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ba285b4c2f3b0101ad10874a4e2bd5487d25bb9981a534bce951d7a2ac9d9c96decbe7dd1681096d63a4b5d55b31a4d285a684d9aa4e8a83280f3e8833258a47687be9428ae143ab9ce0f470f88562aa1ca10f8148cdb89fca27e613da2348146bfbcd8069f3ec8d3b76701c78600cca7cc7c4d10bc182b0679f701731d85ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb39519fe51766f901bb75479a18bca5e2bba7a07316e08169cee1abd9cc438fb10bcf6d3d96e3ac42c4cba79ba770a0d09d790587f77f75b5ff91e0572613bd939d39c68a3f285a639bc7389f9908216e2b7f1f8136cefc60875ae8580e78d1ff08f62f9d47a00a2cc58f7046c5a407a86d7d1d19d529a35fe62bc457817dfb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78e8304c19bdfbc8e35b3fd16a8985d3afbd58462dc535c2c77058e5c0010c71ea754b87bd53b777b784e7cc3a232e9799b884485d3a207f827e47f683ccfb883b6d81d437ec4a09aba55a9a498eb2ee372acb0d7f9a3525f65ee285b6ae327909ef503dfafd2c4df1d86866b5a6f15e3f59ce2940b87724c11f487474ea8d21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he48be06597178379fb6e1e26df2a2337db6729cef18e1bde14578aa480575e73b8fadadc3ead272562e00be050b1944a1bfd99ba07dab7604df2b11417f52706080dce72e129b84cc50912bb2d14387346f0c83f9f5e1dbaa437fc8813d63ae3480268a5c8016f242f51e59d760680fd7dda20883814a391f334bf65e72ef663;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93b5e5900826a95fc2ab8e9225b665214e2a09c3f71117d83d6e27c53720289ad921c7f1fb8921c705e18cbb047b589da4bd758807eba068449a9ee7faddd69d27486de43d45e8b50d34cb345f121c50008f7691ab8118bcccf7f64a6dee6f5303fd498efd7290f9d433235381d6799303a702f5e27475fc4c72671aaf1ed022;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb710de0adaa8ebbdc97aed22f3239f62bc95f62cf5998276336ab0bf66a2435fcd109fc5b43a5cb942734898b2f3145199971707af56163a914d1c0847d915822c896fcfd6881e6c3683caeb8d185be526d22ab5cacde8131a81174555ba65721df849d5582a746365ef157f55acf351558eebf7fe4e3f7aa1d65ed532f7e2f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f93cfed6ad34fc06e1e1c0b32def54b884c681927de62adedafc506104456b0371b2c5d4b5fa1bf128c5c57aac8cd8bbf18d8733943ff9a8fa3c10914d87bb0140c6f2accc5f94e5ac7149c77b57ee27360e70d7527faec6321f227daff3f361b922f43d7cba05a97661f86fd4a7aa0842c82e44d0f53276c605dc544d37030;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha878a2a3cb6b1937484b4d0d25e5faf657114456a5b176cdee2a6f432ed63f9fa3b5343e65601ff1da2195d90071bb61709cf800c38b9d8e6560f6db1eda5e0d72bad438d07f108a5d8cb80a684758f5c8b5be9e2bc6b99d0f574f17606ecc77e9aab539991c4b0c01a53b6cbc25041b22807fd039386b12671ae55c24a7240e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heddc0a4def3ce84bcd054b5ac2700badbf0cfdafbd4ec794020f6f7f611c55f821bb48143a689e38d2124244cc7fa31cd1626b24a5208ea873d1a8fe1648ccb9404152bea4e5e9a090d5a74f300c5bc749c1085719bf0bc596fb25616b059d2176730bf3fd819fa0caaf7d07adaaddf5b1d5c232ca3dac60afe36ce30075ec21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7ec73c734ce769e4abca3d5237d59071a06e8ad6276320039b9f68313576c8548f25d9be26cb5b7b736c1b14b5e27a9f82d616794b31022159355b8156088fe104555be2edf3fc5021307d1dace75219991d54a3f587566e6e7d1c6cadacee470d5bf5b25e8b3d91cff010d608e1ab28d895d4d4990d6aa8ef2c34d7e30642c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6487925622dc04d788e8ca01966e9708f6368f5030b172e584e492a93a79ef97d10730046ea273254cc5eb94fd45c4d944364b84b49e66a42da9eb2304f6ada79ebd9beb4b85a1d3b9edd3a490a5395aece6689e25d82f1dc2156e69d3db6ea887e5a85de33411b36c5ea27356b75426c4bb254d8d590076cd74e3c13069e507;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b4e804445629a636f91d3f61e68244a91df5b4db6cb24c50cb2898d52316642796f1d26b8eecfac41b06f536e76134829f36dbe26dc0d24e683e76f7e339c864b714cc1dba057c2cc030835edaec7e432c21ead471f601c77636c9cabfd8b2834d6f1045e8eb53c72b5dbed2f7ebb6b78cc9381bce88b0179f7701ad4267dea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71d609258900c13f2c6355ec255277fd8241cc96d7f415fe175743b1cf0db21be5d1d833068bce415a67729534ac0cbfb6861bdf05c1a7657a78b0608743e0b7e51e132c920c8deb50f534688520bd2ecd18c83d0d3c437c930c26d760ce3ab0c644e461a9d1f64cf412836f0fc5b586d0d1f0dc54fb4c5e213f75fc2c8e0ef6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e1f123a02ab0e33bf67d5db8f66ef02375297e485f3d820f9886bf39f3a981c6e89ae84f50e2a61ef99fa20ade4cb1b42e86cdb0594d02db2311a3b3e8fe544a63e32816fe4161fa7f546e007014c5a3f5cd344c932c04ebb37cf1f70812ebe7dbd86404e2b476ae90e1205819b79922387b1e8cab315eca98fcf6bf9c79dbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdea2517005e15fb4deba3557f0b9bc7758310be5d69dd61db41ed0e871bc455b041ca547730cb08e143a4f08aeececec297ed778d3e4eb2d21a50c3fab6178cd1575011e5f28eca1c9a33eb37bc3c967f5ed33e925b40716c301b3639b5971953d8bc35f29f81e8abf998ba1b2131bb786d41123787e3eea523ea2ac4bd51ffc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1832f6d950ad412350c36e2f0f6374ea9d186cff9f59a7a6a79bd34aa2be6763fcb7ccd3ddb670dbbc2b17901408923e7c729f28ce0ea70fa712fbf9b3a4a10ac0f097cf5094578103eca3907945d7285c04e22a829f25ead43d48161acf1be45d3b74934ee4727b420ab0749eb5bb74ae58f832198478c392c164f29bd4e9dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fedeba9b6a5b37dd8e917245628faef69c1bf64e51426f364fa5c94f43306dbce25aacf48761312171171cfe44e7054980ac0cd9a7e8b41fb77391978ccfec8af8d439cbe1d69d5bf616e148378d24a5942bce0219028346c9d7e0ba1f4fc88dbf9e98bc24a815c5f5c7fe0db1786a529fd2d94c54114fab3734a4bdfeaf885;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42bc17b50bf4d315a8e826295ff993884c993ce0c4ffa345e6cf244ce685d4b66d4a1fbbdfe0e69b4eb3d46744888fcab73fc66f7c036d10658123c7e67c8b7fb2ce7f0e6c159e2eee4708c694f21734adef6ef3402da923425f33b810414bf5fb662f9b3e61d41ce6d7f9bedb48c7ee20a8f77e963c771e11585cd378d82d45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59466b0d62fc9fb0d6d10183de9fdf5aa706b0b08e3a16b75ce1e53ce0ace85057df777dc6a95ce7738fc45c47e6d88347d8e649af4ef8ff598f7cb0d35bb78584d85b5dc40d915a1ba2d966b231dde0a4e6ad5d165c5958975e00e151e52d6acb59da0e1ea790427442a489b92e9d23ce7498fc105115d0aab4202b896f590e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h100c4b714628b68071517001831ae0a4ec074a80fcadb7a82b07e8136fd2c8579caf1ca49325c11ac133001e0fd8f26c37b642ae02da27d1a91dccf4a3c7570cba54dc1f90194e333b05d330a67d7d6033b923caaa6d587a8d7dc840b6f56b6f1728817bffbad4f6ac3a16f1aac2595e7fdbcedc9eab734142fe7e9f43bdf2b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbebbda43687366eabf0cd99df4ac24a7159447fffc1bf146c64b793ac4c4cb6c257d9afc1e155a30b9c7a854227bb9ad5a8ca07090be302ed68ba435f711616833c3e4dd85c2b81041413eccffe7480de6f458f70bbcf65d0c8ded1657c19b2a45736ffa624222c80b4d37742ce7ce90487a6cf2c0026b85fd87a73d4b46548;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0b9de38348c911c7fe73c295435e3218e7e57cec2130347d981cc8be748c034ce31aef05d9b6e0a925b9debd99100c14190b6c5fdf43ad3594adcd951e098e36d0de1fd6a947e2239659afc4ae0e6c808bdd03e03996023c42ef40a17145a8459fbdc5fa970f9ee0b3a8926f4055eb5cacd8d8dfe9510da6820f265fdb0145d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5734398111f7074222aed220caf48dd78b09100180ce1a3b59820ae59782116a3941c3503ae38187e6b8506ba17e5765c60282de0ada1e1f77ec2f7828b66b8043a346c1f55c0a83c245459200963b58afb04b6849ef1a3cc669fe6374d12107e4d46553592c1495608b03c88f513f7b6decdced57c984980574a454914e1a30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44729428c118c86325e433d6b5dd34c5d641a948672c3437f6c90461b0f1cda22da0d7b3deda89fecd8bb6c43263bc216f68e3cd44dd2016542c809ff914b187d32e1c0ad49694f5a28439e8bc8d1cc6a9e626c3ba95d39ba3d1eb799161bc9e651b70800556545065e006bcde6d281c5134821e8de3ac73e2b54b064562953e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf59e6d01b28913df0c007cae755586abc1b1a93ac06eff70dfdd679a84504acba8181f94a96572c354be0e001d740373819e06ab83abd4db998e93d9e525763d0550b6fe22d3b49a2d28c0af52aa5cfff5bc7cc34464f49f6f9101e5e139262edd44df6bce716d58dced406b80cfea8f58e4154d0c6d201bac9d40edb1fe1c22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26d89dcec4811e768b370f03d0f9238f47239aa917d9d2d7f409bd71d0314d4c4226bf00001d44ca1f0617ff31263994a99a333bd4ebc5bc6ef20c8950ca9b62dcf37cc7461bd676f37ba1d90bf277fc01bb8f46687e19dca65a25104461588cce69840c1f97edfed3288375a32e99ea0d95190cfc444809ba49758628e6252;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9d1d46c31a7d3683241091af2afd911fa829c324ebee140a26fe450c657ce361a561a32e68fc3f2cf22a2fc538eb7061fb27fa5ede663e8e607d9e9d4a95dd13b347667eb73d07076c8157db76189909d290af800afdab36509379ee43cf0074373681fd3871cf128858c0f40cfba4afb83cb89369c231834665224fc878b5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4b9b88991a300595357bb67cd6ddc4889b6b4975e64d1dfb662dfc67e842f92738670e53239f5e43f2d4cc130d216db4005904413492ca4cfd0214621fbbbf2d93ea45cf4103f7ebd52082b583e8f0bb2b8759ac148304124387fa1eb1ef63d4fc1a248598823690c36ae3c25f3e3067f94cd1bf478ccbfd0080a5d9706db2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2569219319b47cbf3ca91b98b485d4ee2a70b23b6b05ca5e47157b5fe738aa474020567dd188ef4b38ddc065e86234ee73cc0e6114ebb0314baf14641169db2d814df3616b317fe292e5c72841a12569294ebf1336331a5a09a6725fcf066cdbdfb3130f704be006c43a5a50b53e9ba5b2aac060450d768532447378761922a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5e9e4154b2cebecce36824c92db0dbd780e50fc02bc7f60688baa9ff7c4155ecd9471d04b0a61eb55bf04900c35f968a205456e88a7e42690df718acdf2ea193f263da5801725d2be5da8c4ccd144ebb89d3ab607be35327ca210c96caf2355756e93ffed2a53743078c6034f971b10e83cff64cd95bb2c5b4c20c1d1b8999d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3993c7a4f58fad23f17f1882e74bd93079ab3e0b0e3657c634962d7d0c609b0c5bca2fc456e8a66fa2d0eb247c74551e7deaea5832b72f809ef5ff4152a66a20a52a5371881686598a76b9d7da117760cc9ddb27eb93935d4c42f8c0a2819dd553674d4b46d2911eccf0c41e6a05a47af167340559d1af5bc9e8643f228ca191;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19565cadfc21a42e41df563a8df004eca3ab02e4426f336a208c091e7304ea95a7e4eba9d6cce257519ef9b452e750fb2541b1817e1e74211043bfa06940201178025c8c41bbb36c243e006293a465571e1ec2ebb8739b0dc42380436b33d6509eb8ad3546c9319d6433321aca584316b44e04ea4eb1111f206584cc88fe46c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8716118941517e6c3f2dd2baeb6ae7058fa4bf77f701a3bbeed08048501b1e4ad54d25cd8fd5209c570d724a5b81d95a89470b1222fd8a1b8fd242d832a5a79c28b8d0a2dacf799ad6baf75c7b1e4a5e780927831adf11c3e3945b9715c7233de7c5c09bd9f37e4e464c6ca91380ed59dc83b29e92201bdc6ea4949ebcc6d9a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h538876d4b9775539827ef4b4e735224d787ba4f80f8b605ecb702c9c24a4ee2aaa49c3281af42f5042e2d9ae72b020fe4cf5ed55bc93c76915de3adda787965e2b3b1eaae6de2c1c4c2f314893a90bf894a9d9d9dff7ecd1cccfc196089b69587373c0df0d1158be349810a18f0eb0a61af50062afe54e36b0146a76118f9024;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70c97ab31b9bbd4d1e4fa504b01efae611e5ea6f88eaa591078518bdd1e78c5ed4eaa5aea035db656854b5c22967cd4f76f80b8ddae7df67f6afbd88b659e9aceb0a0f9f5d28f9ae1f139a629957e86aacef19b5ccbd80e1ba1bc2f53f771d6c1f58977c83d111ca5a9459ebba5ae9a25ca3d6c574a864f4ed6ae339f6ba4e63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae9d51ed02862c202b25c27da442f717f17164ecbc686e4492b18490eb4e08cbc97319daa10f48f3cf1799f7b819b296fce363130b6e3a5aaed08323f1149771f155022078a700c8fc80dbe7eaf296b61e9090eaf9be6b7f92ce38f8b71212ce9f8b69f7cbc7db0b4bae663059f7731a358c8d279631cedab345e93e4f301995;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91f5366fb28c7dcbd4def24ac11d819737e299a397912de1d5ad343957a01a3a7eddee13721206a9eda0ba660812f5f5c42505643f7ad4d7794db58c9517c1e2a2b10fe755e19edc33642c2c2c9d3ce3a4b6691570e589587178dfec06e2570ca4724fe1de0b9e8d5c6e778c5f0d68aef6c28b1b0521fb8702a4ed84fbf5b8b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd74dc5db01aeead19729206bcf1bf10f8d788129e0a1767eadeca2ba2e860a8acd7ea5c0f9ca9cdcd775b2a550e4f0ddb504072512ab779a6e7486cffe93087fdfae8a7d4f5c66fab4348ac45da0288159a0f7ca14e230fda788ebc0d1d59e78d998bde1dbb4e4848e46ee1bfcd52f37bc38109619fc88fc0c74887bc5da15f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f588a6c25171be6d3b79850ff4f9a7379fda30ab5fc0adbaa08e8114a8d63551ebf025ac185bbeca537e59f5e8f7185f7e2458e95373edbd1111fd2d7e9e987c7601df3e3617ad2af165fc3c5c3e316094bc6cbbca48a579980d3f4e8e430f628289cf0a8f9a3ca77249b01b60f12f67aeb5573fb2ef6e2a4eb074a5b075d74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc3da4479fb0f8610e8fc4aac1e4ad3c78c9308d0066aee14ed4b9827d3ee8a2588a17c2925018512e4dc7d1e1669de9331db04940a767dc7a666471bb562db13e1623c8f4cac362f4e28fcc439414647010296fe2ce017c7d41359f30d5f96c278db565d9c78a91017766d7b6706bdb5feb3c4b550cc8ab3c18d54ffba9b5ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ec3b3308980df4aed1dd131ab9c6193bae4cbc492bfa45929e4204d98e08e6a5a517d48032251330a23178b1ab33b397c28365635b97fa510c7810e168db29266db43df001257db2d64ee832a9d41c19da899c00d340b56c8d7d659935b20198eb14d31084d55c552a2bf2ca7c730368f4111010948c1a8edf636d781453726;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he232c6cbdf32d30c20ae6d348c51019dba8dc1ef1c3551429b726ff83f825870891a4872bdb5fd14f97992ef3093c185bc490c14c12f7a771f340e29846d03bbe8ad35dad7149c83c3d726a7443dfab83feec0c9ee4dd2dff3b592ce91296c4db1983134dd0fb7765dbebe94aa9ed2df6afff69e03eec91dbdd7568504929f93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8abb657cf6a0911c657f4b2b4d45eb3a2cc9ba135d37e15c5468fb723ee747d9b884a2eee30316f3d4b2e89f1b28b1344f4a5b33efdcfdcc27b1e435980e9fc514a29a6a9fddf9070e9b8a2c45728a779c7c9806cc71e64ab0462cbf5bcec2d538d6fd5c32e40d511ae1d67720e93f836ce4964b8017788ce29c2425a0aef2e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bb5f54eb79ea5a056ae3a5ddafaa48877384351bddf0209ef1628840284688ef63e3027355422d03a2b39531ba307fa5e13c3441f1586b09a44c751b378114f39622997b8aea080164d19088aae52d1889203ed08c945d6534b3d5167c4c94e7971b044d62a4949fab638a1c30c60c387416e31d044fba4e88952e43b863df4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h984a9c955bbdd62b0b0b1a8fd94684773bf6abcedd77f43c3beacec659cd14ba44b8a8215bbdd496e2cdfc6386c0c3bb289cbcc4fe97c4d322c3c43b6e6d4583a5c27a28b0c1aedf3e5721f4ad98db1fa7ec150c49f29eb054ca60fabedae840e5a8f134d23e96c4a043464a6184399fbf8bd0f9dfec5a700e1574a34b890e49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbd5b67cfe1fc7cfda7ec08e2d6587166e648771592c1326a1cff7a563d5c53bc65fce59925c282bafd760768f98764829eadd0cbcc94b6ba8a61f1376841b3b0607259b986e5d6c0e1a0a0c0772e2da334843b3c7ba40881b2fbe2128e69567bc700458f1141cde861871e34bf4a7edabcd8af72d0139ca49c961bbe3c972a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h782a6c1bc8b96b506c58152631ed1e4c521871c269e3bdc67af8b57bfa46d334180f036236f4843577b2246a2c643c3c208438fbed15789d5281b02c5cbec16982277d828e704c21e67f6091330af81f782099fc73d6e22f054f641bd55f30ad1a566e323d7e17e5aa58cf2a1bc90fcaf97b55af55f76387a4a3e25e38558fc9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51503e5ef244578423dc261ccde1facbf894954614c0fdc3966c149373f7f76af53d1d3db30ca4ffa88ced4b12221fcef251a0eec8ce39e0a9921cba7d3e39e5868f835cda956f5d03a56106362acb88b3fd3d1c8bdad5c6b04de8fb17464a004a551f40c983c77419bb22b47618cb630062557713d4cd7133ebea345f898114;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98b9b0b9711e4bb67936a98593b4625208b07db17d7c668654b5ed6bbb52184bdc3add556eeb6405349fb7789961eba4f6a51dddb9027333f78aa488fd06d07c95c4d3bc82adacb97f59daa76fc01b5dc57afed896192a3d0248329bd3fdf2039ce65b1db98d503a81755234d5f7be848ba7ab19f0e070101f05f189746c4af1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5a448ef928b3ee05fb3e446528c36803ed9027b4649d8b974084b77b93db4c217944ed0b49f8b8a00d9bbdf31d9220d1661788d7d3e75e43a97ad33e0cfac4118c4ea2dbc42710fcb61563c757d590fdd0f1c82f09a76af3b0ccf239d0c9c3d4f47acc352fa90d3e88b9213d5a467ca7a24f77b58a7e74ffe6c1c8083ec8b8d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dce16163a31d6056df81073a5fb044067c629cc1db468b5c267c51ac70b0d7591a1c04d3a60d82fda9d89e8b0a1f5ab4aba3635b2868817b4ac23af5785d1ed44af36a8e71efe3e7a6ded4cb2bd3c867a6d7ff23a20d00c6b27868bd21ec8e049cb517869736ec3e3e5eaed562af2cd56fe6b30c8181832f4f8fc134bf24170;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h482eef9b5c915e00c6033c9c87cbafb38b97b6529359087dfc83e99b4ae345bb64e4d674b0d45fedfeb3a8deeab3b00363a4705c96bce1c9838f6decdb37080788ba3e6a8c80318e3cd3e1bbc5d2f32a4ae02e1d2fd281d74ece72870314f074cae513ba66c37c695c9a0cf8037470fb242574d90ecf051e29c354f7d638bca2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e08fbc989b576f0e8004798d999178d6206e0e9912656d490ea10c25a81ed79fa42471c2222ba92cbd2e1b59da3d749d36856cb3dcf29e08bf3461207a0567162658c3d4a50cd747b5cdea8098489eb5ec4503450f0000e389fcf17965c6f82e5035d5e3434dd58958cc4d8d5c2c3826dafed5af23885e3f85a8af0effc27f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9671141e3cd77414348a2b176c39fc1844204150ecb1ddbd6ad7b67995981afdad60521c752610f50dffa15616cc6bbddb3411ebdfa81e668bb77afffd94048d5670bfd4e150c5cfb247bda94ef1a455d2653b0d1fc679ef84f20cecc02e6650a962adfe267d03f24c98236f8ac9b2e5b730d2883821021ba742501eb84d074;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h116903d642d004daaf56b14c9190d9628d8dd8626acd8b393fb3bb40daebffe9dd359e9efaa890a15d419a762decd6e74a1f2250627fa30821ec62b9e5319c7aa505a5c2f44a67f7a6bf8ea1d8ffa0aaeb5326d670d27230dc1da910050cd5f57546c6f560dc18d8ccb9f5b4d9972c7f16add16561d28a5c8ec29348a36ad02e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61d8d0fc30dc3501cd88a1e2dc1b8bae6957e10512e0d84f64260f553a54cea50cd1fe8e95e7e8a68320a72c04c38c5248517c5b3d15393bd175f933367f2f193f1da02ab8f8622efa7843d76ae699043ce16a5dc8492b2ff7eec912f0fca8e5be9d41e5badc4ea9e446c8da0249aea5b5dddd8ecbee419ca9aefe92de269c2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha04e1206da13c018267877d7f5a9a0fa0718c07a954fb99d39ab2f872eac5bd2a0533bf54c0955179011f6a8d9df08c44ca3773494f5c01e53f447b449af7196830fcfd42e3734facf4b6eac36cd7022ae0992718119267c5f6166b7fd5a370b3d8e7bbe8516b02b8c2d1f6bbbb884413039675bf18d71d5dbd2182be93ca895;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he37d53ec509641dbb150a0134a9eb7b37cc98dd4e9856eea5e51e08b998a13c7e6f6d120b6a84fb46672fac570fc25e2e0e8105dc38adda83cccabeca6ef02c202a4d67abbf6a65a271f8e1252b593343303df9042dd554df16dd302197a06b10bce34d8167597ed667942b424cdeaf13bb380d4c3b54407e378c018ceb52cee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fb09bd093787f022334a34caf9598138a960b52b8d1d4f72f57167d8cefa1b78d33bd2c21a73eccc26f82799bbfb55ea6cf8ec31076530e8b4e56f6a9077e0b882e001494e57f7601f1d6e605bed62d3e8462c9bcd2db5354bc46a430be168b321a8dff2fe35cc5d246edee15dd40502c2d570f307391200877663c6272d2a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61ef4814972a483db022aef7f4d7924448361f18892aba073acb8e07e6cce1502af3a4ad87738d44e1807a3497bf371326f2889debfc9a214942662806fde9f68a08b414ee166d82d02b59d528c83703fe3e78920a44ef64d61cdbfb5f6575be8c3d3d91a9182a528c4ee4bdbd7157a05dac7076e0eee0595e3eb34dd656f7c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h564dc14f0f19eaabeb4a61abf0bdc9bd6ac6c57ff2e55e28194c1c5d03a7680023e01451512dad644b2b602a081ac658255d992c545590620e5a1f135a22fc715a7ea762aa7fd71ec32b62ad12f4b3f1d599c4784df6768eb50582b9606fba44e3b29d7066c9a397155a5d350b525f830bb8b7db783823f51c16e739b2b6bea0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2640abf249c5216305cb4e2d642fc9b1907aae8b69a428faaba4233872901666e8bd1ae66a39e48ff451223db660f36e26ad2c2505e546f6c5346a1444d046caba59011f61768dcee7fd2ec774638ea961f784ec5c2fdb54cee370e5156bbd64789494ce922f9998110f31b46f1762208ad601fad8cba742b5e77e871bbca83a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9778835654ecdbc17d2c6fa8dc688d7e5fcd18e87c04a240aeeba4c1e23cef33b03a4e20df3695b04992b001252c5847086b57bd5287ff8ded8e1e796668c0f7ae9ff0bd268bd1d0c0ba03e811bc59015f4e12088b5f2f03fd321d0b1a74a0e695bcde6a5d61d1a8053f39990ef8abdb50be5d8a9ba63ed99818a938b403409;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf3863f15ec3d70eacfb7d5cd8cb8aef1f3e312a947e5aef6b28d51caa13d02ad315ef30b3949de68cefb9e7240113aa916af9d9ad5565f10fbc902351ea28f436b1654460b1985903cc11ce40637a55a4467611dfd292f5970a262fe6b456145a351306ddd3e2b6d55cccd5a21e4490d76eaa77995606e009707e4970fd008f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6c5d09e30a368988489b1744a79fb290787e51bead59b4f7a1a9925d048d6f1171b69dc0db0d8d8f69023e166a68025c53a983b3d23c1cfd19973626853132889720a3c2bda8ce5639afadc1e4387226c0b19968ab8ebae6c2ccbd87d4140820cef5a1d25860b6ea36e191c644e820948b43ca157f986629ecd65e6413854b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f7988e2827caf32611e5cb75abf49ceacca761a6f810739bbbe8335049ad5ebeebb0b5085403efec45d898a2da4e317e6ce3f5c1da68abecc3cfffa3856c8f49860677fbf599d3e83318238a9614c136f04411169a563f6d79acc4331109fddd382342a7e30d9440096d31bf9a7a2e4e6eed757a82dc50af8f98206e24411d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73c0bfdb42c3f6f5bbf5ae58475abfd1a3d9a10fbbce6b86fcf280733257279128910b7f33a7e5c679b96dac8dad681f3c47cec40f4c35e5900e3fd9cc38753ac30b50e992428a619049dc429e4881f11bb49d136c4fdfc9ff2490864050ad5f319ffb99f90c583297b34597d89439f414729de452bfed373c61b8f37c110562;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2df3015a2b6f2b9054b0d39f8836c08c450fb7c93cf69eabff4b95606cbcc5d100dae949b4cb48227a6f5a2aef5315526b9d0227ae63da8ae0850af585289268b36a5bf84aa20c7059281fa1fb981c5c4ecb8551b1fcf1c9270fa6c7f444ebd3681e95d0552e7a6dd245da1a85861fdd21bd8b8eda72875ed0f06f7c9b9952a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3beb5aaedf100c65bd96d56b78203ba7d50095d3bbbdc9fa76dea3b3ac4bf415daf4056dd9d6cdffa49229cdc23fe6343b075192267e1a29a9b875abcd30833608ecf4f1f1e4e0bbcb961752cb4dd32f3615b6de63e6ad963f5ad42c6508c0c58e7d7cdddf325be0cd55eb145c35e4040eab9a76738c997574d99cda71d5c9e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdca97926e2ff39ffa94b9c4ac892a05507f4c231d51962a4e2ffb061910e3d6b74671c5fcf161e9d621182a8fe358b1f45dfbdf458a9312cba0c86f1330d6184686337692db99704a8865e0e8f4a0095b81b79836d07a42c0451c4305a7d4f5b155d3136f68f4f087dec6a771f8eb260865a27ec9392e30de2d493e57ea9da63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab364b6734443873c04d54bb0f61e7aaec0a957f9444a7e5a10bfd07709ac0702174c8b1d0d5aa983c5cce6245ee7e23e7b1ac4873fcfdfc94d45848a30df8188c7f4e940d03b9f79465f126a93d4ee3d674594c4d2fec46e2bf32c2b4e26ff1bf492be45489e7f1f8c5e06219830d084e218c966bd4008c36e932cba27e30e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha33e9b7e2364311d67140c41ab988a48acbf66ade185bf8585913f0ad5fee99be796f339282b6e41d48279217a4eedabf396c33bbe0258a6a31652d471fee959db41e50218b46421af0976b54b2cb411a2b0786d1fce6d9afb1d6503a949229cab96afab5f57d4524a58a332af116a9af1617412668794dc5a7f602bed55221b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17021835fca7213fb94cacabb3f71a100087e69341f46e7d16c1bd73a7228224b74d4dfe5b7dd5cfa14f0f351171b85eb1445aedd6208d8c1de7420cb6b548aac5487d4fb53c5a00d06c2604b38ed5531bae9f306cd723f28e043fbe4966108375533f508b08e762ded6e6f455522a541d0dc21df520eb182ab9f2a0fa759c8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heddd3e3b3878f18bda60279c2927c6265494c19065928981da91dbbae3a800b6411e0751f2cc0d1996be821dbe290bfbad3e518b8257fedb7cfc874ac66b845765365e35818bebe3e74d2d16b01fe5970c6f5410bb93af27d7b4221820ed5ee575a42f39d786b1e1bd60a875c975a9c62cea6bb25d1d9ac77d58098fec3fb085;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfefd3aa24e4fdc187b8d005318db70c906ac97aa05243139a477fb7eb28a05774910b0e6d2d2fef63e4c369a49f9433c728fad71447d0929602730c5cb4526234fd38b9d84586f1eb8396af1fa6570083e47d3c865b0343e2e563b7c0fe6a7118bf31fab733f1b2a22f5ec346f4a2889c40bbf4aa5b8b496d7125639a7ebe709;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dfb8f1c427dc501672371ced186cded32a1641514be58bf2ac1e5ef088f815e39ded82b456de6610a6481427da551838a4666bbc7f857a0701c89ad261d9bc9ba48b10c01bf60620c7a2d48036fce7efa91312ac79302e4b824d476e8ac994bdfc663e6039d6b6597d0b6dfc473f226db913b6b14c8e2230b687b32deb5e09c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce42d7ad46f865dfb705012f8b9dd3b213054ad76f21bbfb3c16740a9514327e4df3e8be9263fe811f89b8c84224ebe1a758a5451c2fe4d890613f4321a8231dbe38a3b2feae6ff0617885aff535e26bd9866dfbbad1ae432301350e25d7697b21737699325f436cab69ccc9336aaa4099c7dd5ddef99412551866d474e2cfff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4c8cb8f4d31fe8c8e2428bf038617d061d5ac80f5b7ba3642e2c3a73e66da254e250d75c867832557277ea931670b19fa39b19e2a4ddd188aa7ea131bc6618141fa6f7c437896849740bb39283bd73e12218f940cb102e7ebb16afb9f9bbd06defde5a84ac06f5b8d2cf8ef5a79ba345055d70e73406426a4eeeb7021b11a2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51811976c8dd53bb4dbfd6aba9271cad0b0aae177419766f8208e467931139bdb23750ac5fb915836139c33e683baf3fa36ac69590392d4d4ea01453e1a7fd1a944b85607f7bcead56c9a86a077bf50f98dc0d47a9bb8a088f65fb5932adc1cc4f4d8d818d9f02bb7979e19960fda6e3d7ccc3d8d3f161228fec59bf3be8f94d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hceb57b017116de495367bd60db0e02a000226f27144d7a5f61c7a0bb2e569ced205088283ff6dc9bb9559d49eef158eacd5849a89b7adf781b57b9535be2d5140c73a2b13095b630bf841c7fa397d995f50031ddddac7742ff6b7404e3b47c83b213d2e2fe999d120e40d05109a5acfd1ec0cac15c1b79592b7784d927d8dee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacddd41292d1e14ae190bb26278fea74885e09de2790a3c77886b3df90c6bc7f250aa232f8205fb44e8b376b774c6bc1f92a0eacdfbe9d205ffc5cf65fdb02c1da2e9a88540cd8988aa8f69cae493527b612a3ae14d8e36840027e48eb1f583a6e381e9e9841e148081835c744145cbee9f929df06e86e595bce01956eae2d87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h272b9509701be8fced4938ad711adb03089a9554b2905d2c469b370d9ff776992cf655cd555ab35d7e2140218486a7c7b096d38da8f167c0903d8a7a9efdf7578f7d79cd1a32375cb59eabccce6ddf8f0100b3cd9c8f748457654eb60049bf57653aa8566de13d79b98f6d768e5d4b32fcc5e38447e0ef9643115818c16d8cc0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9455d898838ffeff91659fe48b863b05252476e81ccc7d8b722a8de8bedd03769567fbd23280f781505989a2634b638cc09e77ade1064f6ba62c5f113606696d876fd850bcd3e8fe1d5d595a8014bbd87c3f9608a4a1aaa0df1f6ef1ca13a1ab6b25b3fd938dbbee577df9bee6c5473ce98bb2a766d089f683b7f5e902a5a4fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8be26f72233dc17420051afb9f522df16c03a3864083e471112060ae3c43d5979ec24bbb8ae715494536dff12e85f9d978ae3d5dc16d2c88a6bd5a08193c938ed40c726cd4f1aaa0334bba54851814f71d1784fd66fc7b83f0e1f403ae5280867d18a626bfa5011996c7d278e23e61040a26cf7b4e9f083b43b62c64b05e85d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32aec910c7496e59328d7184c5940f0b8c25236b8376b79bd2946637419c0127b2f7f98f62d1315915a3c1ed8b5d783feb7fa14716ab72c257ce76659c21a43f336dc04093698d55a3b73bfe96dea616ac39f8d508b453561cd010ef8a4ae2a7b8c1ed636064bb81152586d959a94ce5ef3530548c20a73a772f2cf9d81c50c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf74bff06b17b9e4452df07b7e85d231cad9a31563018a73efbf3407f96d7b58fbf8ab2005c785996ceb1d9a63ef5722f3f51c872634fce1965d859a557544db2b619c470765dd82037437c5fc279e67c574199c58a7a8c604ffdb99bff2cc3078d8e5d8aec07e50593385c7eee0eb12bfd85cb32b2f2d524f94c65a6df7e00fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h653e275d275acce16630ee43ba16a82f0ca4a288f0b965c85f270159dcd95de1a9ede21070c497f26c0d7962020da87035fa4fd80277a5c58c500984622498d1841a265819420bbcbd6adc6defb52c6c1a2e30cbd330d200a6f06e1b65af38f765124e6c9f468223c09bfc5b79f336e9b138cae9883aed9d76e539a52d7097f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h387ddc086e1cb8a68994720f15c20008add1bed7c8d4eb271faf19d40bd371b708b91feeecaebc440d15971551557731b25b758f758f0c512e138b030d000daec92a1ea03193b9984bb4d8d349477443c7d7f877e5a7476d33830e980ab386caf48619861db984e8263200da928a11ab82da8110deee9b22cfee20071f20595;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8101950d2dfda1c7912b51a9a09c1e11e624112d823effe5ab2606a518f74a7d99e487c85bef518605e5d1b843a25ea8154542f9b861252e23d818b25e1faa4dda4a7490eb003bd2bd2e65b102a6eeee3470f628500cb5721c3c763fda0915221e366a301db8069cec93519470eb6117a9477433340572a857be28d401b203c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48183f4c196791937d17316f88c168fdb8d34c220b930df7c652be9a9910c7abb5576da9f8f63a4c720fc996d0b366df43663da4c9e95eee98b67e9fee3935902820c04b94fef7bacaf8b13ce1a8ab4430f5d38c7d3f7143b860a657f5e00ca52def50b42c110e74fe301fa23ff68547d6ffb6e2df2045206f3de229df23eb9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2492a83d766c63b4bc6692b23dfb0b8805a78b4ae1a7a9e14390c84cd2c9670ef988de0d6169c18ed653d6a9c0cabe7decd9375e4a23d099ec56648eb5681b731445664ce73a0ed166883f2ad9f4b2e6ed90966f6bce3b6a181869112491026a227eabc19fd4fb672020691cdc2618e7013dd30fe0c4765e3ad61bb7919db34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h629acbc20a0d59f7f0527f84a6b2e7f8335faa06b740b39dbb628bd264586fdf9edc5de641859adf23ea69ce8f7b0ab9a2bfde7d42dbc23a059f766f41b6fce71efb59617c83a1cf3349ad22fa048d9fa5dce93d5a1543a10813f226d6b64850d830b0dae742e616c3a230f3193f3035f10c8deeef275f1ebe31a67b6e9ef5da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0a37bacbb2b6e4c406111169890a20734b43dd81bd729bb31ec3e2e5784345d0b270aaec6b634c73d9668578afebf6c2e4685a4450a24a4b2f28f38396b39f1b3964309d2765cfa857a6f493e8383c623ff2b7799f925b1f6baf2d8378669a4468915d2485e225209f8c007b2611dbfafae411e3d55265370fabefdc3c26f90;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54d259ddf52dedf59de3cff6ab20048fac7215bff3ae18b2002b7c7386cd2520a21eb5896e063e3489c4b9c2e2a3dde9b2a35025dae3864a45c7f600af3c787a220cef0ea47bb9ad27c7c1bf9b18641c54d3ee94abea22509a9d625a0c5edf2dd0718036b73b80a029147ecaef416d73b4cf5fa5ccb2a81a73d001843e01b08b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb9114807e2b10ca3be33de430395ae942b0f89d5b38408a192f311332c03753a27669fa6e6522bfde11818ccced25737b144b828fc6d94d6ff59802748b47da9638d2105c46e8f42725ecabec7e4b0b3cbf814138785991757f62bdfd0d21c170037ce3174abc94612d6457cfbb8b08dd8418b7efdfa7ea2d7d545c39fb8a43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5d02ff0a1c3a0f3d58a0ac0f8f540f9c358ffeb6b904d92be13e16e7bae7922d541ac5fd654973abecc7c0eb39fb5b884f11e68f2188a724e0e6574b08f340cf213f390f62025a805ee0f808cc7d894f78367c48355fe21cc39d794fdbf974dcb6a1bba34ee9f28e39a45422a62f9bac318130bafb6f6ffc7572b2598fc43a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc659145183bfec629aa649990d0cd19d28240879030260ea6169fa6bdc380296dffcb114b7a3d387c81fb84db70bee6a8046fd5c77a2ec0bb2bbb9bb686eea633611e192a52675bb74179c7dca950848f5992f82ef6894bb15459dbb40082bceea4c2905f8bce1872568218c4aa42c42499b8eb40699294adde5f3942f15e674;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d52d5078d44f092b71c95ff998ba76a347e455a62aff83d4a693b7ae3cfb6f95f9dcb444fc9232b21c67a960415d05f3974c0894c7b54affbec1fa5f5ee7723d3b6a81664742e90a5181ee51e5d1bd683d7e718465882598a84a029ec46813f068f6b9f674feb995aba234a8a1dc6299fbe7693d9c81324d4bd55fd287f780;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4e6a5744fd8162e03e4a63a0983a453050774e0844f8931600b191d92602a811fd3b4bd8858628212baf926d4d1ebfb3a1804b37e0306aeb92c9f07044ed05f9bcf820895bc93f888ccd72c05ac800bb32bb964e24020cfc52418551a4546cbaa636303aeebe41466632f846b827986c3db30e07d0b6b8f3a9e5e1dc85e8023;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h697e6fdeee627238b5e60b20f2950dabf789aa394b4859949bc947e0f56ac49f2af1676a7e775e2fba9cd2d00f9b5d53d48d22684bb2084afbbac009058179b557317f063432ded047135b9778925a9bdae50a5fa3dec868994d9126d753f3f2c754e14e1d1f1367d806ab57b31b76218ebf7fd9502471896ad0fe5bd7bac2ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5637afbc5cee8956ae161528a055d8c63dfe66af90741224c36c69bb28df9b2e092354673a6e1a6c499417621f5e4e03351ed253dfe560ae7b9bbdf42b3b68a159496348240b673af23d932ffa5c2527c15630b7a9630f605deb6eff5a3d5133111be7da25fbff1198cbdf4f6b2dec2acef4ce7ffc252711d4751291cdba03e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h540aaa81182747bfd9c8d7d9b11b0d51d9984e6e5bdf750319caf4eb6f43eecdb0679c1d7e27bbe0f990a1bed965316144933417352f186ed678d32db3e45fe09483e098da30bf13ee72e897552a2ad320a855ca5b877597b5d3251ffd9d4220a044f7c38df3ec600451cebf472fb882d1b5e0cdbee7524d0af2f396235f918e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd03a8caf66ab794b6d520915947d7922652503bdfe2b777b495aa223d2c6cb0d271ee11ced68f4c286c117431fe02f7ae70aa4e6e8a4ea6beaf326d87c4ef95f441e4ad0d30b9f1d71da3359660b2009c4239b99d42c9e2a3a898fde05b906c521a83b30bde413114efc7adb45663207a0cf09236f831d79558c7fa6f2ac89d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf7565b98dae9f7e73ff39dfd83bb59eabfbdd4bcfec65ec7bce5072d39594d7b8bda0c7cec9e3e67beb27faaf1170661d238aa1e089324c5a2da80492b173c30ee5468f59603649c9a5f7c7076cd8923326f68d6de0398c42acfa327582c52dd7d8c13228ef4535fbfbfb229ba347d6fdd44128933541f5b3147c01bb5e7a99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70b9a00d6924ef062f7e9882256a4a1d0ccbb4bca03e27752eb107c00f30ab25083bef6c1b32cdbf4a693ddfd4daafed75707e00ad39d7208cf95f12d6b0913ab2899e9f0d692769119140726ca7b94573ec8281272d1e3a88f8ec6cf61f8df98c4b2918bbd2b2ff41c4483b9b4aa0b68a8ef6a1bac716f060206e13259bb7f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f447709f7b0bd571a2ba2334c7484df8e6b6be967984fa25ede79fcb0d54949c2582498c938905a2387dfb9a3c09f1d2bd0f57794b4552eb6e8a8be2c2da7fc328c3b36c87868f56b20c0a8d1148d11e259d5aa8ad9d3b79195935dd9c0e46a28568b540781791353b45934bc8505b15f45b2f8cc00fb000e655914d5f7b1ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h653112c1e9499f58d0172269d42a2c48c27516a4dc529f1f209e924ad90271f21b902d7285d1f108baf71865e44a40da4ece169813b66a65d9483531c6f001589b82f3f77258454b1d47b3ae4cb7e605cdc1d856162a8a7987008388b2290debb544a5e0ae1379ab13786680505dea90b3c59e63c65c476b57eca0abd270085b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a3601cf7509737a8f1d584d25283d0f4113f91ad933c1ba44aba70e714f529e9754d59bd5fa415b9ba9eb966b01db0f884d0ebe3621818bac02239bd892ffb2ebd851dbc56d5cfbc4d27b4963b25e7901af89ec17e64347af2509ee919c87a386e1aeb80a98b567ab09c6cf9f5524469eebb2cfeabeed016a2eadcdba696662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfff2ec8a5aeb953c6dfdfcba05096ff8d2ff413e0497e0a87d7ec6a1fbc642db65af5a458cf51ff8a532c42be1e812f560bbdfbe25349b0dab0dbd2541909ba1f7aa0ca814620012beecd3bb0f294d1c17b571641050d89e950ab30d229bd242c34adce0bfda2e95223e024514eaece642636bba101d064b48cab4a7746e3c8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb31557f7199ad46b9aa849581a505bfc1e8d6aada78527969bfaab3b602d2b976739f62b9fa6a54dad41a31e607eba3c5276993b93e769b560d68d5c08edc1081056094a85aa3d15c73ff6452a77719dbb44434cc05c738a0d379d4c595395f3a0e5411c77bbb9f7e2cb7dabae39e8779c3415e1799fc3b8e1a8d4ae13efca0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ae29b2708fedab11ab7424b11c5ad401dde4fa3cd8816f022181bc1a16d56967808c0f8bddcd35976bf2bfc0b488de5120cf6b927dbd3858be874d39a150a4dd70db48eb5241d03760e9a648b6c91a96ebcb69f7cd5c5ef6fba791be5d9d2ee47cc90d15b677e47d4e14b917ba15cc2ef4bd27e51b38c2dcc49df4306099675;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf671d8aebd9058f7727d1c049f9f595d452ec63d6b9129aea7cd4659bb22faf4acc4c902478a7c4f18c2ea002295bdafcf57f8d75c98761aed77523bc5d7e20904a3dc9534e067a8d5ef13114b1bce31a9b3816261ef032bf01b7d8f480785330356aabb77a5794df967c375a88a393f0e0607e40ffcbd41612883bf6eedb780;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4aa901a1839997395473fd20835b436375a3ef80bcbe128b72aea7ddc717f99cac1f2ee8cd6e6558cce83c1cc4c898d441397d0ac937b77cc7a5f25dd68d2530b1284098edc2dd0934d0d7c136dcb9663b2bd7a3f54bd3b87b9535a16d51231fc33b18a8027f06a4cfa6a562a73bad13314bba6bddf6a15f9886ec4e92128af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64357fd0247d2965a9e85363ffdf11c6791e8cc90e33009ed0db509b0dc5b4474864dba2acd7794109e5eef6284647d4c7b688db5ef9973ab12a00a36c84952ab75e6f3be595d045a548d3264eb4c104652134b569ea24285a5a407882bd137affd51035ca8e2be574411c03598bac2dee17c1a179bb45fee6bd3a1ec2b98e65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a88f097db3212f6b85309adc4db077d8e55d768cccb03ed92ffb612a6d7de673c00672a67dd8b31bc3934d209d84c5a9e7bb5e674c050eac505721d1a852a061ce0a66f9ce95142f98b2e75e296caab8318277933f31fc2e3160c5955f07b1f64200e156fa3cec876bb1d034b9cb86c59faf4080bfa33c44f111f0edcf7daa3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c096ada26fe71a77619c9c2bc9124dbef57e67b7591a65b834c590c1575cb496a76542a0148ec44879eb6376356613376371f4c3a7fca67efacce3b4e161fb7b958454d88c90d73dd58fb412fe28f6136b30d1220bbe13d059aadbc2004e30d65819003d9781435ac96a8273f81a18b430f9c40b47ed0edd55f5b60db4739fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e28b2f63129ad5ac28818d40a5ba0297faf2df6bae3a1c407a6a271fd3d290f87ab377deb6b03736013c41c619d78795e78a1e1f100d713b5682dad645fd849e3a70cf233773a29bb0c66b112a79be8c83fee14a19aef3febf3738bfb4d584ff81f16584a5435b83793c5370569e1817baf7b4abbe8801e96a22d96d8bda164;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f0a1a0c24ffdcaecc9851228e1c1da196aa27ca5a262917aa76c0a3bf2fe74dc2d7c66d6d0719ab84db64acd6b0e40d680c46737185378992abb78fb8a8eab8f672eae2a02e90f8620e778cf9149d7d231bbc586daeec6e8bcf8c0325d550f8b5f84fed50e4ee227bd9a3ce6bf28ffc46d5be36e754c73425c42fa59aff5186;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86a495846be651ccedc64ddefc7d9504a1966eb2e96e7dbff084bbf3a0e55cbde4ec6b9855e8d024c62d73af619606d783106b464546058d2fde5896f7675529cf98c48c4b179ab1e506291fff630da3b50cd43e2f243c1e566e4e37024b8d1b381bdd9da92e91fe44ffe8c29cd3121da60e37dc519683c929da0283e193c150;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89f58361196689d0cf7dab8b618e65a25d213d288832d51b51e814501cff600e4704b38b906974de8d4cc35f2ec9762ae3ffd2ccc83f1cedd5083c4fee4e3dc837726f5b433fdfb784d28796eed693c4352110d43c17913aa67be04f7d60de2627c0fe6f2e21a0535934963eab3220465c93befcda672d76f8a2d50c05d55cdf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfde8afec1697a3ceff4ea601b1b1dd89deda7ba3412e58c869c681575a124b55ba78c2f324349555f91561cb4d2f0fcd892846ce2fa2b74dc5842cd05a5991e9d42bd7c2c47d683c862f9aa70bf4ac436e7d388b32f16a973d738ded58ab96a9f5d0a45620af284a953567ebd17999d3e688f305be814b813bee785b90575f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65a029521adecbb17304ca612cc0d140c3efc14211afd31091c63c6aac781066d3af1d959f75b71fd273e4242fbcfb0a1e31d02d484fc67acafe0706d08550c620ce197c0341c79f17a759d51af25dac03b4fec9aeca2371fc2159f4474a7d9052f7ee88bcdcbd3e89ed2eec3bfdda48d5116b615bcce6dcfb53888c2db96f07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc09bfbac97c40b0376845cf9cb03df9fa3af450c34e74e7a157c01724a6fe6c034492fc2fad09478b6388eadeca55e243102a0e6090eb42b3f2632173b21f89eaf144a4aca4a2481044a6daefdd8e037880e4109bcb3c0898f70155d4d2377a838b288464bde3adcf02ac6edc264cacf330ae4a18651c54b1c71ac27352de529;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc54bb1b84511f4db840baa935e7b30358ff920d97f840c736b9146fc00f575320b2c3f8455c738f08ddf049af2b946210ecbb169d52a11fc0630b7f31842ac7aab315cd6cb9fc06f6ef0b51af295c3175a4c94c99a2892c11bf1ad7493f51302cecff375d41404ce45132798a7f9695c7a1201bf5119762aa127b02a91297e75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25e47d83ee05c30f7eb7d5057158f9e463da11e5e0e2857d575023f1f253033a73dde6464c1130d2e970671fa5aca7f463218539d58e9f6c987d593ef934f67007f67c8ba80f826ce7641fdc35c53fa6b0c30f806741b4fc9c0d1acad1a6164bc932bfbe2a3b30ae13bb52d495402590f44931c3af8975cefc25bf37fbc78a1e;
        #1
        $finish();
    end
endmodule
