module testbench();
    reg [19:0] src0;
    reg [19:0] src1;
    reg [19:0] src2;
    reg [19:0] src3;
    reg [19:0] src4;
    reg [19:0] src5;
    reg [19:0] src6;
    reg [19:0] src7;
    reg [19:0] src8;
    reg [19:0] src9;
    reg [19:0] src10;
    reg [19:0] src11;
    reg [19:0] src12;
    reg [19:0] src13;
    reg [19:0] src14;
    reg [19:0] src15;
    reg [19:0] src16;
    reg [19:0] src17;
    reg [19:0] src18;
    reg [19:0] src19;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf6242757b6c28f75c149874e47588bb3370f336f5c5276e7c42ebfc6a700b3310db98aafb6439cc26a6dcab99d73f494fa9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fde414c85f472f30573c33a44c44b404bd7ff2652d4c0e227fef2a134fe944669bc7d77f6e2ca7bc96e95c9bd4e4b3dff45;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9f4d94a0db763627fe6061910c55d994370f3f333d3b012a7ba40a4feaf6f6af19e5ff5819d69f1edc1a54367b924fd1d23;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f7597380bd9e916587a60ce04b7f2332bce123d2dbae05f457cbcf52388f425a91a4f9cd26534825e7cf937f4f7dafdee7b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30bcf5e0ce778366db38d35c0d3af4b96a5a0fae8f3c6e1f842aa9a00c3334d1a09037a2d3031637a8982b00c1304adc36dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dcac2299c8527e11cad6732ec41110ef34fbd0e9a4fe9f0ffcc006b74f9e82efcc770e3e816c01cc4e8c8c07392c73f610d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82b2d60662ef79b75d8d8aed7cce9d78bc9ac6a1788c6885260452921867ade35108bb3c316e02677acb5448e035535f4d31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46d383a8470e324b8f31c9c31ac0a8ec4e34b81dd7e9c40b4a72f06e8e290d2b16c1d174a0ce53a0c4b01aed6c6905975658;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb74e879628613cd8622f17310f848703f459506338b5cdb1991844c0b83da59fcdbb9280afa1f037be1408814d100e35be33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf76519d768fd751c9842e6a9ef03d7fa4062ebdbb0d9731370a6dfc045fd385656aa565e9c2cc8733b162440852ef65768e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heedce81ca00881477e6766cbe09de6debb63b8c47b647d78739352d65488d7cda66964d5c0bfb24300c66c6ec5152d63a2e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc671887afd6b8fafa725f2457e4360bbc7cd3092904b61b74d9dfee7baed9fa80024f334fc0c65186c740571f43fcaecf955;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdad96aba2d2db46c1d56fa3d2f6d970a053939238db959fedd7e30e18919a9ec3f367592f20310a48272afaf1d9c4ffe2fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h175deb2d2308e8e0499140160f9540c6693a5559729a29ad01aa9dbbd427f938a4b6f90bab8f31518f1ea21224844a0c0e82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3c281845df5764260fb1877d54740b0e84df6fe608dd3173acd1ee2235dd445b4d2704cbdd008099f3ca54b953154ed2913;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed8c40775a479017a3db7b88a3e7fbcdda1548eaa7bddc6088d8be25230f72354a77637f9f929aa963fb5ae1294e37b68f35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f5d456cc52f2c485d62baa81342db04b751e2f83402dd37e1b4cde225c284d20d3f901b6e536517c2ee32823869a3be8765;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74b89fd0aaa51973f39290510bdec33226cc62f58649ae8c407feb85ff5ca15d09ff250485daebac627655078de96784a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bc86c50e96b5c1d11149345020a2dd7b683c3f29d6553270401c670a057feb92367ef63b951d35cc0878df7a001a2ec00b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5398abdeaaee470582c9bb6a8646b611632f7283a28c5335a5c83b168236c1159425ab076e3a2ebe276246166cd54a3aa364;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2edb469595edd74efcaf846d10eb25d5dee5712f19899cab8eac7da122f10cae85cf169a3ec335f7c57dbd1a3fbe9c51151;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc407b2fd251655d40e382a0ec8f5a924aa948702d906744bd5898b1ea230ae5e34ab091f5b9a2bee97bc09da2bea81d8ed44;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb5f7e5409b41c8fd3c9591ec0787ae7a187c9c5f6c6ce4cb1da32561396f262712cd3736ce54446e088e1414db05ba65e86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8afe90cd36e067d235bda0c79d2f7a94338d006963ba0aaae6d1c873b662e5afd34c3710c4cede5852244a66d72230f5ee77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27924000611bf0f57b8716cd753928bd3aafcef1edaf3dd30a5f4d421ff00db378daa09da6a1219a2b1601b1974991d7273d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcef3c7432b3237a1a89e579b14340c6e7f44c8f8c4308bb899cbad14662e0d34cbda9e839285860f1f493026e76ec2469cc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcea478ffb77f693d4dd6e3d64411b4448aaa5d3f332650f17bdac526e33927ad54ca717840e10372a653eee216028b9a8434;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h543dc26446bd8dff86696d029349dd650ade9a41168cc663f7990b06e522102069698bbc26e3264491f9ca39595ffa24cbb6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb524258c2967bb12281549ae2faac800cc69c646f37dd167f67e11bedfad506130321b8f566b1059ddc8b013d556f51b704e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15354afc52f700d2307553185b12912c4367711eedc8120647ec7e89bb5e1f87061cf411c1cf1b5c975340a8de6ebb0aba83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92556a9cf0b12e998a5d6638ee8135d5f815b3f032bf7e1353e95773825abbb97ea27cfc6ac4c6f4840ddd26b12444887f51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3331ffead8760531e9b7a2fa8e8937e6ab38b9e43d6337f6db49818ad9bd1c3304b0d97d69e7f751f415d00226ce411abc4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc37bc7ce1e54a72ad261228c5f64790c8ac0f67b2d7826eb7ad5e52532cbcc1e571c4bb8b5bbf257f66a8c903468747ca44;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b87657740c6e811c4628a99e4f260ac896ea7f1b425c89544dd18abbba565188fb76ff205134a7f5f60ce0bf090ae42bb87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a0a6b80234ab32dd02b733ef225de4f6623c5d3c5fe2833b2107dba437da995ba6630a0538b35fe906dd019dd013387a32a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d87a07af8a144383b75b6976e84f0647c1f521f489738e495392edd5bcfa214d8dc175cbc70d21124922c30ec833a2f3a29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81fb8edec6df604b8a3897d3c8ae4368f7579b22e4260123a725b310a20d686bdcfa890aac8052b074109766d03ef1f54f7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c4ce1948fa7bf350e3b9d1c33256fda831d47941d1ee43836e504f468f20107881dc122622e98a8b309c1018fb96ffd8d7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf86715a8aee9436ccae0b9d72c82824d21312579bb68d1f84746228f6cef179a4c4434a5b9ed99146b7b3d6abd71033a541;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45c80187be82db31f600343eeeba8daa9f5794fb479879dbba36fdca9af835c84d99e8cf6ecba810d5faf22efa9dbfd45572;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e8ec3c9e5bf57bf0cbf669cda098f98c35f07ed0ca9405840bfeacb8b94a6859321de1d9459e261f18e81c6142abd08f456;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e781cf46a5fd0632e11bbde9ae5f8ab50125d2c4b4d4b9ddd9323deb2b601dc7627cd1422d73518fa5078270fb8e94f2acf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5810e5fa862d48d392f773c8880c4cc4f646bc9c1b7a5c969f6ef8e2c2e706f3a3fbf3ab720615d530f8475af055348ff6c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h693a42887ee81c3852f3383e5bb1849405cc970066738859ea5c91d9248f8fa1c0cd3dcbc023112304840d756ba7b5e5ef59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15bfc59c47c402f90a00dc15787b17dfcdcafd4266b7954277032404f7f9b7c72372e1e450426b650283c9186d79324da44a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3d725c1e8a7c4811c04cf34624e5298ac401cdbd65f526281959da0da7424950c13889bad3c0f9d5e15fbfbebd7c9ed7ceb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53c6c30218557218ebbca357a7d2b83098e5cd25b398c469ae83d7f6df3ed14f6724b46e55fb5a500501ca1c7f0837de596a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd948715cbd9fd775bceadad47d87dd6193df76739bffc21b21d7ac46611817fd73de414f0f2e315eb8e9da21732dcfe610b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46644e1c2b2f8deb9e9e8806e0636141c68e94c9cffb647c511d5d0305cbf54db39a826f8c3d3b1a034bf6ae8965e9b0bf9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc3b449df43d1ed171a0f173362d2893bf890b5963a33d4299a7c817cef39bcdc5abf999bc34e199f7341e3951994236d6ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3ad93c483a8063aaef89ae9c317ad1e8dbb2216404e7d94a4f3772c24c325114770a7ebc265c16dc45712ca42bf9a758edd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbd8f198bbf1f451589a37260de8a63b555cc49c3aa81e77e6c3836e4cb101d04f3b1fa363c4985fb447bb8dc03b5ce42037;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7df2dd8f7136e643bdd24e67eeb61eb0aa981337e69841765788e7acbb365511af0890a9b88208084217238fe53f39888d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f5c6e61f3bd39268122f9e19704d6d2f251a1aa3d0f0ce998f4f8b9eec4926407e0e5e899900c8d0386639e927e0591f174;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebf53e9db7fc948e372c36e5ec2e67b6984ced2571858ca84c199bf40707895bf1ecfa9fa2ed19d8e71b6a511c8245679e4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3981ad576a7b25a929514918727e02e9777044fb76e3da33b38923799c16c233dbb5061c0c5d0e207ba5b31ecfc18505c0ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6863d59ab9a4972d056d87cddb953d8a9b2b3dbd4910390940f5ed3639e0fdd3a21ddd7b04a3a2f1404b009e2a7833de026c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc89a89ea24508f19577c176fba05141b1983a4ae381ae74817780628b207587c2f3cad496ef406f5a218f73002a1240eeff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3bc0b0e8c781a22a517b0a036019c0bef3129663dfa70f3c2f0e67ddc4aab3bee40f0ef79cbb67d5c23ba42cc9c0a865060;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb11525269f8ef055cab5e90b570f664a61519dee4f5f4fd7dadc246f7312d84d1f8f7f70fc7ff4809a7451e1d7f877b1b19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0c7e5bcbe6d1c5cfa9b1d7a86a6a14eb6e30f1fb5af37ab762e8d60f4ab79d7cb73aa29f93a1a8ca17cd13c02f9aafcfb91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcced642c6b7d43f77f1ac3db9da1609d124413768e5ddeec4c8d575207141ed484c24a70714de65cacd4a7513da3b5704071;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f2e24798c947d90eea80f21f4444e4c54dbd08629f76020c4442fcf7cf2cfe6d20b0ab72d26586d4f7c8b5aed5acade9c33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd45b1d85e278574d9a42037d370d937b70b3cefc6abe254a9f1acc12f53cf86a4d719caaeaed61dbee3234a6789c6c191a50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b3e3a03c1440210e691c52a2b0dbbeb6c5c25947234f0fb210bfdba7550a489e1ba5a7dcb79620193c02fcd3eb1298a62f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e9423fb271f3189b1ed46771362c1946c7c00fe831c64a70c4a8e673d93a3a8cdfec9a2711481dea4280657c7698a8cf048;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b30c727d2ef3399154cd025358a90fc5c22e31a26c847c6d4278a20f05086012d5a18dfba32c81ccb0005a6d4cf9796b82f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h866169033da473aeb610402328e93faa519e7f01760b66b6b39efb947a4571513fdc196dd100a328679a195d5a10fa8355cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65208c1bfd19c9253387c1b793847a23f3230b01657809180a10c1b26b9969730291aa6799882c9a78cb05fe0330253c5983;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h192f8122b2d77c697977624f797edd633931eab8b1d953d6f2b3abbc7bba048da95fddc799153add83a4a9cb5d3ec1210ed2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc01fc7df6036ecaf1b964734ccf30a461a81e02d4aa3de8484aeea6d54474fd0c9002777803c5f23b66b7b76dc38776c0b64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h767c6cb53f759988cb704608e9b16ce353133c49800ca86f794fdd6915400c91fb3af179e67ec72da02bf0358065af85c245;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52dc0793e1f939b7a7eb05362683e918ae7b2e2a0b0a297ce7b5bc7cd00dbfa7102a0b466d933437af85ec59e97ba72cc3a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3c704440e4d3ebb713b239fbe4239b9e91f860d87574e23b6e004de31b1ff4119324400ee7477d5ff8ee05e0a1ae93a38cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h484cb7c68decfea1857bbebc6aad293b152b9cd766ec9eca8bdf60c6537f71ef84150cf0f1b6a5e8d6e3d0cb3d98e2e53316;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h449f13d4cf8a3dd02af75e24139505b4b32489aef4c5d539cf6d96c887f01bc9d814610c63097c9377fda0c24a6dc0542118;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79f0419671de51a47cf4af7ba6e41b42b2c2dd6b690b9491378ca0ba3a620f5950224d8b3f675e1972d43a5f39a456bcabf0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf21b11db2f83c60991e5eaaeabbaf202382d42a4881ec5faa95f9384db431eb10e9c968db9e79efe9a172f2f847af6539891;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68dcbf25113b8674e5dd166eb62ff8b593d18029570782d2faf7d330dd009f738c79b11895273944a102515d1911025b423d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f38012f9722d43d7ec178bb98403b4f167633549d42b4d13cd5f204d9d3b83e808554062eea4eff65c60bc69b50b11b97aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdff4d960e5fd937185cbb99255296c7d9cc375ba07da64e8750d91576ae2a5a31c11ef7080448cfe99a700b011a76d8d1907;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc3d0164c7e19d09a82db90aeb6a745004c0878b8f648eef3007bbfa6dd9e69d2ea73a09437c4c3282870d15f6e0031133f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb213e0667225bea630880b158a80c13337c3df0344ab8ec5685d2395dcc0842342fed87138abad9298cec3a049410958ca93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8acaec351f22cac5e2a940e0690d0c9874201f73d87b62fed298686b30d03ed833034211bdfa4f4f496a6499baf161fb844;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1223b078b13fdf212f7818d52143473c696173b378e41ed0577c00181def72ea838c5c85b9616e3f85a1f37a173e4686e3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb50f0bf10a7799c87ad5ae56140a3a7b2b10830f81b163f6bb23a9b11147abbcdada94368913ec80a87d8ae8262d8f1568fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9360332d443b5cce31fc722f7db29a5f7fba538e3d820dc00344b2849802b855535d86718d1b7e98e9089c2454968bd5397;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd546f3a8d703f35a5444b042fa09e6c87668858333d4795e3e88fb6122cc31f0f5487f88a7c82c620f108d292c72412cac71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95b9d0c28433371d978a05e96ad065fdaccc9371da6fb9bb80a08c4401fca6f3bf6113fe2eaeb645b0e85a980a8417db7965;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h386db8cee8252a72db45c9e945af47c2e3f1eb38490d44089e9694a2896f4955f6ee3132a8d918d5c8341ac69099fa5b988;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7bfdde48a6af3b3390b7f0cee541a9e8bd5ec65d0b8385c31dbdc34f818690910ba9e06146630936171e72a5bfcdca4573f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9586b90c76fe460c18bcac46b04376f200c272a658d1b4d5d14a1671e4a3b08e18922a1db2a105fcf99be30c4847acc4dff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f58c1b00979c58d5f5d117c8dd9093d73d5f272ad152b587aac938626fc41426c46db6111cd2203f019598afc022c88bbee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc452f282f46f9f756a0d08ca6ab8e36f31815a2d73913e1ba822c2478e373efd9f9a5136a4716751d80e72928de76f29dfc1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f25b9db58712b346c85b47a5ad78c69eccf8d64ef45a836d53f6e56aa1dd1b1f179121cbd2ad4752952f67b96595064963a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha547f6513ba78a2007ebe69d99470d6eec86e7ee93d4401c1400b28a9442c26cd6be1bbc42f47d977be584e30c8153be0c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ee1f16f158147f8e1bd67173cf196db239a9c1dcc556559f0b38ee78edfc319a96f7ebe0db271e47bc31600e52f81513e5d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3dbbcbef9a4889debc9c522ac1583c69f628e31706bbcbb4c9fbf7f89dac825ac4ecff2d1facefa5ac9eb257f7f8f1baefc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4777365dfa191bc7b87aa0664f7f7919948ec7558b05dede22861e934c93c15560009bb8f0d4dbb87443823770fc456dc5b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28d37b7c2d137a7d11376f2768f11d9d74a35c28e162972ccb690fc99f1b79cddc8e6baa2059ffbc50f53b7b9af099a9ad2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82111e97a655954c3f0ed1af55244c19fed24b9a7d973757376fa58da3052ede69e350a76a4c29fb8e719411805b6915375a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc53c9954841b9b6666b82e79aefaaca7d6c490a117880ec31c14608507a206de88ba54e563be6a4a9b25612b8a71fcf1b21b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2377e9a3bc22bd27e9be7200f757e32acfc0c5314684886aa1d67f547939bcec2e4553cef33cd117e12eb10efceeb230e52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h276d727f9f5ffbf8e0bfa7d5571eed6776ad5f1851bf9e4f85a9b66c8e3ab63c8ccc6366595ed83b8ab32785546c6c5788bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72e90c1f5014581039109f879bc823ededec106cf6d50e39c7fd1660199735e8e3148e508ed2dba936520fcf77abc7230e55;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2c1257e55be9f4539b6a5c10bf7107e12b8d9428bbcbfb4d7c862adc39ca4f65e6c0929b8365b6accc8799771687969b0b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fe062a4f15b540bd3830f655d90ae9cd93184d28cbcbdbfbfd4584140976d46da0388cfe7921ac4e4abaf34dea8027460fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82a79f7697e15d8af91e1a7a9d0f0e6890b0cd3ed793b5eddcc80c8b6229b0382278d8bf68b1080d160f8946f49e4240f301;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc49a94ee485e18b680aa5e2527a5355b084c53c2433f8616de1f842b92424c46a272575f38e898f5c820aa63ae78ee0a6b88;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h576e8b02a31b29579683438916f84910570eca35a4d7bdc5e872e890fc13a7c856c37f0d54c5cd876224362497d10030e074;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19185b8498cb3401a4ec36f14394e70cd1679250bb58b7f2bded7de10813417959ef51864f59a5115a2b350b82d142a47394;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c5e7703e48c8db98e3f69a34bea3c0bd68319b8557e0722b1dfc8b6cb1e9b633c8d95ccca3be0ed9823661b67241863fdd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca369abe6d105a09e98e2d29688a5768c11d656b1fc3fb722ddd50a5a65ff569bd1a4c8026a2a6198d312d9087ab19dd4869;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e28eb3f9b729e4cce7aa34d2011007c6bb912b91a7f989a466c0780a1f48e1add8e4c5bd43b1c1315f4158169e97b2b4b19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h815c19e0097a8b75ddab9ced48cff8c52e633d49fa439d1461a33870901519ec4bc4d36551e1eae1ca0589cb56807472c65c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h416fdef9d4a5cd30ca64fe3f8a432e8d0dd2dd4fca214850c7c571dd77eb329edff4d161edd69ad633c02e579861f7335d0e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff3d2463668e575b6c2f715271d33f68e13e9af76cd7acea32c151bf8214020cf6623a037c7cceb089196199749e8a6fa0d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34ce12330b9f9ca56a8aedf36069b1fd95a284b0ef3a2a5a325c1f3d3cd4e29952ed4f097831098d1d6a247c03b9850735e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0bc71e7b6e80ed990541f7522acb37b65a554f75bb35ca504b46a309e3f9087433b9f7215b42429db3881d2ea19e388c8b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1919a64204b05b2a0848f4d56e35400c68d29f2be0aea7b94b9c98031891d0cc5fc7bf73a8e34721298c59bfb48c206de18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e664cf5f6eba4d801bfa9863e70a264e64055a8713d62367834b6bdce6f0dd269d08c980d0851cd5adcdaec935f9a09e3d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde0c6c8344990a5a852f677533d7bc9229fa168aeac1ed6025738bd11559fa8c7ce6366403f6d1f1d1ced46c021bb289581d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h717afd3edd480b43fe8f1d24e858e8796d16b9405411ba6d3fee7cf7f5fe7bc9a4097acc7f30b507e5a15606ba2f115e2b36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b87d8700a4adef02616354ad05bd0103a0ebba19da52c48c2d3a741067d3e14fa0991f2b5bd6ea6737ebcb2466b02ad8edf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h247460f118a41bb44b2518aa471d85f9b9d3c36c02bc7fe491c36346f5dedbc855b2facf8873841b81bd40ce7fcb580f3db7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h911349592017de9d1d790c86c53dc14fd31fcdbd79c30b9c1b5a7b31671a3fcc718cbd8927d8de5f824f2dd72b7c7506bc83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92aa372ba564b510f83d91c419c3c906313dae2325b1abd9f253b0e6a970980966c8020f2cdc9481a62324cb061fbd739016;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6e35bfd0e7755a7092d9ca7a39999d68181900e828145bd1fcc2e1b9ab4729ebe75454fb2f337cd567af72b9941b14ea4ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e1acc0ad2afa98d4504be52476c630bd4f43d72f63d58728cb915d97191157343f89db99fe1335339e01c6cccdd7afbbf81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1abf1f71cb115ac5eed321b4708d0a7a81af25082eed044683c68230166865152fbcd486d5aaf5fe4f7aeee9a803fd5a3e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he409e822e00c256383c57aeca74fa5124adef0609994d629a7e4753971cf52a12903f69150e89f87014db0cf92d518793262;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h453d0012249de55faae4a82f0c918fa3af6b4598758881c908edec7bb0441d77cae440d9feea25cdfdb2277ba19e783faeba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb40762f36d5e226823b305451b08f58d50812fe0b492bb970dbb22ea6bed715b5bd4b641273b019d8ff6211202678c9a3ba3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb208e118f7582d319977c582e21bf907137182eaeef95e9cc8744ea676f6e4b411f4f25a1739b893f1691f100f1fe5a8b99e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d4b4d6b5fe6ce37d4a7630fa39db3843cf53c231891225543e562d3ef30dfd25dbcf3410c9dfd9a5782ce5e3d021781154a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d584c07444685387f22ff31317d9b2d6672dcea3fab013e1df56cf1797fca6766dbb0dfd488b72fc2fbc8d09091f1e657d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac6c34e79ab8707d899af13368c38c9f3a59acaf3f3a3c8104b42f4dd9f6bf8391011618f68ed25c0261d8883787f4e7507d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f457a9673a6ddd2ec075ecfb86adc1fd237b6d3cea77e039de2c0adf953849805a796c0f43b8817020457dd6296e9b68f7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5934194aeb087065919a3e199d877717dfb4afd44d2574ccd9a9f061793b5c563d5cafc18569935ed0097e07d4cf6c9390e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83d8b3bcc14131158544e5f632685473607b71a79b52b8398966f244f1f545d827258e373453bbefc1f018dbc4c2ea300d55;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha279dae6bbff8a07805d63b69a7c62e5b9c4bc2836397ab9b58b8a1f45b235c7de61cd0304373b6dec77be74ce3a081dc7d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b8258efefc67feabdf048eb96c2c4481acde86fd36580e1e27cf0fd74c017e70b0a4deb21895716b58dd838cd3c104b355d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7235a1d2c5eeaebc12254e5ef49b3d94c292d2ac462274e1a2ded1fda9f405d679433598231cb8e1e5f000ceff2700c91169;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bb6f90b963e5695b1a1b7c17595e22c3f641dc46aa81982b5c319d677e8b899635552e972a87f08e788e8969dd0f84bcbbc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc77b8e8a7e09a054c25a2e6d64a99bfce77a262e319f006b90fec9fbca9e67387869592e7028df6b73385eec6703f34c2fee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2284e12ccc70435ef554e133c76871619db15e5b6a960154fb09678143d4d437bdaf207012d2264603004c162a45e20be5c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d21a09247dc00b48e4a6de2940aeea212828cb861ff10918715c03c1ac1313f523f7752ee672b0986a1db4bdb95f1060d9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ce8dcafb271b5fb35b3b03c1bba27f6486286c513530483ce8b8f35e9ccdf5ef66ae3f866c2edfc11fe95b41f3a36d110ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h652d3c448ef03ad9ed0552fd65202fb57681a4609cea6508367142064d61bf9500b10506382b86ee58daaede355b468ae9c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8cd71f212dc4a34b9d88a623ac3bfad521e02f5eb1fe897ec9864463810ecdc8ef1e452fa7221508b9c9735464ec86e81b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h484275a56ee11e8880f1267dba8e85b970c68e404bd795df6bfef669209fd1fd5b8d5f7f99e010e624d5f6c1489fff00c6ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70e0eb6791e525a4fd5142dfb6ab9cfe2bc6af640c28e962fc305d6f1259eaebb46945112b927f92ca07d6719774f68f7c90;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c46fa6681ebbf1b6b560170ae4fa6a8508dab970a04d73cb53c03900e5dfad8eab363bb79fd514c71ae88b223483e4989a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea13a3498cff33c86ed0aa5609889f1d23656b01ed7a49dcde04271162f8a61146d86df6ee4fd187b5a6a6ec93d95320f1ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62068f94e83b244c869eae24c218e70b98fa8e4c2dc45c971b12153965a12ef9a9c2272140603b54137a107c2811496fa735;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heebd71771dcb3e0ce2a616bf945863cd0db7747acd836510e6149d7adf31691fdb76bbbef5632d7eb17f69a90d34519e0b54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a08a6eee8af5dab22bd2cd660a5367a0c2950e9a80e42b65c3d915a1ce33a129ae665479720e0db890b84cb51b5257de0f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25ac822e5ecad499236e9d464f62944b01f2f92d680bd88fee83f9d26c6c0098dc94f225d2cc7809075421ed6a35f00453cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e960a6d21fe6b62c24a7e81e146f17b6a1183ca3c82c302e4baa6ae1d8b3124615ee5f0f22c9d82b815740377866685c79c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had2f5ec386aeea20378bc2fcfbe5007e245b944c8006e8420612eb63fb2de178d796b367dc049a3e9e856efc2df5f735ad42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29bbe6937b92311c4ba975f27600bb0581716c419805f814d7ea189ad4bee3de13bdd60eaeb201730752a25afd09739f4072;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5604241ce7ce62861e08f5cb8306d8d92ffd36100a1bac6279eeb5b52598a723fabfccd900bbe3a4ed45d3a608fedae91ca9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h791b8b5fc8868a8fa99659f73ccc5e2013364e33a078c3c5a34d718434f4b772cc42a20045e98e58fb424e6012682f4fbbfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f1d320ec25e120de1c963fdc163019207e2df40a557a5fcac3a02b18fe20233755ed1595adfa38d73e2d5f4c9cb63d1a2ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6f2ba236efff3bbb5fd2add73e14f2c60449848187dd0c9d1fd60dc0cfdbc1cf8fd7d3c5a0286e5f5b4b753cec66c97ac7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3b9d800b979a6e32ba64dafa4fe409a33a4bbc77a40310d8f4e040a6b8010fca40d468986ac9c433df045d80c45e7581302;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea4716036c44cbb6e8e61a0fec9805e99280e90cc3164e793cb4ef261999baa0d1a5f7ec6d02d9c3e60aa247180d57a3f17e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bbec6ca95ffddd01b6929005c3d62dfcd31240ba956748561bfaad62889d425633f93a310ab1a5d11dfa4f67e7afdd4baec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12889399a651b9c324e866469014aee255889864a6f1b8fcd6b86cf4ecd9d620dc2863d2063a59b5c4b002ad5be2b17c3a83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79b8638c4303f522d12e6bfb3e037ed84601cf131f742021b17e5104c72bc25618b5b4a8f361e8dfa33f4c1f391eac051f4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3857fc9283812ecd2982aec0b33d73a28ca432aa081f4751a7226815b4d0d93c67ee604abcbd1a675ba2ff7d60bb1a4ea5f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe611ab6c9ee44760e2021bd9c01bc93652a2e621d0606e1af8545cacabefd7be1b8256d1ade264f56ffe10db784ff94bd12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4c416e7b666f434b892cb1dc5670b4c95689d13c7175aba28d75f78d83ec25dbc877c016f2bde7986a95d28cc3f02ebccfe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb19756924187d7237c168d001ac1443eb07bfb217ad4e95058305595b1f33143617d3592d7a9f026c3829f2798d2818428f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdabf7e99bb81a8169aba15f80fbede4a7617ba4eeb57305743fa9b62ab2e118b583c55cbe266b1cbbcdf425f54a2887aa35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27275c8fd81dbaace8ae94f33bacc3ead9287c1be346f7b38123f2e7a4881dcb504d0f085978d92ae7f7983d67b13468da01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a27ecd5e8d94f9cb06269e5a038af48e27e36af9984f98895ae0066a6b2d88307a39df295924b1c11f13bd6b454ce510fdb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3888b9c63c2618b8ab4ef888e6b9f1e35ffe409f38f8198fc1ee2534386c870365d3d436d8e1b997272e50e316e16c10a7e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5061494db2c9e45b7b2078deb2adb8457c6636d422eef26d8c96c034afad72d8a45f79f4fecf2ce60c0153d213ae4d5d285e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd101a857ebdc67a857483679ba4acfde33fcd0562cecd71287b41fd8f9bd145ff0f889e97d097a70dd2f2c53016d48ac7bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h211a7a55d5c06b70e9b0e211f5a1ba27287667a1416b31e049682ec9649b0b0ac086b3ebaf1841a98580afd37480032f8f6d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc211d389f88cc539ea6ca5c5aacc4be65e8bd88eacee45bf7e8739c2719a34528de8f60c6064980544c50cf84a57ef9e78b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb0f9a47cd1c361a761ad9e1bf21246857fe29655edc745bcef54c45e66de7f2073a85ac01f7d0364cb8c0e7dccf4598cb0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a970623fd3969eca5b691e0e34227291e842d49d00be80bff21dca8bd486b36ae9f7c542355f891a720489abcc44c46778e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e52ccb5706bdab817991b7dd084ba620da6b2e88546c71ad20802b8d45a0d75938f2a6b1ed81213095e17eb65cb30a532a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81955b9b3edd19530cd0de17dc23c3acf5e917dcde88e530444ae9fb093ae748d4d9e94e82ae63250d4e716afdd97f88e3fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8722527f240e8ec4cb007395968098fd4dfe1d83fb62f4e729bb490b906a5118a24e2e45b6382a3573d61f6a6cfc19503f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7587d1aa8ccaf2926b9089a63b09e34629f7e83f0a5a43286aa174e4d3975d2fcd13337631c73b07572e6caba0202119972;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3938b8e18b6e808e4ff90cf56ecfb88c5c61d127659b542b7e208c7d176c02dbf0bda5bf6945753216dee2aba3852ac08f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fa9d683fada78055225a3d70a97edf2093d6f58b3e6ea82a5e9abe568d2cc7582a44c2389b84b7e558f5f33899166053f54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa770dc971df3c59281cbe3119e8224383783f3e94a903f8b53ff87d1830bff7d99ca27a612d152a241d0c9de639691cb18d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d54e59da3710bb36a6bb99a6b161a361e5bc83f5ffef4d6c6c52439bd8b81b7a0c204af08da48b5c5e03d5f66c9688b7401;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d2342124cb6874e2c875d80898948e35b5e62819e94c8a5eb754ec15168d8474462e5190461dd43beee3fafa05159710eec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67838ccda46dc23b09cabbc7e2810b3fcdefa75a3090e4f67ce475a699d9729626ab8ae851088e28171ce5c1fab18d704828;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b82d8ac3fb7f91a02a1504ed1238fb97664dad24a27e6570c09fc5fcfcf0d2cdb20cc79433bb1e29a9bbfed07c1c37c7ebe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa74c662e93d8463d7dc180cde456d0fa16a16c7f7cf54d5a20c79e93f48c1d602d3f70548f00a3947e331332c46518250ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5e457d2a92bac9eacc643cd61c3f674cb2eb9b626456583376328305ac7fd279d425764cb1a97f2cb8e9ce0e575b32520f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h893292a86c9e3ef09001e35d25eab6f8b364771ac668e7f9f3675413c6d59f43e80cc59c250a89cc4cd7f6b584043c9aba3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44524ff2d629c13368d41f2516a4946e986beb98b6eebc29945ba01f6319b4f55d95cfc99f8f3461f5c1c5de143bb093fa3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h760a3b69dc4edcd8be01d692eb1ce47a6648e63909b0bc34bfae2eec2385618a69294798777bfb008a63fe43ab30967ae099;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94a4c12216d70b0589f561d83a57704d2358e5e20f0d266cce7d10140f510dd21be871aeb2efd8022997209caf865cd89072;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf28088e9b98c786407140742c37f60f31d6aa880e3c05bc4c32d2424bd69c03511b7ee4e19a387fd5f8c5d69abf63a785564;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f0174f5e173d85c605e2e0d1ac486b3608db18d0ba20d8b81113fe59ef3b6601211049bbc5de80aa3d04ae6e30299882fc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf171bd921f6b446fdfe217bf3c0c8d525ceb919fdbf16d2d947bc5826da7f4fa2149f5fbd9d43445c995f919a59498f6492c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h382957d65faa8c7ecf694e5c515f47fae0f0259e0deb1e53c35e1f8e069c06ffe9badbb7089c16995172bf981b64b789e754;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe3d41d1e230540cdfa05086a637d4e2709db375c01a87c9c4bd7a8065390faf0aa7e2d9576f63f48e960d5529e57df85514;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6f4d40af2fc30b0dc8ac18371667bf996d4775b4dc1755c991c3eb779ee6c35122344fb9f583bb29a04e9d0bdbed2d5cdde;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e98312a11f40cd4bb433df9534125d861a6d56711b25b9833f53769e8c14b7a10eeabd9b71b3c2b08c7ca05bbb64d310581;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacea2fbb8305b0dae5af1a1f6ff1eed59b780b7db2537ba00a9360f8dc0138e61211c0e4451b9c2606fc95ce554532233895;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fb850e22b605f59b59b120a5735ecf5273c3433efa0075c7b909b08efb5549a51b884152e0be8603b803b81de50287297cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4635b8710624e909f390db45c9634eaa225ca3a96b97743d4598242ede2d82f03f926b3b33e2bbf2d49d10c242da0742204;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5c0e9c7f57309cbef73d22175ec84d6b5f4b2fd011444e235a7a422273e357b5879eae4fabf368a6fffa55133b35a62db3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd87ab45317c2fdf8d860b3946e4aa2522a55ff10a1e5f0b856ce34396986e20a252b6c6a29da638f135bfeef2a5b6b12854;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4800743514c14f624c44ab9648be58386906efef29cf32da08d08475601b65be51fc8a572b463245d69e0435f48acd466899;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd3772c2227b92edb264722040be7236fb74b669b47ac430827e911101ea6b2348ae55120e7f5950413a0b4e651177fe1a64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2db0d3cc9534dc11cf9c579b791be7fc80080b6c7993cc4b0cf4bfa828cb4ba9c77c23e20ce2dc8ee17085f433eb6ffb748;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8117ce142f06d3797fcdfb700a911bcb8a8930898a664c9c1678a01492b3d4a65479cfce0e9a896846038e65c0eedd23e897;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h986aa4f7d61dfab63fb064769fe49f89aae0211aaa9ef2bc99ced2249f5f1633353f6bdf706ebe41241d5ed15e5e57edda59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a9ac51c485b1c8587efb19e57f46a4bf4ad788a2c46ecf2497636ea61bd59e4b353d7c35f113de5d63e804d02b1832315ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa03660be8692e8d5b43b60b5d7245559e192831ef36937d1f30e38abc36a8c51c39324b9e0cac1b7b20ae773923e16a4a73;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea169a1394a05e5d091fc523eafe04e742b53ba8b6dd3ba41a13192a059500e73e1f4264b8883c542f4ffee5fb1f4963e609;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6a18cb713ec0e87858e7ac138b9d3ac4a25ee2429840df24f41f502ac702f52797ec6729b3a0461a643628c4779ce325ffa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8864092c6cab555b0a777638bcc6b9ca57e0cea92642df089f01feef9302a91f7272fc3335f87e659b4e197ecfb49ed44e32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84c96265875967d079e8675fa1b01b4c71f875cc1108d36d3c3164b01d765d3d4fbef199504a855bd7f6da10bb5b1b5f70f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37e83b62b120d45771fcca20746075a4735778ad43c5d79a14074a15d1313f420cf961b2b54508007a2b9cf9f6c2a81a919a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce0277cc7c0b9389186fc90169151f87c20886be12ea26f137761c34165268f9a3381b0acefcc17d060f888d7394cb5f11e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc101219c55cdb8303126efa66d39217e13e97d4138a1031b2dc59adc8f5670114dff6ddc26811a20b10f11783293b6ed922c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h811e6d5b2b17f13499e6e135d92b522c04985796cc03fa5eca4e5a656adc25de82fb13815cd6c4faf26a02acb9aa04c7e61b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a0457aff8991a54fd1582a4e303c15a0168ca761a7533820ebec7e07442798e47be59ce46985946c5d97aabdbc5951a2ff4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8a73bd91c38771c520656b107d265cfe2a304d3e03507d38a21d18e8d17f5f2239d08961c42807918046d652b208ba3f6ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h563ed704bfcbd8f4c43083e1c68035c1f4d0806cc1fd7b54e2e29e5c97de18c33215e2a581dc2b929d6541684d9af6155326;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heeb07daa26de3e67e478a2b3a82014e8e923cc4574b86f83c62641a954890f2d2c58d70d792e9a9cabaee7617f4cbd78ac6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38b9f3ac7a0615aef8c3c38b68ebc85493fe505a6d68f0104778b5bb179775114c94dffebdff0095dc4103213d01163b9dce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee26d4dbcc149631d2be1122608516036b4b09dbcd71c4f1bdd560f8195eaa473e2cfa7efad66b6ee4eb6610f6f06eae6a53;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd48570cd5e4c1916863812f3d315f679c2cd88c1481bb4a68030946882b38e0e04ba7a0cf6ec1dd2f2131846af3a4d130d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h693dffbee3b9a9273fc16a83d575ed1fbfa4f1215c6e51636c46f9c8b268188257dfdfaf9793d606ce446ae20dd7358e63e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc88ac1f8619f1be66f2012944796ba6392b30293b7930589d9b7c2ff44682eea3baf99d1f9cad53e935d979dd658d72ad610;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdb093b6a9874673565c735291ffdd314af0d8cf612cd409dfee96c5cb9ec63ad7d6ddd8f09c3c1c0fe85fbe6db1ec94ef50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3b586ed658d65b0d619881bf24f85cff4250b94c2257ccbbce8acd0257c79f1284ac869ab1aa969c1ee4decb4fc3205f984;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c52487bac3713757c055358a36f221ae97ef7b81d5932af5b22d5e2f29ccb9eebaec3c4535a7d73ca9d2d08a10f6646dfaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa9667cda865037f006a46735a9dc84fe0e7abb7b8adc2927f134a56d0f9481bfe01c3d6f5234456f7c9230bff80cbda5881;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19f874e0931f420d81146e38f3330d39bd5ec76e356cc5ff790394e680dc259f233076326d5b1d5310192b6dd44224c4f4b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef1a9dc8f923888577903e1deb5fa1ebdaaa775ce8a6b4c26ed3c6d6a55b4d88ab046646a1da084f7a403522b7a66208d70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62ed44aaf6160857f3dfb95ecb167330b63875639c919ceaf7a1bfb4e8816aebf01580dcdad1f3029113b4449728370dfce9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80d3547a84dfdefd566244280f6244ab67824edd763c30d629dea12579d69b732be453131be20e046bacff52cc7789d75144;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h290e0b1894687bf0c776e8a82f10012e10d44c71ebd2571a8af03df4cc8b4627da9a12bbdac1292d4f1859805a0009b1178;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55abb5485996f7e785e623acc899bb1e49575ff86e7480da5c059dc0754f32e4b8ebe63dc4b75db386f387a405cd5c601417;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h888e62b840803032caa3d0d24f03a3b12e52f981a6e77ff1194fa9c1ba5cabe3fbcedd6fa379eeead069f11697baf9ceca08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h778946cd822fbbf94bd851b76cc04b62dd0addc6927afc15b76947ec02ca11f9ade40019ce5bf5e2e5cd14bcfa904b2fef4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47ac008ac976cd5ceed9faea27d0bf8ff2bc6b4bd314c31ee7693240abb5bcc74cc70560cae742b702d83dcdae1f869a9998;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49a659bf06a5888bf0bf24945fac42f0b34b27623c42b29a3bcce8d5172ec3fe42aa3de1ebdfab810ec2188ee6c481094f66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b33ab610c67e687dbebec2d58677382382bbacd61a5f62974b0773bf699bcc437d19bebafdef446fa2db36a44276f13d59f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50a62f8698dd26932d3a4466b467e7e892101ed9620be91f303b0812cf4d3fa7d6e717479b1b79e726d0e75bd35f63c69cd4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc57278290202ab0140009aaa39126b8f92daf967fe836e0d3db83306be7c7002aba669cd8a1541be2e261893c882d98613a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8fab50ea6ae30352cbeaa4afc8d3a8befcf0180649d145dfbf2e61e4fbf82cddded76fe73a3e3f3d14e60ee89a1cfe1fecc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3d73bcdaa388d5f76a80dfe8b52d7adc96420b7b6fe3029d361013bf4e7b222ddcc464eb2d3f99c65764e38227baf714bdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd7934c92f5616f3658b38a2dc468901cdb167766dccb1b2186fc1810e545f99f09e6f2c7930fa633010089524fd33dd4df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha66525a85b22057e67ef843438278f44816311f7c04471d586b8d4c299c81ab215dc9527ec7a161fdddba8e3418a123b25e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62edc0a4e3bbcb608a8d66bb1f72910b1a1ffdc8ebe1096c84ad43b8fb4eac08a0dbeee8930b9391f1b28c88079667e3a249;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80f86fd05a04b6c27d97eba4711f9474b39a865ad2b643d5b9ea96e9203bb1e61c70d0081a68d4f05b87ed18034716455cbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he395cf9399095d6b83be8cc1c078f9cd788eb755d72b3ae3969e8cec2e3cf120046baedb6b8be87738c47c8e4572e7bb2c3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb5d1dba1b36148c453a3bf1f08bd3c6a6d62f1fa0f950d51a717e0fc7a327a86fcbb56fc018e5ff3189bca8e8b345146b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d9f9ea7345027091bb0c8d67f1f082bc1bfe3e401aea96c60310099077b4b5f18bce3770b84174dc50111dd146c7e79dfec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99c05146b75002d5dff650fd27065dcc3c14e8f87211aa50fa3bdb5ea90dac592decf76c4bffbba79d0d9131c39c69d0bec8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc54800baa1e8005628d0ae66dd289bc412ae3742beaaabfa854c32f8b2f7d9d630d751170ee8df51d4fa6adb699caf0596a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6c024e8cb2a2f632f8aabebeba1f78050dfc6667237ba29c645b23a1591fc80e41bc6eb3cf1b9be3540f006fd133be77b29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb01f9af21295214ee3bd2f9eecd6d7a935e9169afc0382168ff97fe0359ad9ffef0c630eb1382332e4d609109bbf95c9fa3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58aa22d8c85d8dccde9331dc12fac6719d5a3e727180f5c443114c3b1b234f59214fc14f3103ea7fd6db937a65f83415c714;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc10afee669bbad1daaf240502b62dd66d77232c45c8ab2be73366a4f779d0b7ce1668fe94db28bb1ab7ae44c713c625e14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6a12364c75f9fc6d035da14a9094f485c0b73d487d352211ffe421e0b79664b7a8a653d590003e3ab0eba7bf09171118168;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9717a0eaa9f88234222768524890b66bc21a78187fb297974233e17371124919821e5902720ee074673dc9fe75f5bf480f38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37e5a76e222f5258d5908ae176f15dcf8610885d56dbc6a0e2ec34fa0b151e01a7dbede8884aebe90c1bec9e8f97a49d47a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf876a7d2976a5abbf4efbc65efba98ee91200af3eaf9dbfccbbc0d155b262bda8f25c51fb1338824f10551e13ed323c2b180;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf243339e4545ee82a309f0a97e80a0763e59d06ef75307c6b2a3152ea93ce0bd7432774366c7b3ff32a64d19b30f405cf9b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f068244a35f4ebc6edf6acc2dc9dfe3cbdd8c0048ef9c8c0deb5e50a7e430b1073d9aecad19a64dbbf22159e31e35e1226d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e2b016427c968654524d4a4a7419eca60cd17d5af0132a4777214bae0113422d3b9abe34c28ec5ea414400a5855cb1e2395;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6399b53fe6a53a522b9e7906c7cf5418080975df0b4f8e90c3dc9ee275c0c968c5ef509b2c0179b0cdf6ff311481564dd92f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40af57373923952868f1d4a8c22a0131086771e9014b8e6ec15eec9da6c6e062a380a58939bc8f04b8b76a057a3cb85e7be2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59ed74cf0865a903b4baec228a98bb2686c8ebaa848b11f4ceb9e9f511ccafef582d2d94206dc242b6fdf8a398602b292ec4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h118f6de3750302c7520a349cd58ec6713d3fbeb6fbe7cd3e72eecd0218f172f907cd597d7ff1d45d0e03cb472dc9b55e64c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27063ac6aff358c52cb3582476ce28657a48b3318c581a382e7c858a23812bae090833c4eb95d1baa112616b5db22e0b2987;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2501edd002c6853f54bf3b1d57b6571c8d226234c1e610040706fe52f684a2982fa75f6b17afc1772548fab6af109858d19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ebb29b4e533d10ec50bfc6555dc851b32a996034116ec50fff41a24077d139fb72c93cb330b1b8bf03e6e813be3f37c52c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bf1d1dd2d9e5e6facebd2d6f7e7754f3d073e7a1ca561caeb7e15ac00b713cdbfe55fbff84dbac4a9ed31d20e9008f024e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67e3d15374ea9a6c06b91247a0d28ffe6d67f38ca35df78d5f7b2fdbe4f1f304a8cd0a0d52fbefddabb429b4ef25efb8dd97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2ae7b3bafcd11a4e479acf832ef54a2eed2b1b3420209ac4bc9deb949946bd1d83e4878e0589e9037ff17ec786b65ea56ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4698163fc18948af0b748a9f8e684e56d9f89c55c0917b3d09c69b14e583219a1f4820e8331d23b282ca9d20de544f786ee3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2c3cd447758beeac0e31df56bf1e265a1dc16f83549638c81092c4a0de687168ebec61084af2f9deb284560d4070f8899df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a719e1f31ad1b3bc344c6c4c9fac9a9152f9c7ad59699d9e5dae91fe5a3da2921be4ee9405c53acef6ef97556a97149ec11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75179e3209bcd56a3ebda0a325ef8634c915064adab053f1814d239a8e138a1d57068847c250e18c16d5953e07577b2ed299;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda49f01a61fe8f4f64468c7623da84acc0d626e3126b1decfc26c0fceabb9ad609b0f55df1d1574880561cbc20742988329e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab4f5e890bcc66a983636b37490bcaf4d0d6fcb313def303f26397d038eb3c53a5d97e4cb889d405dd7712f5321175d8e4ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd868050a7b1b072df5ebd59a1e363addc2f65dfd900c83e3168f7d7dcdb747ffd4f2a3e2a9b7f95ba714b095d643efa3340b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccbbf22001369b5b78b0f68998b2a4ebf53eaafcfc74f2745dcb2b53c904b268cc3d2a7dddbec97be2907bcf8875709dbbaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d00001ce35c2738430973cc6a1733a07a0b2426b9b393cd4137d785d22d52853b6534c460d155719fcde74791dbbe872aa1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbae46ff43bc0218cd55b7dd8e05b1a88194c6cc604d8be4833158f2fe46f0a0f9e83105bbbe3d44e1c2529503d8f93c33d4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf15227ba7280e70462a4d7b5f756d4079218c850958b4d5907f8edf96c57012c2fb99fb34bfb710c7dcdda93c1c48ddb26ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc61c31b573bfd5df17a059898302a754e771d972f736a502e596ec3598df53bbf8d963b8bfa712d5b1ab5b5986135fac227d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d3c29eb6584d72bf7287bfb8648bda894bc54b738b76f6f72e3a00f42b8dfedcf16cb7f35aa2dc887aebf916134c9c336e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d5fc9ef5f5761655b52af8cf1302e83c3cd8af956ce669a2114a4ad803f4d5edd1aa7afc7cf13b388340e63f0b6b5082652;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cf96d0cf950133b1e72310e4ae1b313a758ed55223de37b624678a11d4f4649caf919f1a95495c890e60522e763d812637a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae2a99d2c089840d73b421206fdef427e4eb3a13ea3e4579e34bb4fff84cb4fa6de166938d3d14f388daf7a75101577fd989;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd953076ec684293943e59b5c41ac5312ada118f8c18f3d44480329917d0b3a806a564534d2c822accbd5fe33a9a20a63e86f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3454f91527fe25623b49cc8be532778707bc819b61700d81aa691c093308ff419a991354040f85476f48b132e48fd6cc47b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf876afe02c440163e90a4373de62e439da9cf8af3f1a4847f9d5366b3db7716a31d78bdca3b3f55ed5c87ae31f6ad4df6f71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a985e9b4b8157873722094ac82eabbfec3b423f8e97f0fbed8985a8a8720cbbbea1d0a6afec2929d32f693f75504def599b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf190aa61bea0f6f78994c5261435aa81d4a2129c7e5c5b45fe22e9645492059bceed12ecdfbb28914fa6735b175cd8a97a28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba0d125a53611bcd6d2a71ca12fdc9d6beac5c4969468f8b1ef81b7d6cdf36387db388d2537bec4a35452e72ed008fac081a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18d16f6b2105d1723da216dab23b1bfe9d2972ac8bf87efe8eb637a13960544795386cad98793ffad582ccac036db55c466c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94c940e60d6c57d18276c660b322a20036829349292021311af6897529d214fd396e9fffd4db40bb4a8be45549ae92ce4084;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ad4e8cd6e6db60a840955b06cd6c7c9a9d4291767b58f528ac1aea2c6cd2b11fe451dbceb6ef92675e711c27f1fb466632d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd36f52b93b7bf50894d2fc0ae1165f45b8105c4c29a3262658d30668bf873a2d83d816d9a4b3a14ad3496ef041493491a2c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb49045f128f483236e0727e9216180c71a0ef42a6ce9423b4c38795c06b3d30ad55110a69c825c0b7276e53f9bf7f0809730;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73ba320c830d06c60629b6b992e9e2dc0adcf2f05232f60acc6d3a954597a083db0da267e32bc611de82edf6bc72e0f6ec43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f6aa0037fa6583d6dd157b84de1c0e7bcba3d06156de44a27e625a174a324bcb802afb10379c510bc027c3cb0a5a2c24ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda981bf14fbfb1572f37caacf557bf22b717fdb436f37c159a1800c7a72178c0155fc9851e2c6bc8cce4d58dfa32841ca692;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf88c4f68d9816c8f14ff50a941c6f088c56ca90cf5eddcf51f64790c0da1c7f85301ab2be4428e3d7d75c8e8a6cf0e0372d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23f26f93019ddab266a1cad5500d953dfd41950c36b4c30cfa6c0272a7ea9237f915276bf9caa6d91f209e0ce8721c8e5b9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaa9393a50c35c7add3c8552dd3d20bc0dd1cc8065e84f096f00922feacdf3ea59beea402827bf701aeb0b1ec00a39ff0348;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5e7c3688ffd465d57b781548f647665fcdb3692f2801da136f75d976731bb973907310b6b154722ba75eb2ae84378910d95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdb2e082853ec6943787d0ce9384b314707900b95eafc11f3942be7a02a28f661e6b116599f274b353b644067eea24cda94c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b8d780a9637ef37e972d877de86032885462bded65846540feb30c434b60dca99926dd3802f042812189e7483c74367553c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18299651fbfef7aa45873cf81d15c4ce71b15b11c98c0ab3155d15b44bd4b7751ebbbaca0c54a20b09b360ee7d769c01197;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44fb270302859fd0501ac34d0263bf6926a1c255ff845546f537ca2f883ed0bd7aa91bd2dc895844a9134b2eb5864457e87e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d5432717e2551a0680da9809472183ba9d8f51a6bcd747e24ce9544c76305971892ffd1d88a107c7554fde9672b0e89e358;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31ac189fc7f0e40c5b60108a270318e7794180da4d2686c1f5c4ebbb3d051cb64578d5c398c8e23517377eff1587d8f22552;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33bbc86b5182a948148ca6711130a3cd2f95652d633e89c88e353fd4b80d002ba3a4f5f617fbf83735ae782d966fae9c1406;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd337edbc3d17cfc58dee86481ad8f53b1e873f349943ef0a27ec1230700d3e3e333b73e08900ea387904ae8ed2e2cb6164c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8011d5e8927965efd3e7fa9f1098b730b15798cd2d2ff4931a19f5a32d99b79c3d70d8127b0c2ac083c79e6cd5114a68f313;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10bdeda10fb97a1d36619f408733444ab080f652ea1150dd514350010cc8442434ab48c5f6f5428a8b7e89d795325d46499d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h852c2ad85f54fb07caffce9c08d5cfc13f747ab3faf6623b64fa3f45daafaf291c1b3a5fae29ce3a55a3a12f91d1c8ee2df2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefd49ba1648b283657def819162f9a52d628bb83a36532f801214f092493fab39c93403eb4d6213adededf84be22d2053455;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h868e14d8a4a8d07061fc23259046a88f50a4da3d07cceaf59ec4a1d7d7a7c56e1386cf8f7b037aa9fb1af1fe42a299a1dac3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf79d4923fb25264a805cf0ca61d292004bbec2ad36ed45e40ad83db1227cdce7ae9f071a01502233a16ddf2f05a10a7d115e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b904b281850804ca2f8fce886034a837c6d6a92b77171957d70056d54cb8c0e3eb7ad33bf7df6b216978b71fd34160d5aab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b4ce3d08c231c4595063e50312d4c5c3d400653221d13247de0e0a6f3fc6db2bcf38bb76312b8a0735f3ab47890b3e43758;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc23c33bd012333076bd43429c942a7ed3b5aee31ca13e4524e06f12647bc94e3bd9d45d710852bc79a5ea43550eed893cd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0c145bf8dab9400c38547b2b90400adafb63671ed9b9ce692011da91488ff30e7501b187e73e264f727517ee11af77c752;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb13515054f16f2ca65ac3eba2efe11179b58cb9b49bf03b1f5cd8588fe613d5671a1ee0e688238c09110b949119b99d383c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd60846f5feb9ce948d5bc7b412331e0b15438130e232b41262febbabc2dc24048e8dc4fe010b5f3ad2d28ca36217fdd2b8ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a71b07d9fd239bdb59b96156d2052598ce3954a402263421ac69e3bd3738b1d8618cc381d545c2fcffcd832380dbb9a9011;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46af46d648276bccea114b4071052a17343b83d6cfc625954863a5e74be89588c63dacd4d7eb02f43f54e581f8254cd5b19e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h197e6c81fea22a9f043279f8ffd33fe56de152467518116ef65cbbb2f708f2286ab257f7d93efa98696e4e86f18ff5f12100;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a5fdaa3f5accaea5392ce0b40cda0a4291d808345f52e4dbbf0f83da194b4426045a8545a2d67dd8353dc70cbdf50439025;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4244151b6815b159809ead7c63610bfcb498ae0bcca4a1ee23686143144bb1ef5738f3d7925c43293c457899eef17b826635;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7648125e81b45142034053a2c2c7c14d5ea1fecc579ea97e934e3f2eb455e25311e421bf3c6f713a74a5ef6e224de58ce490;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfae822a1a24110ffd452d37c093af413c8efde9636efe6af50394d0b378e84e7d0b379a8f076ae896e8e60180f7ad4c552e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e0d230a16b5bcca345eb9afe7c4e85067a78f36b3038842a3a386263b92e2ef4576985eea680f0d88f8e6697b728f9d8e1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h385ab1d0383893581ec38e8b1c1629845597e6f7f3af244d726374b54576f216fd033ea3fc29e559b7c0af59f3f7a294e531;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2a15b6e37a2256449657825b079576240a08aeb8108af02d3bb94c49925ac61e2254203ca5ae5a3320b7b77cc62ab080ea2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9436844b660d043f849e16a32d498af70950d01810f28ad359497cf9a7227fa003559655a59fc1e3881bb7631d4ef7dfd8e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9afe6a39e789a2df2a4c3ff86c69c2069df09cb92eae5256da2166f4b55b2233d935de10de3f5a6588b13c5863169b22b84;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb9a5d4cff290abacb9e5eef38a9599f07cd68f097025a63972e08042d5d70dec128e6dc540d008d7e8c58440ec14a33207a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h253a5aed26ff452b960c31ae591d882b54e05dd9406eeec54a9afecd6021368646f6a202f2da0f66cebdd8809f92712343ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8980dd6e8545eddec9208dbc7873747cb3c34481c474b37440d69a43bc8b7450611cc89999639c6d084ff47cd5aeee2e1cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7b3dc6041cec7da8df736b760f50ad706610b373f312ad1d4fcf8c52b2265d1ca6202fe67deb29d0956bf41feeffedb3318;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39881f1778c444a79e949fd2b8d56a87586224d8ed0a13586ffafa431f0bb56b6cc0cc5eccfcb87dabbbd4195ef4df88250a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34abfe5b508c7e53abb3150f0e8859b4118000ee809d480bb1663d8b5a02123ee9ad0ba5a0bb3be0a1551821e57ad0cc0ce3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10a0b3741f635755a079ab6181a0f5daa33b4927d59880f8073bb3ee8123d10e59b90bb39d4d0fa2c524ce0227b9ef312220;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffd12ecea3f9fc8709a481be12ad5df07560ab260eaf82be15396e854ab07631105b254380fcd7f237fd7eade1addf3e8732;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7f443dd6e699777f82140406eb18dca678fd958f473de6e6ccb30dc7fe3076a9462ca322d438d04b7f03dd0cffb7a82348c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4987520b44570d6935a67528635aa07f655c505a85e281b292c79dec90f11f0025786af89f69cad4ac5a3804e854c64a2e94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b32a088597a8ac2b17977f3e3c8da411a92500af95875feff398664674723a5591234b8f924bde8ebe2ec78d33d30aebf6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ca054ef26d611fbd018a159c7c5e710ce07f1c42a81e414f1154137ff6555978d5a91646c4b831f6902b6d04b854953d128;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0d1e34a43fb8514e2010316c1201598fe3b29cb152397727c5a95f78b8a3ad76051b9934ce809d95ab4d1ee08402d591836;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5fe4c8de7746fe7e924aa58f76bdcc526647d5135e468cf0e4d264a55f8847711841a701a31b063d968e0ace62e10208acf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18e6ea3f7b3e74b87c9e6e247cec2ab8b883e01754c10cb884e4bcd58364e4495c9c5c10ebfbb1613c77ea268e2c8f5f4b02;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9d5941926af0a92491ad6a6e0cf2df839114bff22bc38c1d26a12eef99b6f945fdf11ffa9fb1d00732cf4bae1adf33e16b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heeb1d7d2d87ea054f1d0347d0e483070970b90d2f9244b82248f1cfb19ae9a2c1c5d2aa6961be5d717a8759c057f857f82de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha186af159cac80ee3654a01bc59bf78833622c7ee62cffa18be40c592683ec03caf13d53606d43053750e5d02f20892f4115;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92913f7bc713ff03aae5cb19b1ee5b54af955d2c1ecaef8799543abf1ad9ea33e683f4c2712b1039e7c060548c8c49a2a38e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7d24efa9270bd41b515b56b14200d5e53a874f8e2b8dee36979c35de9da1deebedc413f4b9908e7d94400778972781edda5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bd611f5c567e03f022344e81e0024485c15e1eaa4e32669429eae188be8501aaef6b458b394292a574604469a5cfd6efb9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h507501dedf3c573d158395d8a58e852fbf36c6ee478c1d6ea8971a8bf64d09e6937c45dc50e9321fa7e1355230da86336d73;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f2a9c868f4e17e70284f4699fd5894cfa4ce6ccc61020e4f4e0943f60115c7846b4cbc0dade96fa0bbb6f92719b2087d54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd51da841b144fce52baf4f181e46d85fae089bf19d1aed9bf76ac0b72530f513bf7ffa3d562c13b0b3b8ef9fbcf8554488f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6d4a1d3df0317d6b9bb8ed5e6834a2e4581d7fcc29e79e75cbea8741345468e5b80a4626e15f612ee7b372ccf810e0cdeff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5395c6eb1e068e6fb33d4339ffd37307df8c602f371d61430c8b84df28b63473a4fc8680bf7633a7f8762c249a0d4f7fd01b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51f53ca0145e6026b56212ac6f7e01aeb53cbc649ee9930db822578e4468170b337deb5e4a864a244f6ad48fe70bbfe84076;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h608ec7b76ca09946082b972e50cef28ed5566ffa2885387d40647b37ef2fa07a13c92a0ec71e625473a245d84644080c6255;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h976e4ad58f1b8511952a6ec9bec819d0849bffd0bf1c0b0b3b2d7daf6fefa546bc47eb6a3a7bd5ec86b7bc7f189ed574f7a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d92fe165b6f7c7f78c745b281b55e0bc1ed339c3ff3dae95bdc803eca051323227b1f7eac30a7fc37f464ac61a85645e6c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43edea89f3d8905b6484afffbd3c96fac1a76cfc81c5133bccf5a1c9d65b00659db37aea432bc039d5b15b8d61028490c91d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffe8ebe40fc8e0771c2b70f15db0cf8036a28b1f7209eb505cb4be07c70112e798bcc40e88c414517fd185e19cd66276df28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha796f5660da8dab90d95829b6a4b3f5e0343c2aaa2ba763096110b5b5287833439d2e06e3cc9a5807c7357c4185e1e23e088;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfba745da3ce662ebb4f4088affc7eb9846fd5a8381efba0236598bddfbf3568720ba9a8fb05f36adb9ec4f6ea70b5a06a5e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f68a26792eb2863e9b375cc2f2597e1f0f3d48925e3173a082a56177b94298fee0a9be65e13c9c3009083d4d4e972d43203;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6375cf31d9608e4a00897f48284a04ee4ebe5c6d2eebb67629a25585916453ede6d971130aee96e9cc71191d60aa4b43f774;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89a4d12b82f2d54a9378962cbd08acdca6c0511db1208343ca66402c75582bc0c609758a59deca0ae71acb889790ea29c48a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0ebb303275d176d173f881430f71b5b827fda0d8ff6bcfd4cc39beefe3ef037d4a4ba5ad4842882322f4f8bf6284a1c910f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba2a0b685070eeaaa7cec816896bad4e6b4f8d2742cb3d26df555d90603f8ecbef62dc82a988e1e0fcc8c6b7dccaff358a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64fc4c0be2d26d2db4f4245a01d727400d94caa9975709a74d0bc1c9266523bbc8484a7beb0c6472d6f379225e2ef38732e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cad704ff6eca2f29dc1cc3f7346f692a69c0bd62bc69b1a772bbe56d1f612eee07a7dc2841959bd22ffa8e5b2d865eb63c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc57ea816bb9fb26e0f1406c0cb93a0a373e2b70dbfd14042281afbfe97a270506ca520befbafb6a4bdb67e03a4788bb7a30a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcc3dc6ac0a49dc64495a1a8cd26b1533a899d11585dbbff94a4bcb86e0bfb13b0a726599aa9899a1d30b7a0cdba16102321;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62608638b4ae2f1fc30750bc63fd7f83db4b8e06237a14c48387d61b804b5004eca6a490e67b7d77da40b3d8250137814938;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4847328dc1afae254304e14aae4865fae9cdc5a6d7d9d77b3c3823ec5e8373bcde614dcef3509dda92135e4b7de8181a787;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h897972fa9b7806fe8e84e7f3889e3ec48027ac1c1d2f92de356c628347ea5376fe8ec572a5071d9a61c872c7f790b6d798ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7244932097e8f0b4a38a5d9f1f399ce1f68c0f3453c2433eb176bc2f4079d7a41338c24cee9c797c8c31eaa25109e6b16647;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12bd4467632e57692da19156e9dcb0e3657b11fca53231a1f560a8ca0079ef89fecd18823979deaa68744d2378310425aa05;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29eb8ad98edc6c0e99145358c2bef5d594adcd3b2e5775a313012fb2bdf47dde40276161eb7bc28cb0abb613f1f483b3123e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebc472b32bc709c117042340ac5516fde20b3e99d35d6921dc2bcfe7283ce9a7d0ec8aedf9ace0167c5be87c3e0b4e6bfe95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26e2b12edbb66b857063c9ad3425001a1ff30da96bf5536594a26e9b09fe886d45768eee4e595f5dc964ba3827ffd49dc8e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h871ba6929212844c07236ce5b0638faaa795a7bdb80ac0edcccda6dfb31125264882f9ffef6a0689d4c7e6c6a1c18e1b59b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3949067b3458cd4da338eb90f098dc4751543bc9a64015f6ed3a88512cf2093b244c081eb6f6f2d4ee0814178cd33d739aa8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac2b3b32a2f422db8f915dbb07fc393a6608b41e906a33681d368b05d3c8ea909dc819cc1bbd2c99d41b3f43f29294ba4851;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h555f200b8009c876f102a0e9afcdcf8b20cdd2e83caf7af43d08e86a823b2dc78c67b728b5620bfefd70590840a1ff0a63e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c2b157d88417864c682a706721f0f11b47cdf356d444961c165a81ccaed32791ea3c91090bb6339278bd0fbeb0a854c1778;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h343305a2ae69ec012f5e9980e864adc31dd1ecaca65123dceef31f12108df55c04fa6b7cdccad4edc3eb4fb636687f5f4bb9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97016143dd0f28b1db6ec7ecaa79576be5d6e91729d09dc1f580826c385c466b497d686da3a8709a7aa1d413903bde20c4fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h996f6904207f21685cfa5dcee9a838d9b18c333a7e7f17c89bcf360ca5e1a11c170d25f8f15514a709568dc3512d8a9b3186;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf1e48cbb3f9f14d32679cef41a24628a0ce265ac6ce83fb16fe6b74af00edcb63b02e3308c46a2f626cf9e770da9353d61b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aa94c12c23a504556112894058d039ece7bce3414fc42419b72fa47382e5d4cdf46c79a9d5a23ed452a843d62c6f66e3c72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d7abc12ea96e497ca4ee0e56c7cdb395bad64be3bc5a99fcbd60792fb3717daa8bd2574fe319b11d461887567e63c8f6495;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee2b777e696f499e83dea3b95ae9e6c0c96b95841833eea2d46b0b1f1bc26364ba2bebcf38619863ce3c6250ab849d5e5d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac1486ffee8dcc25802b423052f901d5dd33f2d6beb857ee92aeeee105d8657880cf3b4375334f6f643db63cce575928481f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fd783d7697a4885154563e4fb56e1f99e9280784caa09f9e2d69d57a14584d9a3deb32b71928ac75fcdc3ec87fa63d56dcf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfa353f869624064d75d61f4e5de5e4a997cf893ddf5e7a51879aab040bf6dcef8837c311ab16da7ad9060eb4f7942ef4d36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc25e5cfa5bdda100b1797ae0cac066cc5575707a79785214ca3cbffa46ab34eb5c5dcd7f6375b0302179439afbcdb04d2ab7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32c5268fa9c0e4eedb40e6e396248bb78c279f1cd2ef81c8a557b9f08614fa046dd549040b44df23ae90d99b8b047afaf4aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e1a847ced19cd495aa9e2264b3eacfba46469658a2a93b6313785db2185b2399dc39fcb7f4ca527867a6aac78be39141c08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f5291f9789610a866691ba45598d8089b24e93fb108a1bd866293599ba42663e1a0e2ee2d729e6cea5c636b87d76f4d3559;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb33f311c468172838119b348a5aed6747fde4dfcee30b9a21265686a19f3c03b9a74368805b7c62e9f37ec7008fda0001d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437f4edbfb19492b29356c3ac67f7bbc272992f11a7b4d60a1121512b926c5dc9f9bcd1661f6b524f58de9c3849568e28836;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h101d5645be36259c955e08e5a859fbf489d2f9582aeb7e4f776a92b67b392c7cc27571c41e1ee62bc63ddddaf9c228c57a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea62a88efe5d7b4429c8d8406ccdc668186ff89eeb183e18a2ecf0e7c8cd3982724417ab32439bb8bf3cd5fedbb4b9a60e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h694acc3bf6f5f807147b632e209175cbbe9a74484a395eae4aab61dfd03dcedb9c55aea4d05238d1b8589f90ce4ced325de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7825acb05d07eb32e8ea820eee048791cfe9f8bd18c880a86e90f6ed177a4626c29ac718b59458f2a66d4a199594074b64cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h527b3e7f682ad2fd3814bbb5bbb8ed6f55313e211a6a6924445ca4aa243a49af57ba9f49a62bd64b27db209cfa2addeb178a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9038ae2826bbccda7fddec9c1a9e49bbfe3503701b5d6c194f2c4402c55ff1d6283161cf56ae04ae856075884a7c62efbeae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec7b37ffd4a2df58e85cd145f7eb63d5f07be0bd5b2436bd28fff961f5f64ac031e64ef3e6a3bff43ceda119c0fbf4670ce0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ee38cfeee58b8eed5bba7bff1465970acddeef68cfa9771847e9c1f95676649c1371e51ffc376d90da3feea2348a7941dee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdc862af8b68bf97e1c634ac4a5b83f0a7041df8d5a928ad197d53808a7b014a30c4f939ae09bd7e8681f41ca1601114cc6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e55a8da74e71bd5d09d5643c904bb374ce1b3347a54711a351d750484827d04807bf6ab2473a5a793d4597a68e9e3a8c7f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb37c3756e5ddde192f70d91be0eaf83de4eef0d19b3bd908005323bc2df4c04581cb05217aa484ce2fffcab76ca705cb0a60;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f3979f19ae7080cec6f105c310adecde091f2c9c0d2d7e32af02cabe827b267711806964ba25654905ef6cf9276c9f2e58b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bfed2dc6ff629491f80f5a595fa220fb071a1c5bd5b47926f5328b3f218a380b8cbf63f2494b06767b991b7ec280ea59e86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb312f6786547e8dd87afad5faf0dd883a79af6d20faa76bd5c1655e0ac364db00c1c87ae9474f108321e6f4f14361fb627ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4e345423da9143691275281d13a768f81b958dfb55fc2b063f8c0738d033f6740a92b3522d40d91195c35e31a7ebb86c6f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b6afc0ca11b04d681d14569aca0f500c30b1c8b124a563bf7796dff34ee20808dacdebec3b25da92995899f859587bff1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a862185a2bf462cb51cac215132db0a30a29d6330baa785059ce1f5e40b98368ca0668664685bebf49c6146bb2d6feb694;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6966226db035e5c361b72b05ffd34d1176e61cb9089f21546499ff828bbc1e793b3d3259e981eb49da782154b8841b12571b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9ebb966fb0753cc14b3b3b8d8cb4f93107ae7506a571fd343448ee87c99fe2f6d6a819394faf4685cbf18c5843cf634eb88;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a82a9578d0b154dd9541628c8fbe9e60075a6829d4df9cc750aadf90d3852fb50aca9a215d6860f25133b7a8f1bf19805f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62765611176483eca82c81fbf51d7f161ccca240c54e48104b199454e79212f8bb2958d9dc5382306b692d43674db8754b0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4036a2a20ed61d12fe8ff796614a917114bd1acc7e5e03970523bb2638733c01696586bc3782499468f5b836590774fb69fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde25fcaf886960afa0376a26ef5fb5178aafe10d601b56ffb517b440c44a1a41ff237e98c64cd8a39976797a4369d1f62db3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6b389e20166587961cd267d6a98c6acf4a586aa7c25757c8e4d72ccd7fec4e9d97fba9196ef6aa9aca0b58a31fd08cd1fc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2241631a6d002796649c6a74f3d4cbcec676f579c8dc0b09a6d1c690ba0cb041c220d1d0d20d29ca3b473c1bb919904df3e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd008b2ae0163f75c89aaabf479a42aceb3130bfa3586bf618433ffaa4ba7cc582e8160e243221a00c1cb2c8482fb4a68bca1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fbdcc0e858926f2dcf3264efd43ca5225ed5d78b9ae5ee73f293110d7e9fe83894b053d6afa9e3a0bc0065d77121d776593;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc33e82d36b2437cd143af031d72cc929def1ab7f0b9fe0c750cb32141e5a6bed4ad97ef93ee69dd7e5628d62a72300facc9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3506ef99dfb77a5bf09b4ccf65f8b0caf443900d4031b948611b2ce3d8680a557f2bf856e1398d9e5a2d3f4ce751129f11d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52511e0f0d022fd7d30b609dfb42d1c0aec7288f019a69355ccb1d61505df51b3845fb3b7c9cfa51a90533e77eee3c0f4951;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaf1bcf54f17124256ea89c7d09fe18cafe655fe8ae53dd0df88117021519c5e532b634d2767b6af37ce9f18ac8c14cf38c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b8e5ad67700065c47f20ad67503e0da60eecbc12b821154140acd7b890299459aff04edba16d118d0ea7805efd30033c715;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58526e41a97c278b6dfe0b1696ec4a1723c41ed53d8af8c05f4228eb5877fe9fa51274a6bc86a22b1e2ddef754ef20dd8ceb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h648ffd6984349f4160b9efa9c7f5e663f4764826f5f27dc85df618610e3494c771add389c62e95edcfe327d48b33bc64b6fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0284274805b4db573f76fb37627452df0f2dbc904a7fcb03c90116fbbc8012405fa0bf59c3e33c91708fc8aa56ad8bdea13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f5d845586540857d39d53e5f91ef9351b47b6ccba308d08971fb859090430388887874ac7bf420d85e4d113c61e95ce0dd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h279bdceb23b02917729bc91cf65d671e6d7f4eefec62c7cd685a7b93f7f194ffa105a8abaaa44f4deaccc9bfb34133fa3fc0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6d3d1d501df5644b1a57db44ef6fe2cd09b4317cb06a8c102204c983341c6a8333c9304947c2ba4507ce399d46ec31950fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39377423e9f6c59cdeafb4b78c8aa122d61c177de80b46fb95911343c232d68881e03b94cd099f37edf3b061039bbffd6ab1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a7b4581a5808cd060eded6100552186b14e6ca86c66ade04bf916b337e4e5b3c0fea86da90cedecb5d838ba21a50dd45688;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48be40118370b84ad8105c7819d44f5a1642e8f754cbd4a1c219a735f70cc5a0417de30ff712c00b66d2f0cffe6496ecd9fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b49b12be57d5af69c6f809389bd004930f42d1cee1eac450f57a453cc51351d8a0a0b43c3516f22e3f5632511a0eef3abf8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9728bac5e7e12481f5ae0250042596770589bb7ceaddcc2c6963e5613430a4e803ebc0d794f66018d0ac6fdd238f7e61c221;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9044f25e99c698cecd208723d537d87076788a2bdebdc31bb750309a3e8e9cc67bc0b00ff09f0f4646de0ebfbbdd19bc2da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h674ae6670243a1c32fb90f2d5b3decb30de16418be3f0843b7d80d3788e754d6a88c3355ba1dfc332f8807c35b28a37de1bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7613e6a59954c7883c73871648e0eaf004f32cf5f97c8d9bb5d4af3311ea2ca0529e5a88d7a87931a52face1746d78c9ec0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5acd51f524d1bdfd99a4b505f9a48d8a874fa8c065d2a6d4f2909e88100c7ebd6fc7eadf2ed970153d8b650ecab17ee51a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb40e55a9320a9360d192d766e9a3ad35b22dbf54bdc73af290de06cced16a51b2bc870ee13e9402b06bb7cea86830d211783;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13d39a040128e57b0235c12272db99765586140680941586bdd322f26b73b92ab01596039d45e3e25945767cff704d9bba58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57412f203b62926d264c11c02d27e1a5a990a85f3d8c5dc9986fd6aaa2bfd23b824726dc71eb4d0409c47df16978cac15029;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fa1f7b0d968f7effe85f1f3ac596e794d0db1598603b9086abf3370ab9ee0e4475bd375687fca53e585c8892234c21e72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ec2190106aac0e4b589de648dd314806bc68d6dd5ff05ec7400c0dbb1ad97b716527e11ecf699787fabca6dfd1c97badfa0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c28829edd5f591dc07d15ad33b8d15732d35d65cb7d516bbe0f5afbd127224ccaac005ab778fbdd10ae457a297754e7323c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b52f3e549b1a79379e8a4825e6cc1a49e53996fea18c7f8a420b268d25c3d35ae281c2d68b0789ab193da1257897d29297;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2536cf70c346a3cc36aa81f61e71639aa751d719bd1b23c41fdd77ce2e54cc66be542c7c45026f25d8a387500a7032b9b3f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc54d274d0e8eac6666da2bc96e5b23fb186bb3ec2ed18307df3eebd55c5564cb2805618c0e267a0d432818ae746268c36166;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h312504f5b59239d1b0764324ade18bf6ed40035a3921a59c42b78961ef9cd2f97d61d204597ac9936f7b4d2585f3f521ba16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9912605e41e41a723736534bfd1d656c39417c77518c810c5b6920c64f6533a2c0f81fdbf4a3464f6dda4ad77e0f9399e539;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2512b22f5d9acb1829280b09782a4be1cf99be17f64433154e7872930512329e4ff203dbbf944ca50c46399d5ca7f8e3b3d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h886f43b3aabc2ac6c318894cb4162be8e0534073d5ba1bcf4d3ad9041bdfd6f04e03ed926ac301027557504f48421b892999;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d7578a4c00b12b67a4b7730e92bda1ad4256a1e4d9e830c6258bf884249230d121406a00f1dcd5510571db2f77d420948ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6089edaa4fc594f626cc8c8d95b4aecbce288bcc20313babe91de65210f4272eb4187785831d6a14d51d2e5ff1cd442261bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f2972fec70aa71c2dd1b14ec6ee6f7d9d7005058b162a8c665b067495aec2c6ca462f5718b20e4bc12559b68dcf4d2a629f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h207280df80b75ea81f2ccdb8afdc67fbf5eb1d2fe1e5d724e282dffbb8a21ca7c12fb38b890ac630d053afa42af188738482;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffd01fbcb4b845c32b1fcc827cabfca2f8bd90a2d9653191e942bbee7747fef6d41b26a7d3f310b0dc18cf42f9b550c9a11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a380a5f46f46616de7ddb06bc4c6fcbe171feb42cc1feca977a17028cb5430520645ab26dbd272ab58407a1085cbec351d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc77d475e07fb150456bd4e923728b973212ba29ae6a10076e17d86e4f38ba4e941574ac429dfd80af0c1e82c687261a52dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23718c644375eb99f13474b943c5fb3b27f2f6e80cce8ef009cc9112a3b97a95b1009c4a3dd49035490d7faf8e5f18ff5fc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7753ef97308ea14d9b86104022af4d7fdd6696d0212fde85d2b220488e3107fad2a590e03aa8694845babc1ee192ce8c2cd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc07d1eda5179b44c0c2cef35e7c7e7e5ad531e0205e67f3172f1994b9ec394e1c157693c3f71fe90515859f363767751c7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd59598151f44e89a5bd966a6b5c2e1d99fd72100ac832743d2259dbf7e80a45c08c9f3d34bf02bdb2137517c89a77dcca95a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf13072ea113143f6a8abe0320fe66ee71864937c242f59f3e4809444d448c9e23df7f5dbd3796a697e3675f7d0a6db87de37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd38b408ae980d11876e70b5e2c1a6bf7c6164c946d885fb60d4a46dec1aca68d5f50d21ad5765bfc5e83a34612460ee5a53f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57149cd974bd1028e3f6245c52a82cfdd9e5dc5d7dd609e7e0c18f36b3b9de652c715e2f529ed192589d3c5e91cab8c340b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d00ad488b7fd37fd878eddbc4a9fcab5149ff3ea21822c9aa3d3c8b832a67ad19562d033098c431586bd6f4d80b9112e99e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92ced38d1b016ea73f4d91ad67155845a4b13cb2794a865cfb387732f519635f4494c2b312145290cbf83be5fef3f22e32a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha52b6dcf4f31850880d5c8894fd2debbdd652359316415a2740e62613581370be59c14874f20fbeba270ec985afdf482c275;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba07445304d895d09d75e68a755ee662c6712d174d35630ef5764f4f83c42fb016558580932e88fa822350ca29e13aaa17f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7301dc4f5da3d5c46c9d600603b7d5fdf56a8c5fbcf0bebc99436df4269d89416aaf7f1ec0029b3196af99870dc81d0e4a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bbba33c3ed68bc8e937a98fefc3d8e3cce4825a2cd969589e55c68fe42c51bfe28ba07d69074f7c33d65bedc2056985022a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fc61fdb2a3ce57b2449f5a4523ecc1e82a9ec75d3ecbff2bb08ec6c1fd7b03c4af63e34983f94df13fdb0c1076b91c8dfc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc16c7eb3687cf2ceb3b60afdc1a158d1285284e20d18ee228e08fd9d3a688efc1c372c38bb6409232989adf28c5be0c413ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h121bf0e843d46a541c5ff6d3ac11c48adc79372bf69922680d144c51e86b72770e8c5c2883d1e40751e1db2a381ae368e2ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c5fbd432d6820957ac36504ae3cd31f56cd48f93a0ee1ac84ce707235dfce342b748b4de1d1b95187a860f632a1a7ed1b7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9609a69c9a06eb21ae987cbac72d880acf8fd0fe4a8537967fd99e7934b6f68cf6576fd17bf1bb07b70fe6983e7944e68ea4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52fc879299ee76c684d1061bbea6b94f92f82a0426f8e659224c30e50f901e30f1fbc00dfa633475b1b5c01c472885fbaef3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h577a8a46064846045e0e8d9382594026f30ed407bc7bf98c990235f30cd81443a9436f2b4385d143bf185119dabda9631419;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cd86969e8561630688499f662746bbf202bb59563125482ab993bd7a27c5ec31377d4b56be4f6d9df422a15b7883de9772e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cd6e5f015edf052ac08f0cac8f2cf3aa264d83551a17f1f55f8f1a829776fdeafa66aa2dba4a316bfe9f70385c798957de8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3ba86ed7b90ca7f673972cdbd13d5caf453194c4edde77c955ee12f3bc48bb9d137ce8b9efb0395a06e5715918ea2c9d4fe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6728735848ad5363c417cfdec7c89a395751395546ecfd19f40bb66e5fd5130983a04a72481ef4400e51e627e34fdcc935ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a2c6802547d8872896b45223003c3b9f5d21b9cee653eb76f0c49cd12165f52023b1a4fdad0c713d0a4933224cc565b3ef2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1746280b3987ba98a64679384020a298d109f11dcf16f43bb788e7d6812d9885680b8a6d3c8c5a228c5ef53899c6f60df879;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10b8bd35e9ec06290a88c939a1cdcfaf44951b9a6fdc77684193a5b5e73b62c8c0c2c730b8f10b6b24d8fc1b5036b0f1e5c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6b80de41709aab3c2dc7958cf255e6412d8e57323b3a7117d7256e66d0c12a8c3a32c28e332ba357de5a6bb0e35d59140ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ab580149c141131c9acf1113200a7fb99aa47c2443056b58d548bb303968d38d679e29c8634392d206524dad06d6b710c1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a7e75a41a2d39518799fe4bc90bb6bdd448e8d7120dff88199a0d18b02c0367fe39962a0e859767625ec7aa9078b4b8d174;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47047f903eadf73e81b1e4f8b6e8065394a794ce8f0ef52e5779f6f068c8dc7c2a98a7e7520e6dbe4cd3bbc115cf4922650e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8964e65ad4ec849428017553bcd6ae2c141ce2236c182f4aadc43f7d94b8e35d61e9267b87ab861a5cea4a55f0baed58eb8a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h191347177a0dc430b0e5b36ff903067b1be1d3eea4913127844c706f6ab4e5f92a258e17d51cf415d6667b73192543ab57e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e7427213ed785c5572317662a160688152f6e92b6dc48e53317bf23de5fda8309fd6ad9ba0e916aefcf1a817baa0e37223b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8b6a9bd68ed90dd258932fbf9ed851fc6017f13e97183bde8d43233d05812d31c02015177223ec8223cfcd877d7e0196834;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0a95e97c64a49c11e9445a95282b71919be9a77f5eb5a85ecf16766354c53a6736d9e5bcf79d0bb08d172c965680c51fb1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66876d841ef083d245246827dca75877e2e5b617e3b787e3b73934de45e20b28355dd21ac619230aae3a25e92398937a55eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca221635c13a7b7c29de194df155f9e0e445d929a82a7a71f5d6d234a4d73a469f8f8bc25ed3312995339a5e3242ec0005c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h542832d24e40f7b6d8ac456db09e997a52994146fb43843fdaacde25599d4b0c25c0ac0c40ad058821de026a135089fc3fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h658e73e617907f47e957a6415939a39482c39ad1cb30d6390bdd6cc052eb0e9fc965286f3065517db4878eee77f9f0cc165b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcbf86ce94586630004b70163f8fa6933e884476cc409e22b7808a9d7daa96b8bf238f7d57718462b9e8866ec3939cc33ef2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ed483d127e4c1fe3981edb093bdb92c55c0e4de4a8b86235e0eeb41f38f82543226a26b597102ba9dc59481336763103962;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb4ba9e4f5f4cfc930755c914e0209451f59e95015dec3a6aff300d8c64e3ab51ffc907e81c072d6aab2037baf147338eede;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3fcb92a7abe8d0ec3e423c8e7a74dd05133b08fc6cb2459093caae9a3736273a634ab282af604becab59cbdbaf56066af6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h737c6538b109303496533eb9f683c503294804a35dba919ede81d8009b059c801e6469341d1f573a97c04cf079eb890cc638;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c4bcc9a3039d36f04494fea92ed8b076f365a22a69727f8000215aa585e027dbbfd70006150c4e63b4f5c6c3239c5baf106;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79ce27945d3f3acc07325eff060addefabe01a3f61c827dcc6bd31952f7db3c5b77e28a698845879d6bfe93f084071687c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8262afa08b45f03e716f8668793a31b97c4eafc5f837baa5c994cfce61bf603c1d2a5874bdbc0602e317b4102cb8d7389fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36cb73194edbb1d9758a710d559c90a2a8a1904cb4fbe299b5d3cb19fa8b3d017339ccd56d62a97537cd0682b1c3312e0ab9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23cda98a2221696659aa60dd284e2cf0977ec0e9ef8adadd5cbb1baa690ea2352ea8ea5021534c7ecf8979f152bd414082ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h707f059b19f1a673bb2199dc39656f707b42fa7edc567b5c68805566305941ae9a324916ab261827dcc70009d68a8a950f62;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b865ed8d3fadfb630843b12261fa23902a05b7288dc9b2b6bafc861f0adfa62f7e564cd6272c0acf6154e02b9772fe08fbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf51b2c40cc2062791ed4d2914faaab666fc8e090da6acc234ad83c858ac854704c21baf6cdbbf9bce4f138c5b5f9a7b7955;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d39766062a3361d34b70899be53be162de64bed7ff836027d97d09d1e4cdc04ef74e76e7ddb93809685808fcfda7d749372;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5578d9fd29636d249bb7587b4b785d8624b5fe49db74f599482d6431afe786addf95d1af2ac18400989e59e76a4a5a18a5d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff912c8c4bd67e82892e1fde933d360563aed2cad46e4805a88d9c3aa3f0ed061fe6f2b2041901969fa35320df3e35fc192;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d22c3d9038a33e5b62312ca20e0cc2532be01f6da1af811aa73fb081124f32e43b97e4b61d71264435ddc2a3be73ae3da79;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cfffa6dcbc451d5b48b7a6878f9eb9d3f5c928e31f868946b3e3895f1ae37a5cb30ea7fc6bd992345d7066b20c0abca9da9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1225310ca69f589a8f559638e3ec81a5f260e706ee477805c28fd6441e26d23429f3d47576f7c6f07d8364c7e57f838bb635;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fec820d7a60ca8f9cd430c56c9818062f44215367246f8963d269675e2d096746aa2a5e898dbe8e4e2ed61e1da8b6e485a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe1e3dbba982ab2680b8084205e448922a8f09734f6b6aab1eb3911cfd888a5ad20e544a2266af54c5e969e2d4a5f0552db1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc080daab473ed036bfc5592c7e4401d619861e74c7075b807a6a1284a565499ef348db557d6c3d8f9c96a91664114d3dc2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fcf4673d4225fc3104182d44066ca5b3bf0c1e8a47aac4f93ffabc9e27085262b0035abe80d9cc118e72b83b8ce01c748c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h344e06bd0123a4fc6b1ec366b5175a01673972310a993ba7b5f7a3686113e1ff09f1e5e3f802ac3122dc70479cc647a1f674;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a26fdd4eeff39cf008f90f2c1ce88c6483e909fc1f50d16b9facb6a962246c0026cf55ddabf01e91be33428fe6dec6f12e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf72906e44b500544aa8812dc50dc36d1f5d74dd90c642e78540368568e03b958de3af1a5b33a68205456c8799388629e7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3fbef3a0f15ec1e93098cafd5042808e9caaeeae5c14fe8099c0b4defa5a28d266a862889ad382a4c91e458fec55a3424cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde2ec200f8f2c6bd789463392da36a6f7e7f92152a0c25ad1b1baa841368275a0fee43f6398f9c13366efb0c37d93d4e65d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf93f9e03d1705117fc96f3601586dbfa976bc0a8c7b9b45f3ff6cecec3319fdfba375907a1d7b6c3ed5f1cc2b6a25e4eea13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf98aa7a270abbb5046433b5b420eabafb37e221550c1d6e2e3c6b2014be351cec5051c98984539af2096cbee3ce45dd80eeb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d3df35573e590212aaa529acfb977f91e3acca1a8b320f76ac15371f7e13729d3e016d20a19866d77a2378640dd275757c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0180fc1a07563d36069bb9fe0eba787f0087a53bb9784343d131473f6fdff56fd4802093897e5b6082743e155c427893c12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb41d683833983cae04253a2db291a947ffb3074fcf46a0d752683dc952a93c8181ebcbaf6832656d5270f9654deeea08b525;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78247e92f9de8d6d6098076c5690910a894915a9a32be7c6bc3e73aa509d84bddc27efb3318c170fb756d9a3543b578b3b32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5b8ef9339ad9d97e3da3dd3921e026c011b60af28c59fa43d32e5fb6ff25cb42ccb319eeecfc41791dd57ea1ebb32ecdbc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd83d6f2fed55a9359ad449d35d1aed70472cf9427ccdbfa5a826304c96dfafcc0659d4eeb02d5572e81469864ba09d2568;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3289f7984f1e3919d940c8f5a904d3a704b40260e41af409d1648895a0b34a0425d06da72a75b4428076c273a88e03fe9aa9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h193d0f9670b21b029b242364a88af9313992da8a6ab67228cf8f9cc34c74952750fccbabb08554adbbe7b4c76160c0e7cefb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6692a062c75736935a6ad87c9a8f1344622c4614451b1c02453465f7e807da92a722b4e1c63620580cd26f74f5cbd7a9f5c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2e23b6e62bddf8973b3da76742ad89d610de97cb7d4b85c95c83308d88c84f4f121f20f88af611fd6c2203db8abedfbb2b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fc42d79836daf7760423c243d7a58674347b08e2a94f427c3aeec56c3910012727656f235e09bbe1592d45f5f599381c50e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3720b50fd8c5fb31e5e20604c20015d0ad10b4b545d89a73e89764281314e2105801117daa41fba4c741856264eda1df905;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ffa886bb77614e39b676822334a5f166d862b3c5a3cb6b9ac33be02cbc47691fa9ef46b489c2558a896d0af5cf0d7511a60;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb76115cb959e62433034b473d978949dbbe81ead3dc21413c5a30c12924a457b8b8808dab61c536cc27ed1a4831f32023471;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf65875c149514d92342777ead16d4f5d66db934b6fe87998e3c059040cbf27702191f31f937cb6b6a5da3b04e046b70b29eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac5e12793b6525a83acab3538ee75a1d5fdda21fd220bc5c771ced44b93faf9c1117993d5ec4424a87a4f91d0c8c20a3cb4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf612568b07760abf8ece2060d8449bd02aabaab2d815d7c7d411a5812c34bd31d6402332450dbf148c49f102e10b7cf330e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8bfdbc390d3d064f15a0e28db49fb214e0927473027fed0d13b9879c995f481c7703f4aebbf6424f6a7b342593da3988edd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7993fec15c946fd23bfcdad0f6388a03a48e8c330c0524175e0c406f79916134ada225010eb268829e6574ae854825055290;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h609d3e1196240d3aa12e9223c809b3e3647fbf8ead45517058ec8e432de8842ca838dec4cb425aa1532974bdb39c3353cc99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c27d9c364f08793c9856b88cb6f6bd3b475c8a58707299093564ca8dfc01bc7e71d3d49843dcdc76d76379231df5c162867;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e3d75b21bd706714953475984e28fffd0bbb9b3e9bc2b235813ea44607a0a1cba9c6be13fc9ef16d4778ece0c05e9f8f40e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb305ff74c740303297aaebb64f08321f451d9a5a6cc8f24e7e638dff7b97936e19084b4d3f965f9137735c41ff3eb3ef076;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7095119f8a4a9555be30a1d79ae3acfa63e45fbf93fd93de6221e96bc17397ae4a94c0efd3750abf4b3c870bf4d59e55217;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h618685dfb3148568d701853cf4b783b061813db480b1b89ff9b09139aca7ce1cc60715bf5cd45022f9b293782b7bc3948b37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3eb2b1852b2a9cd16d6c0ed59304f1cbb66eb11a91ec9570f86ad1d6081fb9a7e953551c19af5b81e6d9a9eb33192af5ff32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a5c47e687b2f9264d36c9e387a96729af5896af037dc8460d5abb77c6c61531a8bbeda8d2ffa8230e6621f6ab25166145ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b11e6c9799d344df2571c1f1b211ea7900d3694d7803f3c9539b07caac2dc45293b9e4ffa912429fa1ad8b314b512a32a34;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h965c2a5a621106113897aa16e30f167f315061a441a03f71a2497d45fa19c70d17f4bcdbe0b72b5dedb7d46186b8672f164c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha28ca63306b0a49af55a9d0d4c236a1eb43009eb142797bc141678119c49e82e2ba09befa122904818f4a436d03dd272129d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48df94e5122ea25d30da6e4f5ce084e6b1c2a226c23fbce3e497408d84ed8ebdc2ee44c725d1b44692311658b9a0ac38646b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a1ade7766913c79a3162417c8977be76f08b531adfc810f509447c1852054472dba453787ea286f9e06f395c89c8e9bc6e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b07a1f9c53b9a1ea0e8af4fca97809d35e678ad15c857772493c543f01f38e620eaa51acd4a44ca1dea048241a8a25cbffe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefa25116896b95409e8d9e29397640bbe31728504fa9c86f28da1a3f62fb6ca35f817ecf0a169654f4da02252c813902ee8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74b5c4515ffcafd90451552e4af6c201776550d699a27d1ab6689c7a64be069a55e6a84b9db4951d2492cafd5e209f934ca6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e29523a4d8ffca7b93b7bf10e51738fd07a625d91b8a50951cfc07b6404f495f0f4f7bde3d3e76c4c31f1f878885a72451c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ccb3454f8f1d4ddda7e4b9bb29cf6764a434c835197fcf54730f5171358ccea6769991acd1937d598761ad447a53adcd26c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8ef15a450ff6fdda0e5445f870f5af73d9a5b8318e19047a0a648a3e5548d77fbe5a388a69a46d392910b9ac6cb29b0d1fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd01232cc77a44cd13df7fcaf34fca9f1b7c840632907643ce1a60164e3ec68b4a276fe57eb22a6df5eb6e7b0b8de7f22fbb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5401ce9a2d37dddaaa0118dc69eee642915178d3ee8d0e3f04f83791d4b624e20b11a54efcff2439465026c1733b244c4b63;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9088f4fc693f7096c5d99273e761bcfc4db48e2e7f7060b221bde4e66fab3d58913db3452692115be2667624f8b544b3d589;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9be16c40d63a97453c678bd6cc4ed7c7bcc8a158c9db518b1c0edc525a4745c8135d59b8d8c8a42165c46d444a7dcf50671;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e9c5ec4962749baeff8ab2bb5e89a30bae92e493b479faf9d94c586c6c9c7a8a3ed10301757886931f051be96781716370b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59fb4b7d8870a96fcea2006d86392f1684e139317be86ea9e6a1dfbef24558575ac7b6fecc8d8a5e3fae8041009310880207;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2c7a55a27ba832ad92ad9fb923390b6dc2fa98e81f3346b81e049642168abfb4426b0bdeb3f32a7ce6abf1eba99560459e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6991e13b696c66754f5f879be8e4a0c7834bb34dd14bff1843e75667c7c88d520d292a7745c36c90a93195e73718b881367f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9b29bc89723a642feb5bccb14ed6bc5cb075743ac16a572b06a971b2758112acd7aca8771d1270ea48e6ba4f41e6ed1f5bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc40b527c3d3c857257f61590048818d3a4e1715c486364eaec6bd47f1a370d3f5b2f71278a869e0fa3860dd69f41015804b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb706ab23540db9fddda7209e9266303c80e4a68fdf97418160fe131b8163ecc8c46e93c2e6282d3db4f51b503c30899947be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8d546b0e028dc2da84adb2387380907192c77dfc334058f4f2817c39828ddf5e3d132845a4e6ac03f63c6721ec220316c02;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha636cbfb863d519a86c8cc4bd9efa3b157d990c60997eeeaf6b7f30d79842e63bc8cb4b5d465b09e9bd85562ce833559dfd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h733650888a1c0d76a4d9fe6ed489f8a82985a4fff5c6b261b7bb74ddf4a47f36360705bfe8db0ee9a3ebe7d7c8bb17d84f39;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7aea84b9f27c2ab47303dd4f5f11945189c3b268d3fe7e3e7401cdb2c3d31f16e545fd5dcd26b993c4d9c7a4d4f3814ecf8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4965a6f4c11b7a0a7a2db1396c85d55fe052f90e9386f14301a2cd5d42ff8b9745f0950aa1850a0a7c722803ddb02648ce01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9d53cb8b93d6188b59528a3674e23bcc3bee23ed8cb373a606ec209b8ea9caf21a2facbf1cee8d75d2aa3293da8173f5dde;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a265fdd95117891a21d699cae16c05af0691df61ec08a7fd7fd5a78bbe67ba0069360c72a35d694f608a8e276ba67eacebe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f7e100e448589f743f26cd07eb628a169f2133624ecd278fa78e16b23637aeb64b823a15b8309d191cd4693ff7a284b81d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15318eeea9e8f2b40d2353aee342e87c4a521a058bfa9de1587639ede40ddd274d5d4c83365f5894226fa80e4853445e1f78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb04a3943a4b16742bf11e6df07e37a38fd44a80e56281dc5653606591f716a1ae9a3cb4b7c418464a79b1253b6fe6b333c2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha150b059a4ee6cfbb7e27c343bc780d2b7b1d721153e48d42c5a62dbc85be64b43e5fc42f4dd47557d7f23dd14a309571aec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed511bfa7a8c225833da693383ce336430c6b538127e2473e8cb28a8a4f0ebc1db43a3ec36d4dc031f896b314f9e9496f7a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he823d0c7afa6a6ff99128821416d358ce4d73e0bb2426ab346dbcecbe948ccc4e6356623927086deff750abcc794fb87e43c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h235224580e3d7ab6b39b8e86c0b1fdf16abd3ace13a09e4bb840a79a915210abc2d28dc70e4efe225aaadbbd63d2c8430ab0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5010870b09fb60410e5594ca6374fa51aeada2de923250be51af5ecc62ca25101188d4ddcf9fd18364e4c2cadbaba5578ba8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb47a0e33e1dd8d6eeeb856144cad606a284aae6dc0094224a8949b7214ea34d0a83e0652851371a107466147d50184c7a54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9645173d6b16555a9d45728421b51fe24e8c64b578cda122e729453a2935986a415a9581f83b6027b4e6ee9f6cc74a65352;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13ed4903a54efdaeae402a9c2b28a3d8ffdac438fa96e80705a64cf4647da5a3e7e73a84ec626a0c16ee823caa6c2fd6816e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2fc6ce877807aabb390cb7001f899e93750e42e0eae26edab8b6e16f9a4ac797c259a1de83e2d420ed6ec96e26b8d661f52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fd017c70ab28c821233743e34d67bfb67e1ae382d6cfd056adca497adac33a6aa5992972a28516068970322897c55cb4f58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27469bd768d2e761f1d814febdd8023cc2697902caf78858b921d1710cb7ea6b780cc74feaf9a51fbde4db7819e76c8c8126;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd8b7def697d437c8a07cd1ea08444fe44d654f2cb929a6c0207439a06c2895d213d7ca899582a597b302b122e1c6125c984;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40e6cf717ee3c7dc2bf788d3c745231f8624a720c7629e33a8858db4621dc2bc46e3ca8682dfbc7e14e75e295fcddbf3aa41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dabf0419d5a37a35c2a543ef77922458896cc08b3a62d085d131986ced5769ea8c6bc2af211301f0684d7729cde3cd3923b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43b89f1a449c92d6f0f216f140f430112d31afd2341b466a4cc6f596430d442d158f40aa344ea63038c1313c35754385ea80;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h840ae9dbf2ec7c02ce1b2c82f133031738e95b07c39b45203baeeb1e014a0faa20e64eb0e258a7c653f2d2fbd649d0e3e8f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h353197fd42778d856e8717c4331d7ce1066aa0440d2980e7cb62263e303657bdf0c70eb2d7a6ea719aa9f4c4e400cda604e4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbeb4d5fd0b020114f45c5f522b6dee29a72a8b52ca33e143353b13b085cd67bf938b61dd6b8b29f59565ac935337fa4cba8a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc257bfe16358f1a4a1191cc52120f096c3d3b6e31978800a53b303c39c8f70ea18f57a22e9147acb64b3e00cf74c2ef0219f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb58cb656587caa43b39766f95de1566f85e32570a48640a89c7e815a7da4e249f37d56614db81f4eca60edf310f1648a6836;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d75b147881588e7115d0ba04dd2188a0cef89259bbd6dd59ae572efdb016cc2ee619ac038795c73b9928d8b91d0a3a90a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3f472ab19ef03a695235e78d1b130731e09ef14e9e7a0799912ec0ae20646aeb984f29128e2bb3ce79a9d1440b0ef1456f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50c05910a0fa3b6d63483c5f3441b4c16da494136f2a4a30657d49f1b42147c1aca3902c7b58f0892fe441cc1b3af6d374f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f697f27171bf554ed5bc63731a728304900b897073bff1928be143d0d828af5b762030cec800639e7c4bb36fe1fe986782a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a40fb26d775e626bff191bb1a1b800d131af1c5921f566164a3e031fa482067adee9ff37797c03488d8946f4c680651c060;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a3db636233d5479ac234104db3b9ed060f4d1995c596c87c7353cc7c49cb7bee8d308c26113b73a7694a76ab7072c4f4ef3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d4bcaf7f87c89e1a3f030c42a0cb9118fb900f291ec66b10c26074b039101303e3dffa0c111db21dd0a74c88573b5acc9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4adb88ea8d38b1a85976da05eb3790076f4f0ec9be37b36e26691360202c796721281f0382811760617babe7c612badb4f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85ca80ffbe0df0f7b13a5d9f1c1af8d58f903a7ba6b7e9cb27d6b8e5cd81f5c0e50246b88fad5f3226085e9b75ed6416199b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc84f4538dc511fdf94fe7795a26bebe4c3fbc2c467c6d7d6fbd0aba6ffbabd3c1c5a66f0bdddad0a6f008298ecd5d6245cd6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h866c705958d6c24e3aee79aa868a47e80ee62f3993b0da6cf9fcdadf4bf46c80517c66b32efb441f6c99cbfbf80b08a5429c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb4a84b91d250f29371f2a6ebf88b719b936d8004cd213b0b569edf2e58dc00853fd1ae24c632850dfe26da7dac42f174b29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c88b012877315d742f8c862d49decb01e9ed3507bc47d486cd9f7956734beb22fa6f24dc7d0302763bd8f93c7486da63cd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dd344ea1a622e90780f52ccb15477cad315a5e0218e4b4a8039335f326e84db76638ebb96184da14cbc3c10036bd6061317;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d79164abf776ff2d1995af37a81cab6087e8a7864c2a0664f5fa390c7c50eb59715b0bde9fe9b840801d82e9a94025e92f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c9be97add82b3a4e5e6ae274e2273a5065a09b177972a3bbce09504bb320d6d5c9b2434f34234eb032f2ab0373a6503448d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9330b9567ae75cce75969d63b08300b270f7a8089a073350cb823969ad4c37e8419009a7bc011bc6cb0256d8d28440f53bd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he03cb48b0fa3c13e160796f204c930fbbce80a5e9b4d7de539be6e0fa1472b950da5360225d8235b68f6fc90f40348a7a758;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc36c3b24f5311c46354b660828eeb82ff80d40456a0182bba5fed75d92789fc2a312496bb977d9982c041245bd76cc4667ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7475a40200b2ad31ec0ed5663e1a2c164ac7a6e4b75f5f4850f3fba646d761de615f43a0d01584bf04dac95f375fbf9903d4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd560a4679cbb3b91b5065e39729f0f4af820fe528b7d592503fadf4c99676993fe2989cc60dfc8013b1e23d30b03f9fe885d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88133a13f670c76567e1247af69c35fd6ed0cc12d7e4e9260521e1bbd6e3b4d5e275d78e809e7d7e261d0f325ae43396b6d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca366bd6f25a7b238620693664a585821be7e28fd272675c9a77502f8450f7e38db9121d01a533a893de7bd13a852917d2cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3d4ce8b061fb263541c8db181c4030c16dde628598e4ab03ee5d0bb823e9d81cb1e6ecbd626aaba0cef4fb6630a5fc246e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h391c7a2c85b2cc1b1bf1460d60c995ec39724ab6c96bf7710da2b250f81a073546b16a11d99ada389e4d6f6aaa8505ffdfea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3799c19f113c0f15fe877a74c76dd311a7b566b8dab58ac07feedb1a1b674ab45bd128e34727925553fe74fff23d2cb7484c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2134cb6aa873d0f99f01a6df7ba653cbf7d9c85b0e56eb24ede555b991d40683bc87a651939d00b94db168d7bde9519bc906;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h772cae612d361d73e3b4ec68fdb0f24dc2c8feadec1f8a75b708bd5ae09adbe0b0b2b514603ffc555df00ae63f6dfef9a682;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c77cc215edb30dac2e35be5ae0e7e86adbb04530569b1e8f76c290852a9eb4a6b9f4cfae3128ddab84b64552bfdab522c1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3144249e2b36c28be84d01385c16b9cf454f783809e22d1eea8a6cdc392987b475168df68d65f1eb23bd5d0168bcdf09ccf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e0db09be7f38045965b65a8340e257d56c7915959746b7dcca5e8fc124cd0c27e4479c62c45df8c45708d888d9617a54cf9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f731c608ed0a0d96fedec048ba4e0e9f90fab96ac581bb3c910b7cb58f7f8d7cb7ec73d4a9998836700380764b7fe43bf22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d1c0c6cb945b58dabd9a8c8c16cd06b4bfbb02fd1b4a56949f847d47fa96322d5ac8043e4b664376e73f77f011da74cf4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha71b412afae05012f51c53ceb19794803f0eaff6c82b8572b158a3fe52af3165afd935056ac97130ed7aedce033f95ca36dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2ff3a2eabca8f42a9f65cc99b875f2bdd0eec0ac22252631d3a8391eb176c872ab3f2a7afb026419e8ce7f3c9b67b21c8d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heca1286c5becfe79d2d375bf2cd04394ce0bdec59fb49d95de1c83a2823eb41d0330b15d171045eb12f23ebbc7d4f0398516;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaa8411bb8045d09c276a194e955853fc6c392127d2b3d4da84b5bd4c29047aea954ed924c0f0acf385bface8f86e34a2b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45a3c1bd4c621e2d8d6e5af429a8930dab565f03bc19d7af5f97a73373bfe416f2f3f43b5ac403ea16a2ed0ffd530a4e9376;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he44f00f10abd38ee4ccfa0126a891c17919ff9c519f384db95c8be34e63a2388a71b82adddf83cb648d0970fe41d1a9ba0d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h842dcca8f7a2e837d48a26c0bffa0b5cc34ee9827c4e060c59dabf3054784f4cefd1b54871fd5640584e6a058db36108df1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e78a9d187fb8b6bc292956c82a250f403b1aae0067ad8c083943e11401dd07daca023ac356ddfc861cce81967a6e330cd2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99817519eaab36c6d5a539e1d17b38c308d35c7bf364f2c971545e48b7c47573f4553ee84f53390884a5a6741c610de9463e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e0a229d1fed76d956385284e0dd764862fb850068c7d32dbd907cd7a764ddfc8f920334dab8362711400b184a25c11be4f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1efa86be9ad2f6f4c740989576b830b99fdbc7bc9dc9f8d25e3c04f3d4ec784021d0f1e7f65880349975ce5bba7099b47e84;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7d9e3f1e6bfef9ec9cbcf35255007802eac8ff06503b4dad22ad3122a1950cf7c8ab7b83f6f1f9bcf41c6f96caaaf51c7f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h619ccc81eb8ae4214ca8f062263af920e7436cd1379e0d97361a58f84d1e2fc8fe88fbc3ecfde68c2a6fcf780680a4b94c3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71d97eb74596e5712815b05df8cbb9017fb5e49463ae5fa7d5b826623cfacd1c0f65be5576de73d1915139aa0df4f8d3f3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h859cb34c88dbee6c5ce6aa9f538a4a1a73076423000420010b1dfa97e92511c0aee3f48986e93267ce99a8538b7f7a410df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb6413d8c48894636dd941b7f56a7696a862232c0baa553809050d5e7e358bea6d935d882903d077ace4d85695953050b415;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he41ffa2a5a60eeebc66e4703325ee6a319a7e8e1e24cfa6657db81e1f20920a52ab700c870f46995ca875664a3cffecca56c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8290de50295a89fa0f5adf7b15e32ea435baf3f172db5f6202b8000f018059f6f50e2730b77b6ceedc55190a69f537db2e25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f9671c1fadb169ce1e4f69effb096a678def046f8d794c383ece4cad66af6ff3f23909cd24041a3bfc7282409c3ad730eec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd1e706355ad44077688e0ff2d3cefcd237c2ac3a755c067f1a4463b190a453a1df285043472aaf5141dedfae95ac4428926;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb815b7ac86e4182ae6c4dbe3484248e3b25fd486fddeb7be127e2d5674325e340a786a4b17a2c816a81d6905ddd30f76ea5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h585c8157a2dd37ccc8892237268c47160a78e8adbb024e55f340da7e850a696dc4121b87369515af10797eafce9b71875663;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee19e963723ff2a274eac7002b280ab6cea30abeac1bd7e28e00689ba2aecd8127ed7aee33ac5978c5a678d89cb8991a6667;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc23c1195e6bb0ba2a6811826b05925cdcf74c98259badce087a7eab1d443b95bf42cc88d97c01324db8296f2dfd64eccf51a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aa7ef7c0927722b473717dcff5dc3cde59b9a80a1e3860b82945e3f2e173ef18071fed54e4491db824aa35576312187cc00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f4d45c4eb771fa3e25600b1f439370bdeee5881ab04d09cddb55e84c363d18d0d8c70e970a133e24c1eb325dfaae911a977;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h413f504811b896bba33e0fe5a3a2c1ae6dfe460560b3902df1c9b552d4cc229591ffcb1df729def2d57146110c02f93a8c40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4df21a5d86ee8532a2d0c83236f4b776e6344e3b1360d1b97a078b4f3f3a0c13f49c702813c6458b3004a26b2f879e2c7a22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9750b8476fbf8ee02bad579cec510915bbcaef3b1f5c1f76c8f69c7a7ecd935eca2f06e4edc3c14f66d75f8c57992233b449;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ad551cd4365eac564e77deb62998f3f26b0b8351e546af695e5bbc004c2deac78c4c80265f9d739b3df70460e2404908cd6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27331e15ba9f513c2750782ec7baf425563b15681b4e6157399be013678dbd0a508ccce354154112d09479b9c9b7240b672a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ea3e70889e0ad2e85a38c7b7ae865c78362fd66a6fc0784617a0d2ab13728dd0e0a9b5abcf4be71aa7597eb03440da642fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d06d9d5caae94aecf90443680ea2a0f0810cb2f9cd9b83bd02eeafc67a3d308b1e5b45bb2689aeeb89dc7fc7028a4ba74b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h268592c3774dd03a2a2760e1ae77cf524bb573c458cffa71582ae47770c90402398b7f4edc751450f535bb803818706c84d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24d338311b2e894a8ef85195eee71c6b2488312d287e60286ffdb5760028741934b04bcf4b6bc3ddfced730b378a8a1cc4ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77f35f53b2cfcc16ce35995e598df23493e5fb3faa3dfa3688d236bd8c8f413530c5cec2f6e1960937edf1dee85f723a744b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9e893a5a27fe7be205fe6c7991120bbd7541ec797958ebd8056e1eb7576d098611720014749efeed6833fbdc2c9dadb1d07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18ab1009c2c5914535f3f51c91bb3e10714580b8be6f9c512cf2ab686dcc13c1731c3775a46367d60eb03c61b9ce34b3fc68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd632438af9bb299b10fafb16611635905122391a3e23b1001f0b0c1254c135489dbd540ff441829fdfc813bb9e8562f2596a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76bcb96a991bb73cdb81e61b6ddc833018ec68da8b36705129d5370d0fb8cfe3359682b470ff99fcfc5be884383a0c34af7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h613537a8516e0b8a1996b60e32d6775af11634bd3670ae7921bafc69031b3901e86d188f9f2a4b944967e7a33b0b90038ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h731326142a0f7719f255222ccd3b0a593b21c8e72f4e0982186984e3d3eda924f88fec252eb08ec2f6594f5dc479f5953d16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64fd7a581149e07d2ee3b76cbe5da3a0fd907306fa558588aaa6a0ba0898697b43c7248cc8c65b7f3428cdd853fc45f40a34;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1d5d3154a2db8524369b3d815fa9df617fd13c3ccc937268e7f82247b7781d6ed7de6f3b13aa4cd525d779edbae883d2345;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he47f309865578439f8c1f44b15c0c9d97517d13bb761de9dd2f0041af6b4cabbabde780b2fc39a870f7ff2ec4a77a4ecdedd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d65633c9e3e700b5c08d7d35b2acc6682e26f7917c5529b32e02770918b3714e5c091c6fdcf38bb8bb33c4f9e314dcd467c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8faa3cee8b8e0673558f8b569a67d4db8b30168a34366db2767153e4ed230fa64fc1ed19219d54e82b9f5c00b24336f4fd33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd46af6b1f1df6b2e0bcec52e1ee82a56b803e0316621c4f2bbd837a1c2f453030e52ec3396885d13d39d03cc3c4e595da2e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82b135df8064c0c50ce889d2d22993a6f5158fb7817be657a68bf2ce9f10828322c99df197ef74309d1ae9a568c0625f8d1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb4aec3d69bdcf440e5c314e1cc6f24bc6b9b734ead5625f4f9aad4388d8e66db5121dc2ca3b0a6d6fff949fbda7a687c34b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ad6d7e53e6282c29523773ac95baca454daa6f2d42afd5d98a9e3b5037a00a03e2362369f89c3ddadfa53cf6165f3a6e193;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb345ad8bc881b8e6b78135e95ebf30b54469ef50e701311b9b2099764367817ea171c444f77d2f935bf2f7c6af9669afe21a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff27edb9fb66e46f5f3e4d8e83ddf833fd99277d0c18a9d94476595092fee416c015eeaf5022ae684875c6ba0beb142d9860;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d2487a5b6e92470b18fc97b15e65b4c27d777a274852dc3ff1a58c0a78e4fca4fbfe20bec515c38a0c527020a63f7381938;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd213b482acc59a17364b398eca05dbdd58492cd6fcba49fb27f8c34454b7d18b71a2d482caab1ff63959ff2de4f3363222f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7dd9d77523ea5dd636277b3633707b328a0a3911d7281833308320f94a248553300ce48f7ed9f2477efe7cd7d21620a9b7b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4727dc7d03a4a12b122cc101e3031a29f90447133172d793f9fc5d248174b894fd1ea911962993d4abf57834a83f7d901199;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ea94f4909efa179fb016b27c5c45f2d6591636a4217c5a3ba753021dbd1b372f7d3606d1d1e194252014daa2e71385d60aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0f545990c2e39b37d8daf1590a1f4cf70aa3ecc8704e03f0fec6825d42dd5fcb2161ded393318a1909610cf1034677330d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fe3e4932a99a6861f9d1931ed0d3ca9839de1a42a88cc3eea66efc7bc1475a68eca460460de431d3f2c194467058fc9a8aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h455a488cbdf959a3a5dbf826b80d56127584770f85602118fc37b71b525ea7bf202c5d24a6fae7bf331422a93be3870a4735;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h126112caa6c4ad453540cb6af2f37029cdc47f553c9b2dbf062826ec82760a2db0fb5f6544a2a7347845573d2a211ba8684e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5e16ce1ed29b00a4c80fba5900cb0b4c37343174465554a7456f6f40824611b7b6f12a8cb122fbd9e94c8d86e4b8657484e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha48fad4c934edc84d798ee78e72baf2f5c9baa08fac419c51cd78fbe24be4513e0f53b01bc03d73ccf96ab7b94a42823a93e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe2ecb3c2cfb4cfc26ccf8af22a8a8a5666028b76a8abb5589748c46045a3699aa8760fcad497bb36ce697bcc11ee8125873;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h274f3421dcb5e9ecdd6ea75699b2c80d28e8c9fd60d4bbeba50c20ba76b3678f78f1bc27a89b4cba00d200524d17e3f4441b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7b0ba8006bec2812e5c65fa6180644be4a16ddc0a6407aa3296636f9d6a2069c134ca3db745c7ccd469a0e376104427c8aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he25461a896173aeec2cc2e03f682360c9d7f459ad1060e30802be0ffb41ccf0d057b2733b19998147c2db01d9e0069fe16d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda7ca2ee3c54d5d18af96661f3821a0eb187a564d738a549a8c4cf9305bd6fbf223775a872167768549bc49255385fb2b4f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d7e056b896d3fbf114f68f466b0a5f063e94a48f38782c145cb9e29c939edea1f5158f7e8766f236630b0a9864eab2b202a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbbbace33e3080f7c05d7a9ec2834618e01625af0224a0c7f43ec92cc6e5bac3ca8dde17818c38d6a1a2f846aea33f1fb883;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfffd454d0318fc1c680adccba63db12f00fa8cc6e40bc0538f6558e23fd2d35f67cf152b9bcac15599ce86ed4ffb1ab8c9f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f02532ae12259a022fa856306e4002aa3e363c3d649e6d600f42aa8ee2597bd839e57439772d465edc05592929225c4c9a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0e2e2ea47d7ed4e251d3111d47e051e613551a5a451873be41178264c4219861c8e2351009897dc945fe9d1d639cf1839f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef038bc7db9a24d7b9e078bc06ba248b04c281f79253da5f577d813a2804ba3ce155a4f3604c65f2720bce3ab2f226c1cae8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dd2fa8f71445d906ebc813b105459e19997267bedd7a08d019f4ab1e961300da3f33cc8fcc5203bd7a10d80a09bf662b17f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f56c1304aa98d188ced0789a720202a8a2e1e99210966715e8a80b0498361d339c4442064aaddb023dfc55a8d77c0058771;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f6fb4b648ed2a0d398bb4742d85834b4fb0687503cf9c89004d73104c760e502a7b74cecb2770b6751c67c879f21fb36f33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a51145fedf58a50a420dca95b6d97eb16230b5548edac0bdf102516b5c426397d328b5e60fb1ec7b88fbc739365fbc5717b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae93f5b4e111c0b201471ab918faea50b500a37869e5d80e5ae85a142e73f8c05babce32328cedf53ec00ab62290922d467f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc887172410787d60a9ae9df8dd44ce608ad7f768637b4b26bf2c5e9316684745489cbadfacb5f7ae99961589913ca514b35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45025f8e94a6e7eb97f30f79be27de2495c1ee49785b23b3041a767c4b3c31a25ce639d7ea32b8d33cf1d671f81982c9cb12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91d632bf1e27ea77877785ec27a93e3eb5a84bb06183eca50ba9a616041523cd3ded420bbe38aa5114708e51bbcc4fb185a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8851be29711c483f84919f1c1ef3e80c5886abd3407c09d645c6db0149fe8adf3f0d38cfe77544870bc2f86986372b76356;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63f4f16483a6e7ca349ccfab097ca554b5077d164241b1d15938e11e9a28888e2875f54afbd5a77cfd681c36852ea49515d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb26d4fe4ac9bd753b7d5de6dec3ee71616242b5dab46c846963b7f16808fa8da794f30aa32d902bc426b2bf776eb4feaf40a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72eae90e627d53154dcc4357b685c6bc0b14cf7133eb9b2c51f50d0c2e3eea82fc92e17d843e0daf758042dce1926cb5486e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h944a5def39691aa1cb387aeb2dd351090d8019865663d00106b539f2eca6ef453c9fd520f0535d383a80e8792fc5d72e7e9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b2b1bda72768a61dae6747c024199a9ad1537780bb5178ce1d139e20df4f0ab5d03b6a57e2a85ce369758bce4be69c04f78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7af180138d0370ec0f721c8465bfe9beb11a99a8f69ebc76cd037557a14cc5be795154df84c69ab9f8fdbfe4f71a10fe6420;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h333e98b0b4c63c57319292e70d3492a5f7f8a562a1385a1ba5947c0c9a9f877f2805e67aeb72e3a2d20593a4f4a5e98d7599;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedf927cf0fd0d25b44a8271c5cdc0bdcce1ed320e81baabfaf006ac89acc17ed090927675c46f73ea8d47f53a4d58dde0e30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80dce2e0c2266bd658fc71c2a6cc3097427d039115b35db9339fd72c15c881e7c21776f6eee5748033624da4216d463ed415;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1141cfda00049afbfc966b88ae5b6d73dfeaadf59fe27a3fc02da5bb580a9f50424497f73aef802d2240e9c032187555b59e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43e3357f0ba5ee90f15f4f24131d04c3da24c981307e591af7a6638eb118968011906ea4295324d93b23dc608a66bfe22a15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2ab35dba98867ad38c7ffa4b1826c2d53315e850bb53008f2933a0d12d947e49d8fd6a122180a684f2d365be4800884cb67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20ca9db9584ab54e3a2d331f12a5ff54491c01a119c2c1d636bb0b01e68005db0f08d4f08abed684140cfffdcf75a14b0c0c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21d8e259403c897175b54d5584161bd28a8ca6cb6e52c7f48fa37876f78e39d0900f4e9f1a62d1d211897cb1a272f9465d6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac7f0bc53f77f5be0a26e52c4f76e2a478ea1668bcadfe90f6708fde59d75df3184a5f655943bf5a74645f355fe75b5d1335;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc35505a86d048f1d79f3e2ccb34d6ab74d276b311c2a47d0ab133df46859d5bcfdb40fd46e0fca6478e6ad8a8ab302c7ae51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3853ef6073371a32875e46f07ea0d3849c61bf7906aabf51f8894b48fe334f147d44ae0fac27193f21c3c6d300fa4e687aa4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1454169739dc0c5a5eaf2384b151c1b19e4a0512845c987d87d2c96c7b9677882a4a1527f7f2e0684b20f9a75351f42e8d45;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had31cafb86f9dc023cba2a121176ed5ccb5d4d05a2d84243205a7837e4e3f188c0579e90d895ba15051fcf41eb3fdb177b06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h857a01676b6b2e29c0ce23ef4e8db1e1196d3fec3999650ad18954191acc500d879767cb8ab66dc87b54b814b5d47bf80766;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d471423f999e7a5e67fadcb766fad25c85b544fa3b46c012a8e3af503ca01e6bb0421f8b5bc4160118587596d0bf38534f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2f427addc2b61a10fae15cdd4abeb9b9ca82933e22321f7853f21a44861c34d1f64030363fb8405523558a9cc0fec9d1006;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacc23e5c67236421bc587005988f20f4d2465b402eaea0f8355d8b070cf2c8d191fa6595d8adfa9e2462c0751df60bb6c523;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb55b23241534d5fa9e0232ec17eb5904438db53ea45c260cdfe9c7af3e8129f8ae0fc9d8dce72bafa78d9273f86ee2f7772b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h844428ef3fea082b8c0c22f82453793d7e15c0581f576788eb251dbb7ff5f9ca40ce5a59ca0a852a66fc9d3c5cbb026724e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h241853fbb0b2856d59cd2b23438c88533097da6810c6fbe9294e64d35e37f17430c578829ba3c6fbc8575154d228ef78436d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11939084842f4f3ac587f2ad989cac9d5c22f172959178a4c0e67a33bc95415f65e3d843eb23da39b89af9c3d425bad0b75b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h969c0a3a157b096d0de5738e95685d5f228c829ddd6d74beac2a83d365a1cf8ee56f983628ab350cfcffcd95b4a20c9889dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e2dc22d258c924d74dd3cabb99abe6aa11b2121940209141873b69a68da853efdd8cd65b0bdff10adf92e26e8d91887174d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3df785a268b65676a9d15ee94b381845a35efcefe91ff1b075bf6a6cc25d45fe6fc459afdf1aedb4427d07472c451313e383;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46c1705abf8b038e31ac785d620a82273a3214e1894b06ab7adb6b6dd1343643d3fc2a02fb908d46b68c0922a0c7b3911fac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heec3b8d66df94b82eaeda4ec6dd0204f447596482e10b328cde2f8388c3aa7d66e44afbe72690d71c62372c61d23d8e07af7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3680ac33ce20efcf345397b7abaab4f21b5e8e8781673ca6ef5fc90e2c0e96cda2ab18d0d787927e6ef6acb298c4458041aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1683797b840b56b62cde87e9f6ca45ac9f22564aef815942c2e9b2751c648b757131fd90c9c7a2d1920cb2636887a5fa8bc9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70f65375814c573a81fa64c4dfc39dd20682f939fe1defa82645c23da00fb802f260b2e397e946bc6db136492c63b0dff11e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecd50a0a62c534c975d1dbff2f6b80e1615cc08f57d8379b858e5e1f9933c16155d72860a267868ff96ecdc689a5aee46a9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8d0f465839cd5e68bc32505a4faa3def040bc7bf8464786e72e3c094ad1c077c5c76b0be3cfbf7532ecd52e5a4d23e16a28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9165f85a501e1022e06a4ba9bd7da265d9399eb65520a55e6fb44d03d4af6b42fdac36bb67e9d4cac39056cc6896784168;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6daa7fc6f78a4cf100aaf398c339b94bbc9e9cd80dde066b0c077999b3ed91eb05a1ce2c6f71e3d9a569568ed28cf5746a2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd018241bd55fd536eae4a7473b5edfb7d5327c5f3f6bca35d346d69f4397820793d5ce4b0a53d63ddf2848410416f9de10f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h766f799e3c3e9d0e1cbfaeb890c341384f3879ae815d36bb16f21ff75da33593015dfa5e1810c15937b9698d29a0a9d6df2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfc7af99c700d0723e4907456089ea48972f701546fcfc369a0310b619443408aee6c714ffd75798d18031b7479398492578;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6430fe3abc4d502677b99e36c62e3e972fe0d0a7d04f25491bd858d5d5dbf7a5a74cf9dd69d9cbde42083fb7811842cb7ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3c24761fa3b0dd839c7a20654d7f229a23eeae1789d12669644b685e66cba45c0e36aac70455e621f743fa288213e91224;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f65810c404adb10df63e90904f74f89b2cc90d9208fb921890320f0d42df33bac05e677fc7e970526878463e62cf365c722;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbbe437175250794119666d7244c94706f8cd3ca91b7cf38ef58ad4743cd04deace6c2e16f7c7bdb30cb3aac732ea116f3c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h373867e32dab1ab945d3342b6d0c717cc576a87f252810aa570054ff4e4658da3c598e55c186da568f2080a86a65bc2daae4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbea36c8cecebd54bd62a7432bdcd21f7891871fa2805548d744fe39baebc0c24af2870b048cb4e5d055b533e6771199dad9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h231cab1f2a9d2ba875a28a78fe76fb41ee8dec008fb594d692a4c5a9cc86a2c45575d4f57c826984b5dbb639518d9cfcae19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4e3177ba4d10823588b6708005371c3cad3df511f73c9d24948c175f2140f77086e08ef429d3daf3337d3a316a063d4aaaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77839810dba04ad88f5838f4acc1abc6cc86a90826bcf824368f076d2dd2594e4bb4a7d9acc863131b5b8712cfa51909bcdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a63b4e74f7e974c0116b305869d18349e8abba8d56287758026f6d25e3d3c7b6b52af731214d13ccdef1a1b06faa396549f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fe1c9168afbe5b82b871756dbd11021bfa8b8f9d65d627069e7a9274e8afc6d6fe735a2501c0e63a7aba8dcbc927709f726;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87c209baa69266fbd43830483cb573d74b05260d3d7fe862250670956b313474e584cd2d0ee1b0349fc91535465b73a2ec3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f736df5056aa8986e3d1705deb7427c488cc86a227bd87b44266d6108dfc9e9ee44c88a2db3c0bc32121f386c078d81775e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha90075cc2064dc747a8eb6f796311c8983324a2b3766d7e5fe80039eb1ce498522d5c1bee11aeb4efe7ba988ad1f872d5547;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23b84f8065413818748f713fa31aeac76cf85854e3e9eaec0f5c857b5028f7480c315f5cbd7595e355c2bfadfa04cd55f259;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1691711dc901a69d51099e0ce26e2ed04949c161d8d04c24806d6f30f84171d4abef8cfc32ed65ba6f7151ce25a5fadc7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b87afed33dfa18c3fd4597a7820497df270e3189d8035989330cffae4ab18e4b050d547e27efd06532d7496a41ac6d5c205;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8841f76519057aaadeba75d824fc134c252aa756897810b790240d4994a1d175da823737df57a17add4dd2610ebce4c1c52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebd302019bda1fcc4ed3cce572f1b0c4bdb33991cca151c9b901f97061230c54d4583f226415cc2734336cc2b74f96c8bd7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a7100896ed13d037bdfdf25d5c006ff8c2dad6bda75e4823fb83b155bb93c6e5f3e9a951b24769aa1f831544bea30f2bc54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a3af61c563f314816a734366c48fc3ef16df4698ef02ee4945f74ce2ee5f9f0bef46ce7efddf8191c953dfc6ea7768f4b15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h664147f0525032db54aa17401ed06455ad73140c409acb5e74036a5914bc97fc7e97f20a3a5177026143dede5c9742296ad2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h517369816bfd42b534e49b7f4f2aa65a5bbaf6eeb850505979ede7de038f38d8ce9fd7805974224039bd4caff3b6c22df507;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cde833c6c17fca7bcfc6d388b13fd6e50f9d84b58fe1cb81070427c647428dfd9aeb1d804708a5b1d423232eda9b354bba0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h961935904af396ad922463783f244cd0a74ad5a68dbaa033f1d6025751882c7ac09787aad09719c5db8e264926f04dde0d1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fcf074e7bdba20c481abc319a1ba846b9dc3bb67a71e31278f0f5387d49eddecf27c908fdba57f649dfa94d170579733790;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h637fa9e9c10fa1a2955872fe6791c14f36d4b8f8dadf427db952073d464270bfd56373ff7c5bd521f1a8e3f71ac1b66e1442;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98fe23d02ad10cfc08765cd63f64f30170601be9f6c08433bbc698a408912c6f3d08f66d1ea5f6502340fc6021c98afd529d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6327d5c382cea2d6b95c960ec1b955c1b4e8117f4b6f9ddfb3d58e395440b16c815c5cea2121e99d17d6862d4cb072e1dae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22170b4d20193070d07d7b058490a33e221469379f45583d303b3af43e07d40bc04c40745afb2e53a4edd8becb88a13e12c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa5a15f44648217e301eae75b799d67cdbad3f4805473aced70d43bd6ce7042c75c55908d56734a222425dd92845c832ff8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68c205dc76d4d07f1f849e16084a36ccd0bef10c7f34d2df8c329465f0b0b2c3c0fe289e8a79ef33b39675a2e857b63f00a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf2e86a33c32084f7f72a564d7ed9d9c274f1559d4b04f9af1a535ef2d37bceed419eeff69dd48990f2df929e8e7ea072d96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha263392106d9e011d620bb5f094a6da4b66bfb4155cc5d6ef0512779795ce893ca561ee3f5f109d671eea0602abf9aeedc18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc065ed326afc4dd4d73ec078fa2656344627623cb751bdaf83e184d88f7b8bb2307cd4e96640c56902f9603eae2c62cdd228;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd55c279a9713d350cb40e15e43c725838ceb9eec3b93ba980723470e75b13f7ae7cbdb9cc35de6ac905bbff2548e5ac3e562;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc2cdfb342d89282a12fe0fce6f35eee259bdc47bf97dcf20f48dd78e29c24f3ec0a34be2fde3ca18e21d3157e623c56209d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27d0b4bec4155d6864218dd611dbb9f32e4625b8fcaa8fc2681e8f1991b442119406e720295d25dd4a35f9da50108671b10b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4450e4838c2bbbfbe8a0ead5981ef07b398d63557e16bf1112b0a31ad4fcdcb5455f4acf398931fef4c7c4dec5f300b9327e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cecd2b8b0380587eccc8befedbee50ee7364ee0e544cedc1621f0f168f420a83c9a48a9911ec06ea856070ca359e9ccf988;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17bc4c9029d89b7903f3705ab9730006ce5bd8c2c7782dc10dc9fa4774674af631487786d461582a756e5a93b98eaf300f18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7745cad29453ad9918bbd590cd5a5c00f367d7f4ba3322c79cbaf0913ea55276b5e2d70ce92b198f946aed9e5010b817cc0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66cad0ce1fa78e882b54f686129bc14e6775625627304d38ad19c50a8d9fcdb9ed9c713b0cdf12c5c239fe55ebd831f57420;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e482ccfae8ee51835c49db3b3d938d3f2819de8a4be39e5ad7e4754556f825127df78977be041c8f88795b44d82ed2ab939;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf78b2812380f7471617a975b0fec78cccbfe9ed893d607f6a48a953d9f6a135abac5051ee11b0796ad94004e3b2d4b9edec5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha082e0f9dbb9205162abf493dd8d40dd8b0db4d2969d7b6c61e2dfcf2fd297d24aca71d3aaab728493e18cd9a18afa04db6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb9caf87222ad378c358a8b24ed996fad2319bb5cf26acfe6d1dd184f0eb6af1217c289a925690b592026c3fa483f60839c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9602640b2e66d25c836ec21f64e93004bfff6206892f4f59c5f8d7af8794e3d432f3f71f154717d0cbfca8f34d696d20a6e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb439fc98f188784c217a8010e9d9e3f8b057a680738de1c85dd02fe321a25875ad45fedd6b38f675e35ec4a8d988d35ba80;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ac8d7a83dafcd6f1f5abb4c11dca8c644ce2e032e115631023c39ae4cfba7144ad70dbf0c96dc94af453422fe2eab741987;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6c2a7b24528dff7aaac80baca0cceae7ff20d838532b8f42c6dca674e05f68daea38e344d5a5ef77553c1fe458c685b60d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd50e163fedfc71ec1bcfdc9dd2389d573838ace9bb7ef00ae313b94d614f9d4c045f49e5c8eb7d5c7cd22f83f4df8846b952;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d6fe736f833354c76ab34fae175e65128293b233a80aeeff50eea0974c7b4f492693ac908c4405843abd4b12a91dd1107a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8b7c69de806e4f56d639924d5acf5bc160d4e882088ff73628d39d206131b28cb44323c86c1afa3a9375b89adfabfe64e36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h118db460ee0875ce5b98742e1145e15d441ffb8dbb50bbb225815c629ba867954edc400a0245799d826270bcba2bdf2cdb5b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf96db5a59fc236724a21a843e70d0943a3379f7e95bdcd0c43474cb9723454fabb77c8a10a5150d41c224b1fafb5ac559e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37df749c5c5cbb85e79df3e47b2a34d86e56ce9d5c7ac0c11a38b33310994a8072d254dc33ffae95a529187dd2350cf8e9f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcffdac859fc234c3a91f276dcb945c85e1e222227a5b595abf11a49c1280603a4c22ca1bdb3f7df72f87240171da054904f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2e661e2aaf82e5f2fd1780b336658c2908fe8eb3bf1f9fd9626363c724a18216b5b484bc66ccbb41b7a59169ea7835e17c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c8489b69bdfd983818e01afef1a41addcd66358bfa3b8885dd94ee707cf15e6f5c9758037542c12ea1ed130b5eedf3a7d8c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82a919de96f0827f7aa1ea5787e2a3866abb5f2e6892bf2b90eda50112e0ad42a26f0fe0f56c724b97f9969d87a9a436e7af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed8a2fe2f25ca06a2158f8d27d4f858092d8156e2441582e85e23d0d1e77680d3513128b896f18cdd2ccec3da764e3c45f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bc32b34b950d26be967a9035777cbc2bfe601b7bf820ca6a2a3b48338f730b1f375e6ed74e3b0166564f2812ee8536fa1c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5d761a79b707f69febc61574bb12d126eaee3e0f5af419b3b2c8f78413b1d2bcd3105a329c6313e02119d7e8a6bb2f79b7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba6c590513080e6b2f542df7b26a0acb9a7e320d4eae1d86be6e86675a50cfa8b2f6097929aa036af668b6fdf04858375128;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb10154298dee1ebc1766d2b41533fa18dc05416994df1cf7648fa5b37c19d005e5f0230d6e16b1a66c3b0f4379366833afb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha81626c58948b86027416df5b4c044658c6cdfe2755f3b13cce4a6c4e747a37ef19ba83213664509bc477b2e57dae98c5455;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecfe999e96d5863a53827232cf89a9656ebf3989be4435bdb9abdaa39b008b5c7b46cd82e4521316e6c0f713f4a8bf8e64a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e11869358fa6b0b26449fc93a061f6ac0f5661449a9e86231cd1b4d8549eb35c0fef2c2a2208aec9b18276794931900d4d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6e81c775ace80c2a04c3f102da771fd315c5d020a6b1184a653667f3e1798687c570c434b4283cafad68d6ac28739ad2c1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc09fad2e1b117c6d39ec3ec880af245d9ed4279e4a3c152425f0c8cd08d7ff618089cb7b67a19cf7c4800b4e8135f3acd1bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b512be88d13b10cf265c5e067b322310d51c5ff6a02a5a990f5a1692007922af26984dab87fad4efd2f47827b94eafd0d4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd54f456f7461ddcdc3e4b7ed16f9eae80d812b117d46612e64f706d4526f444b0d602be95f59d858ad75b497bcc242986446;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd517506defbe361f3c212a2fc15716249a9edb94c2cea11603d5fe68aab39c06f71010f623ee35105b0c286c422c63e5e3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6b8396aacaef2cc0e79ad01db0a2650f2316ec0a54569c2c489b205dfff7409e6ff68d7fb2ac3208962014e1e0d63821c35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4ed6437ea5c8c9fecc36c1475bc068c6b39625a0827a917498bed07e53bc16ef4e9e2e7fcfc934634467d5dd1723ab803b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a6d10ffbe03f13e4715c1216c69e5cd38ccf7dc2d7400ac908a7e51582ee779e1ce024beef5c00c888dbd1e5adf53fe9e04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb9ab829c51d80a2eea04bcb2d6b7174df52ab4d314d7fa8a3a9b23e3ba1e7eb1dfdb3cc65e5c593b337eca745d9353eefa9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc76359c227c961c2f1efe63beec835c91347d8ab1a752544d2156b2f4c6b87667f86fbac243886a67244ac8c2242cb0a55f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc557304cd402a67ea4d45ebbfe2aaa4c4311ecfffc41ed22262f55b26b38951bb4547482bb82110b6a9470188f0c9ea31290;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dc5dba861042193424d443a28d8100da44d089d5dfe72ec60a2c94e4a1324a8cd0d6c0303857e4a4404548496418bf0a222;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86c6cc6044f3105f799810a5d5ea0c17ed3a9088d3aa8db91fa12eb33c1ca7cb93e335bb7215ed8df2cd086969d1dd59d9f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfafbfd5d71c71b64ce31c2e4ad23918cf9071b9f58e38e7a836e30fdfd1a1da34844853c92ae7a3855b8ada7dc0609122eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b43e0b7bbe943c6e6271301d1593056a033a2060dd1998cd1a1522420b3a41b8f3d7f8a587b2bac2f890dea2e368f71d52f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f21879ebf9ff0e9745e17626b0ba0fab73cb80eeaf1e77be08d2cc16a68c4b431afdbc78aa71dc232ed462d6e7dd24c6eac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f0c29d93e9feb64fe789b8bee203449c6ea653574363ee8f4ac4e957520bec45bcbc78b6610fca9b1eb7aa35c03f38dc67f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b098278dab53729ec03ae4dbdc1e02f3e1af7bc0c682a2b695534858f5919919372a6e29285dba366b9dfc8199d20e5651a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h600946c6e072687e6e8dae1c8b6d49e4bb34796cd55acfd42387af17ea22e524973d55d63865b04336e928eb30dd29cd7260;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c0b27add971b90eca80173f53d7390cc5e059c9142f91c3dfbc34e09bbddee64ef8e8d73e207178d7c9362145fb1d40de6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec00efa07a337985d3330035e3c346ca4beea174c0ed86084fda090df84b24af72a8b180d11ab1369c1a88aa19168520ac69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89cf46cc46c3580f5f54cfa50fbbafe785339e2e5bd348ae3821299c828bf5a2c7377324271c172282b6c0770c68f0c705b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6606875a52494730e7ec68fbaac8f693fe93407cd4ed1a755c40953adc3524721bdb029df0422c374265d4e7cd3201c2a3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6af0478cb66d2fc2a66c53a8fbfafdf343157427354190b511b1bba2bcd093935966bb075c49452587ca4e4c3ee2d9c6da69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39b30c236257c3e41c226d47d251f90a5ed6b08b7f443c9b24eb0a2c9f127a66399ed186843bfa5aa9c80cf836973c3fd16b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5054970074a95529986d3eaab8decc69bae6fab62936711441528d015b2279df2531fe62b5021d2db0cc91c8478ef81dd1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5472acf2b42d9603709bf12d838a7a2a787a41eec0650f6523d8ff44ceee01c97f125d0ae066211e3ddeadc5176cce00a810;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1bef245e1b2f2580717be19599e11aeb36423e39a896623e46f460785224965c73f56c5e9d23402bcb9b8881ad7197ace3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7702899486e88aa67f43bab91af619167d67f6bb1eace8b8f57971835523f07926926b70ecea89c62555cec865f064124fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff728db8f40be5ac419f05e64df2a8e5f0a4036b913e186afe6f03e5066a8c0de08c4640b7c7099530ddea806dbddc7d6930;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ef760f159ee94c8bb2d2fc869b049466fa54fdcfa5b1906a6174bc86e712b7d7d1d248a0f6db3368241899408c000fd14ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72cffdab9a703edcb4ce7affdb401ac67a389953ec7fe517fbac1b88cad0a5658c8be70012010edecb445d55c14856babdd7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84247ee9267afd3d1e671332a279637ea21731250eeef13ed9df4159bbbd04247006557040265c7368c51e8f593e83f2c178;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf68c5f4095c49323208c5a521ddbcd841ab59d4d782642b1cf267b77831df411f8688ecc2ade78f72cde1a9eb2f280392a99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02f4cc89e336f3975f6f4717fe6ce0b608883b5bacd63c0b7644e9d06c7908528486bfc3b6eab578dd534c91d308f02f9a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3da5bcec677db84e35320afde35e56686dc690f843e45cc5c0184001f4354f348c042dac5bb157749ef672aa6c0a233e4ddb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h893521f02d7ec5d2d6dbcfd5a85a0e64683f807a0348c2e55c67873396670df0ed5f8b1f6203412d340135ec3dbf2b3669a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha523633ef32320e08f2b36d844fc9d6837bafd5d968813267c540f0aafa2d66e02b22077afe97c1b298423c28ad3f21be333;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf59ed7bdf8025dfafea61e1c4eb94b9fc10d8a48433e60846493a0415a198f654fb023f47813af243fb8b7ce11cb4d6351c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9886bad724538e0d834d964e43c94fa5892cec0974bc6a52d6d000e525fd15509eb53d9079201d1cc0fddda2cc280dd06fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h816bb93fe800ce688fccfc577675d7d5520a9b160880a34b34c561d0c64491819f1493a2015954ff2c049385c0aff631da00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h957f425076d86b1df2ea9324ac698797752b22a953dc17588b8c003257fc4c8a52196b1411490b372d39ea91a7bbcb114434;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50fa2088ce1ffd102cc396c8fea8e7ff7545e1c558b4120aa39211d0087811dd030050727960753decde87f772acf8edff0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd56ba2ab04cb1ff1f84708e298077c8293ec588f3be1152c720859f2d818a57f2a2b2d8fef79c8ecf7773c904d04d0c18092;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf97aae6ad8edc118f80908612368b5e6c44dec7a5d50a7c808434a16ec89ca98a10a77dbdde750b43d02439003b156cf48da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcba3f833f558109cb68608bee9f5950d700eae311ecbe85a69ddf4017c6e7f5a111039d65eefb12e71d33a524fd37d8f7fd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56107ae67ca96f120a3fa5aec2968720a66624106421a48347a2ac02d61a058e25836ed1c7224a13c4d77a78c2ae86cc917a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2fd83b84843a8d24066c570de6ab9de09af54c65eeec392a526dc1a23bf966aba929abb8ad7fb5e7853bf18ade1d220ed54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h638c207d8a1c892b2ae2159ad112512e55c66a5e0dbc893ea0e35e10bf6ff503c4eb40afb00daa147086a3732212450b443b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf54023a35af5898899e2f0c55c16aef3faec9ea7ed9fe9ccdc09ef9c1a4150d252dfd40e7233277b43821d8f3c865b8988e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h707924a037ecb7a8c5679ebc91e2bb2037bb59546879aabfe13312ecb9d63c39f06f04808e82890546b47884f4dda4452df0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79e4e60a16c8c08477e495575ac27f97c2222b038f26f6b5a85bf289a93a8e9e7ee52d7f20526e94488c9c0c68b0949951a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3511f756e81cfbeb65e63e0df2da1d8e1465f746497ee45b22e1d28cac68299524c4998367d036748ef4dcb0f6c682ee94a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a440c6fec3a6c6b83d12d11af6b4c1324eaec8b446109537a795dbe88c6043534d9b040063e3e58c37511486b45a0ddff8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b57a3e1bd78375c5b8e8fafd5673bd82919f9913d523d9c324a9fa9cf90860a137b7ec8e1c2480253e72b6e5054b905e239;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdc2ed629171869c94046fc15444617e6f22ae85967b1ef2b0c6a90463a40be8816e0da8bdeb847c8a1079ad26fad4c39f17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1783610ed97ca600977cfa480676c5fad50ac46c0f65a7a574d685cd2f78ef0bcd764127901afee6346f8142afb9431196a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c530459d2dcc0df5a33ae8957a959cdf05f2f7efbf8cd9cf77e0013df0b1b13cfa0182fce5f416bde877691a27cd9b6958a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f5e193e49bcbdd2963adb5b6a2d5819005b9c57bf9a026beb526f2f857ae1a7392dc2090e916a96570f7386a7acf79306d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ae6a4c26cc53cdc3d4d40137181aee11beb70484873edcdcaadb9459840eca3316c9ec6f7f3d295ade888eece1f86cfb15e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fc1106922d0f497f42db8585aa8023300e6e4a1da3be20f185372fdedbc0b7d548acc5498b507d28003ad07d0637a677e46;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfadef3c9c1e3114670aa61057b965ff4d0a28e1055bb425f9fc20e618fae37c31ac1184ac95fcb16a08f0afccfaa28a6a250;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4dd8df93f7293fcf447dca1ac57b7024e9749fd1f99549ffecc9003cb1db0f72d3ec8db17581f7ae93450a1a06fd5cdec3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f9c12f0d775aae9f7bc0f3371efa678d6ddbaf9de96e0b396ec8436b23d058191f6d6df498498c862b58592a49881ea55cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2561364387ae926deb1968c8b0aeadd690d7e1b9fc5c6ef9d1bf8953f68ea72b5ab9078ba6b6b615877d27f1c4a66203b9e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h873b7011997a8a5680492678e8510b863965f9f19d75c7d3176d9eed6587573abe63a1880c4dfdc2122c1a4f0030592de041;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc46dc8b09c8fdc44e32989712ba9725117d043fcae870b64444e881c23c2448f9c71a5ab66b07be27771221ed3c83c2561;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb56c22e717cbee48a528772ccf3cb97c2b280bc0db5ac049c795e47fa4f22ba1fdf762ba7c26084642a17172d7f2d5cde846;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e95fe66d7b6afaf0eb5d745621eff7590b8e4f6d24c74a05896e01e7bf747a6c8ff72980be2c2c999b858691645345ce4e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5de983a1bca0591d1a20eb30164efa85a94465cd9b99c97304af29453414942ae40df8cefc1970fba9d74a37180e2fbf79a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h732f82667a0b80d90095feb9df30815b9e9d55ca9992bf31a0c24f5c4c6db637531c74b0c2ccbf0b90584e713289522ccb3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ec5a27e2b51d12b363f1fef2112fd72a72b78cbd6b82f6c938e2f38151e17f27de1edbf52901cf2918e5cd021eb52e08175;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78424badb78d617c077dbb0e47000ef227b8c3b643536bc116120b9c85774ea7ade66af98878ae1969063f98910b75fd6205;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47bda749f0b4e2486583a8d32d2fc3ed252cd13f896c03b2979f3557f08da5bba05ecb77291dec4daae0d1e910a553dfabae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h258aa446bd882ed5bbc5d91fdb962ce97d984ba0f336e3966e2c2b76e13b919d166e1a95b3eaf310b022fc512195d85b1ba6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3197ddf811a4559b96b543e86ed0dce4c86a28fd62b93a030f9f72e544cdb50996061acabaf69f561d9f922e6569508610;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e890469106dd9c2ea0b0937788c610a40c14f4c83e2885916fbd9cffbf8acd9349c3a058e75bbf686c54af235e91eee2f10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f112ac2462a68fe51457fe37a1e309d5f26f3e656cce593bea8a0f8ec22ff0587e685c807b04de48ea1c2021a46244c8939;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b68f6a0cde64aa1c52cd826972d3fe5753b2e004d00523d913f692760af96f9ca57d71c4425804a94593a11087a10d464cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h105059637f144865ee44cde4b538b03252a44a47793e2a380c0341ad07a4b602d7e207a3ab448a4e77f42e80963ecdf7ed65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha95386526805323205a7003dd273650a50235c48bf7b84a2ef4a5b29b503e49c989b0fb40ab6d5627ae2f075d2cba581870d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6fce4019ddfd11f0d1c6cb7459abd9ecc88304c2ffe8996368fcaea7f08ebb66ab45d04585d4e4d81eb9420f9ace994e565;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79b68fc632a3ad5f738d67e102e16bc53243577df709626cf3d63f11a0abb941ebb94bf66561ae53a94b10c7081437930fc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b0603b539a71277b60e8750d9cb5815ea5ca21edd55a1bb3281b7208192411fd261b280b7dae6b512db61e3dd8540eb526d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6c111fb696f06b1f3ae9c90c1d9c0baf4a0dff90ea6bdb7db7ddc3e3098a8847ef233e7ad93413675ddd3c91b884b965514;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4882367fb26d9ce5c5fdcff3294801d1f89dbff56fa9cc6caa24d17ea76d67f138438d8f0eb8b15a26717a3d6d388a69f47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc299c9f8a38052469a4b96b8c5e1b46968081db89ef33644b737095e8b41d7f9d0fe3839d3ea1c2e74b3f8bd4c9a4edac43f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ed21b6741f6a6417901b316569dc6f69558e9ac0b1c7bd3d29c811fb5f0773612cbcfeca514662a15463d9cc843a2c41123;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c8c4911bb9e5c4bf844364c032bede61f947d56fbf72427256bd60429208d7dd25286de43807f4b710aa1899eb81ea90c5d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa9f687a9e10dd28988fd0c93439b475781ea0f7b04b884d326bf85f45dcac2ce89b8e4253d8f21e77b4887cc36125098950;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8481b4c4b95dd23e8459dea7db3dfde81db6f11580dddb49961af3a6ed195405970b9b4fc8205c2406da0e69135e47866f0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16915e764689bd49f00dc0fe3b7fca62109f83fb6d781f8ef2d9a33e1eba3d3fb0416264ad758708d8ce1aa3a6b7f2d4f015;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59ef57e0204cdf94a4d6bd39c6bdd236bf8bfc3f12c1a225965e1f4a73931ad0e113cbb9904da43857bb920931a79f986019;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93d371e8eda0c0a49dc4278b0b4b21f0a0089b2d919d8def781c24305f56aeedcd17a5a2aae733d13fc0abba240fd9825ae7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd82755ca71a87504cec95d5cfb0055445313be5554c552b360dcd8afe37cc47c9b65093ad2098f207cc5535dd9b2f14eb83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h293e7649b971129fdd5a08698c972106c3eaac81587341675c83f3e6e847025b7bd8b075ba734db24c655b13bd4f6a96cf4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea68d35688155417b5e223b56e6e5a013f11f3646519069cae573c961d10fecb45ad972e8d46698c067b70ca67ca429934e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c24140f2208fc8eed1271f5bd3d69c811d8df8ea710b03e0f8d4ed7fee87dff3c1ff7a737f150c27834ebc944d6d803d706;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e065cc0fa9fa9edc13068bd8dcbfc19197c2ed1d24d06d87d392d5e558ef87adf58ddf6fe36f1518b237d6084d2c485cfc6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c29701616fefcbc99f03d8873669ec55d5d1b0801a57b67a8ba65923ab20d8b750e0c95bf07b7622a0bcd81dec356d4ecb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb253a6eb27bf9880a5fa090dad942ea58debfcc49a7877d6c69c645a15b7e89794ff29e6296e38a2c9596535351ce4d0c74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6c6744072aa44912d60f7221c998c75c6036752b75be55b760b8af1dc3f58f3bbf4e55beecbda0033e20a2a433e525499a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe43a5536608220f5a17230435e3c385a919a60d36c49df5d6d3d92eb22f6215c5388634427d651c688cdfa67f77d045bfb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed9e96af5d03e1df9ce142579fd2361a44e4a51e87507709aff8892f083e101c2849fac822932c708e9460a57d791e6d6bb6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha77ca18aaada7fae4be3d2f6b229128cf97b02765a7d9de021e0a295b5bf74161e0b2a42d4f2a8f9ce3876696ce563910aab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heee6843bc13ddf4cd5dc35a71cb8480c7eb53d7e1cd959bc203fd75b395f6e6107d08dd17c506f5dd92145010d386c01265f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c2a0c47ddede386f56809e84bb7f55c6062cfedbe5bf5a6f83af4021c724631319c69f16c357a18053374d3bc7ad26b2c7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf57f534a4d4fce883404543bea9ab3b434a30f2f0dd064d34b1f4479c7ced4eec817babb565aafbd54eee82b699fcc3ea5f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f16c057e5cfd10e0efe8186b46000e83b86751e882970db0df6cda7e5c974cc6f8c3a252ce78fb703cef98c186c65ca87d9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd258471b8e24b76b5629654c2f87d0a093d74bddb16422f5718bbdc4839dd18e43305f90e5e51fec8217e3ccb92fc5ca0b7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90d2171b694853fe890700a9c30258959ea4099008d6a34b1b5e2f94a8aa793ec14ad1ecd122697f4d53ebc09e9060a7577a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfa835d0e61439feb563fc79d9cb9659486cce4b9ab1af2dc0cefc444375e5914e28732110451dcb84ac06763f0d7bed8270;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f2eb9c16126dc5062f0714d28fe79b480f78a612b0501e694410a03952d3b5d87d8e443d5766e8ad796b05387a0afb165ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h122fc00eaa9d8fd013e5353f7f7d5458bc0d4c0636ad9be654a529d921d6a090cd75b10e77e256c6d2b0084b08d1898c8085;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadcb44ddea2736ce682be53322ddcea46c3545aa7a6d90ec39bba54eca21fd0566a606495f515ec8d98198f24c6fa4128e36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2eaf57fdca240fdda43f0715154114271d3006c16d7ed4bb7f38d8c9338f9df94d9876b6d328110fc26369cfd2677143358;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fb946016ef7c068cf393ff39c1e7c2ae487b3e350154d53d32ed667fcba7625bff03571440ca3359a5e6f924c4c507eda32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2b19d7c7df0545b430d58de551cd19eed2d92f1da264f8dae1f63887cb605a981c2fbabc425b29a16f1decc710bc0890eb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h310910a724ff1e051a1bd55868092690e6c1bf506d888421c33c524eb995fca31dd0f7407ee3d1d5b50187b51a426adb8671;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa3cf4e88b302efb3998d98113b57628623f9ce2894d96bee2041a84333292993ed536cbfb28d6fa5324db06847ebc171293;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dec417c7f437ed8dcebe072f3ace183aa88a2429a4ffb8fc8bc5ae7d41a079a1817adb86273f3875c099c468e897496a2aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9943f24a0a544d602f3bce929ecc5a52e3648a9bab5a42aef677b8b2f1df304da62bbaef7f20ca5e4e798e3ebb4646538a4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf421f4a392ee9365cbdcb4a3c3dab10834c21b2ed820d6c14d56d324c989963f8686bc3fbf50c1d12c6d6671cf992514e96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3aef16fc68dc70e70ad151f3866b2971ddd9a8b37c12963b739060b069e2fb3c555f0715de54c5c38dd7e71ad9ed001441ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4d54561a21b177445a68b04252c98cdf3f2b0536ff1665c8ea64e2021cb5f697722ace89bf0469af9b848941e496aa416ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d00866d36b3dce52eae0825acf6124dbccf9a7aeb2d1778d820fe62e8b86b5515d9d24fe5f65327d7c74dee5d82b2e12020;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc304202ca7bd03f06f19763b12400b6f1214dafafc2fd7c4a2d09c07173af5535a9f28985738bd6347a160a2a305d4b990d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1f979e75e78e1b73515d4c0700206a39d1b54eca07ab2b1a846f3b6c16966bc7eb0fee3dc584e39692b537df5c68ff0700;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e5fe8fe261d2d755f995569f5489c257675e466c8b1e22655fcea949e36168b255c88a80ace606639e43065693a021f4e19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h241be79441a4cca20733c5266727a1137dbdd19a3b32e74522f08bb86c8f9b7cd40ae189bc978837923f22bef32155b70d5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70eb1a6b6e3091e30bb683a455f5b5c20961a7b47769c12b879e3599cee4a9556889005419dfb63f07a56c12083a690c5a8a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a865f8492964271a72202695e858987a96a3e61ee161018cdc9bf0059cd4e7afa30cca438dc1660298a718e36539c3b4278;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3428c9a6a6c0e3d3cd098caa39ec3c2f0ca5f1ce79cf907276c09374ff2b86860944f5b2ba4a9419a35e1d84c371adb2290c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75a9aa02fc985eed82276ac32a2e21df00134321d3aa6b48ec5203e073820fde87409c632d98a8f25e99eda6220ec8fe8f74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaad1293d839663f6a5d62754ec92298786a67889a176e4e3a25d67c68d256f1eb3deb7da4e1b24f2a96d18a2db2bf3b6739;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfed0aa7f58ae3702a4cddcc26fd8fa4d06764b1733486b76d4c235ad8fc1650bb45539798de943523222f5a2bec2c389c8bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd12598df282b57eda2c2f256f3c4510a9c2bb6b259c613a163afbb1b23d45ab2b38202275e9c919e32d80edb0db22c19732b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb80a6feecc7334ef4fe99905b313c0493c14784dd26023b834c7bb80c1b99a5791acd73ede1920220a1c22bd11ca488c877;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b1c04f59bab44cdf5ed44d49a9b839c0b47d4d4ce8d0acbb6dff5545499af734e3297e8aeeb73847d6ce276fd28bc75748e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdbbabba08c5d7d09b3c518ee025b5cf0f9c999351a168fc36c1aa5b35af7184311775515640a6826e9280a986ccf3ddbeb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb651cfcffe99ec67a466dbac0f517aaee42ecd10e08eebca08043c9ddd65ce27f999f5c46e1b8a6a8387dd375053c93f9e72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94444d7798008bf568e70d7b41c25a799a6ebe5b360a9fa7f2ef3fc85041fedd8976caa26141e1dc9d2719f8c30cfe907470;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81b0bae7661d74334d1e1ef378a44c3b73f2d14a5f0aa5b5116b4e648d92a5a915b9cdd2ad5423e91dd8eaea1249e83fa381;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35c7e280b867090e728f23113f61c5cda6885ee0a073334ae4f0505aec4fbf4c15e10ce9457bd0bd192b2f80215881a69362;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7896067d00625e95ea3a50e3228c229eda06e965e32439bed4159eeb1d1c3932dc7c6b4ca69c4048b125ba2180f2aff70fe5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had1c5f8970ffb8cea7b35498195c8ff5485eda085c442c28fdd3bb874c66b34ad765cf6c7d1461ec77c1b80a76251ac28a19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h871e29312f306cd0de23dfa9459bd52cafab8ac7914ea13ab0c8b77e11f35ad8f8f72be55c288c278177f779625c7b707854;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf5a92fb33d02d86269d64137cc5f09d483558974c35ee56855244129cfb8f198a4e98df6be7c8ce57b78ae1d8f7842a9a7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2fb8d252207393d245184bec08d875786e7aee4fd0cf9d2fd4f84e706726e82955165f30ddbc7e5aa6bb9818dc3c6161ea2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcfdbbbb50563ae02e2b5cd4a8f0ca60ef7663085d23e24dbb51f609654bdd2ba0bc0ac41b260890617eb086cbb2623d0823;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d03247bf1f9d770e5e576488768a5bcef6b5c21f5e4e78320a51db38a53f26a1fd7afe002010e1b87b00562f7df89c5d99d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h755547c8d044d5ffc85986fff412b9bb60144c05be98d071a86190e8f5bf42dc1312a0916c680bdb73a22b6f25588ae108f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3fc9084505de2998bd890ce875d878f522e1ba11251751534742ba1381b435f68ba58fa26dd7e51ccd40402be3a229c7e26;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f5ea83db9f2788f0e1dba4feb280a7b6730c98e82a0b0ada03120a7f62b7853e6dc2e6399c08f779d312d5f254cd7442527;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h582635d30a45466811965c4398283d581e56e510afc9dea7e8369c6996d679a69d58b75fea6647f4424429c855a6d215ecbf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9c3a6cea36e0ac9c6816ef0308c60b641b69dca98b5fbfb2ae79d36a4407e16ac2d19a488ae0005ee8b7adbdac754dd1f7f;
        #1
        $finish();
    end
endmodule
