module compressor2_1_32_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, output [20:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    compressor2_1_32_16 compressor2_1_32_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
    end
endmodule

module compressor2_1_32_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    output [20:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    wire [21:0] out;
    compressor compressor_inst(
        .src0({src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    rowadder2_1_21 rowadder2_1inst(
        .src0({comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[20:0];
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [14:0] stage1_0;
   wire [9:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [14:0] stage1_4;
   wire [16:0] stage1_5;
   wire [18:0] stage1_6;
   wire [11:0] stage1_7;
   wire [13:0] stage1_8;
   wire [14:0] stage1_9;
   wire [12:0] stage1_10;
   wire [10:0] stage1_11;
   wire [15:0] stage1_12;
   wire [17:0] stage1_13;
   wire [16:0] stage1_14;
   wire [10:0] stage1_15;
   wire [8:0] stage1_16;
   wire [4:0] stage1_17;
   wire [4:0] stage2_0;
   wire [11:0] stage2_1;
   wire [1:0] stage2_2;
   wire [9:0] stage2_3;
   wire [6:0] stage2_4;
   wire [8:0] stage2_5;
   wire [5:0] stage2_6;
   wire [6:0] stage2_7;
   wire [6:0] stage2_8;
   wire [7:0] stage2_9;
   wire [5:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [15:0] stage2_14;
   wire [3:0] stage2_15;
   wire [11:0] stage2_16;
   wire [6:0] stage2_17;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [4:0] stage3_5;
   wire [1:0] stage3_6;
   wire [4:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [1:0] stage3_10;
   wire [2:0] stage3_11;
   wire [4:0] stage3_12;
   wire [1:0] stage3_13;
   wire [6:0] stage3_14;
   wire [4:0] stage3_15;
   wire [2:0] stage3_16;
   wire [7:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[4],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_3[25]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[5],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[6],stage1_4[10],stage1_3[10]}
   );
   gpc606_5 gpc11 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[7],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[8],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[9],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[10]}
   );
   gpc606_5 gpc15 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[11]}
   );
   gpc606_5 gpc16 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[12]}
   );
   gpc615_5 gpc17 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28]},
      {stage0_6[18]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[13]}
   );
   gpc615_5 gpc18 (
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_7[24]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[7],stage1_7[8],stage1_6[10]}
   );
   gpc615_5 gpc19 (
      {stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage0_8[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[8],stage1_7[9]}
   );
   gpc1406_5 gpc20 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[9]}
   );
   gpc606_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[10]}
   );
   gpc606_5 gpc22 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[11]}
   );
   gpc606_5 gpc23 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[3],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[12]}
   );
   gpc606_5 gpc24 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[4],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc615_5 gpc25 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16]},
      {stage0_10[22]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[5],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc615_5 gpc26 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_10[23]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[6],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc27 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_10[24]},
      {stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage1_13[3],stage1_12[7],stage1_11[8],stage1_10[9],stage1_9[13]}
   );
   gpc615_5 gpc28 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_10[25]},
      {stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30]},
      {stage1_13[4],stage1_12[8],stage1_11[9],stage1_10[10],stage1_9[14]}
   );
   gpc615_5 gpc29 (
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_11[31]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[9],stage1_11[10],stage1_10[11]}
   );
   gpc606_5 gpc30 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[1],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc31 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[2],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[3],stage1_13[8],stage1_12[12]}
   );
   gpc606_5 gpc33 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[4],stage1_13[9],stage1_12[13]}
   );
   gpc606_5 gpc34 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[4],stage1_14[5],stage1_13[10]}
   );
   gpc606_5 gpc35 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[5],stage1_14[6],stage1_13[11]}
   );
   gpc606_5 gpc36 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[6],stage1_14[7],stage1_13[12]}
   );
   gpc606_5 gpc37 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[7],stage1_14[8],stage1_13[13]}
   );
   gpc615_5 gpc38 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_14[24]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[8],stage1_15[8],stage1_14[9],stage1_13[14]}
   );
   gpc1_1 gpc39 (
      {stage0_0[21]},
      {stage1_0[4]}
   );
   gpc1_1 gpc40 (
      {stage0_0[22]},
      {stage1_0[5]}
   );
   gpc1_1 gpc41 (
      {stage0_0[23]},
      {stage1_0[6]}
   );
   gpc1_1 gpc42 (
      {stage0_0[24]},
      {stage1_0[7]}
   );
   gpc1_1 gpc43 (
      {stage0_0[25]},
      {stage1_0[8]}
   );
   gpc1_1 gpc44 (
      {stage0_0[26]},
      {stage1_0[9]}
   );
   gpc1_1 gpc45 (
      {stage0_0[27]},
      {stage1_0[10]}
   );
   gpc1_1 gpc46 (
      {stage0_0[28]},
      {stage1_0[11]}
   );
   gpc1_1 gpc47 (
      {stage0_0[29]},
      {stage1_0[12]}
   );
   gpc1_1 gpc48 (
      {stage0_0[30]},
      {stage1_0[13]}
   );
   gpc1_1 gpc49 (
      {stage0_0[31]},
      {stage1_0[14]}
   );
   gpc1_1 gpc50 (
      {stage0_1[30]},
      {stage1_1[8]}
   );
   gpc1_1 gpc51 (
      {stage0_1[31]},
      {stage1_1[9]}
   );
   gpc1_1 gpc52 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc53 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc54 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc55 (
      {stage0_4[31]},
      {stage1_4[14]}
   );
   gpc1_1 gpc56 (
      {stage0_5[29]},
      {stage1_5[14]}
   );
   gpc1_1 gpc57 (
      {stage0_5[30]},
      {stage1_5[15]}
   );
   gpc1_1 gpc58 (
      {stage0_5[31]},
      {stage1_5[16]}
   );
   gpc1_1 gpc59 (
      {stage0_6[24]},
      {stage1_6[11]}
   );
   gpc1_1 gpc60 (
      {stage0_6[25]},
      {stage1_6[12]}
   );
   gpc1_1 gpc61 (
      {stage0_6[26]},
      {stage1_6[13]}
   );
   gpc1_1 gpc62 (
      {stage0_6[27]},
      {stage1_6[14]}
   );
   gpc1_1 gpc63 (
      {stage0_6[28]},
      {stage1_6[15]}
   );
   gpc1_1 gpc64 (
      {stage0_6[29]},
      {stage1_6[16]}
   );
   gpc1_1 gpc65 (
      {stage0_6[30]},
      {stage1_6[17]}
   );
   gpc1_1 gpc66 (
      {stage0_6[31]},
      {stage1_6[18]}
   );
   gpc1_1 gpc67 (
      {stage0_7[30]},
      {stage1_7[10]}
   );
   gpc1_1 gpc68 (
      {stage0_7[31]},
      {stage1_7[11]}
   );
   gpc1_1 gpc69 (
      {stage0_8[31]},
      {stage1_8[13]}
   );
   gpc1_1 gpc70 (
      {stage0_10[31]},
      {stage1_10[12]}
   );
   gpc1_1 gpc71 (
      {stage0_12[30]},
      {stage1_12[14]}
   );
   gpc1_1 gpc72 (
      {stage0_12[31]},
      {stage1_12[15]}
   );
   gpc1_1 gpc73 (
      {stage0_13[29]},
      {stage1_13[15]}
   );
   gpc1_1 gpc74 (
      {stage0_13[30]},
      {stage1_13[16]}
   );
   gpc1_1 gpc75 (
      {stage0_13[31]},
      {stage1_13[17]}
   );
   gpc1_1 gpc76 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc77 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc78 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc79 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc80 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc81 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc82 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc83 (
      {stage0_15[30]},
      {stage1_15[9]}
   );
   gpc1_1 gpc84 (
      {stage0_15[31]},
      {stage1_15[10]}
   );
   gpc606_5 gpc85 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc86 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc87 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc606_5 gpc88 (
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc89 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc90 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[3],stage2_6[3],stage2_5[3]}
   );
   gpc606_5 gpc91 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[3],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc92 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[6]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[1],stage2_9[2],stage2_8[4],stage2_7[5]}
   );
   gpc606_5 gpc93 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[2],stage2_9[3],stage2_8[5]}
   );
   gpc606_5 gpc94 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[2],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc95 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[3],stage2_10[4]}
   );
   gpc615_5 gpc96 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[4]}
   );
   gpc606_5 gpc97 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4]}
   );
   gpc606_5 gpc98 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[4]}
   );
   gpc606_5 gpc99 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], 1'b0},
      {stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[5]}
   );
   gpc1_1 gpc100 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc104 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc105 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc106 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc107 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc108 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc109 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc110 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc111 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc112 (
      {stage1_1[9]},
      {stage2_1[11]}
   );
   gpc1_1 gpc113 (
      {stage1_3[5]},
      {stage2_3[3]}
   );
   gpc1_1 gpc114 (
      {stage1_3[6]},
      {stage2_3[4]}
   );
   gpc1_1 gpc115 (
      {stage1_3[7]},
      {stage2_3[5]}
   );
   gpc1_1 gpc116 (
      {stage1_3[8]},
      {stage2_3[6]}
   );
   gpc1_1 gpc117 (
      {stage1_3[9]},
      {stage2_3[7]}
   );
   gpc1_1 gpc118 (
      {stage1_3[10]},
      {stage2_3[8]}
   );
   gpc1_1 gpc119 (
      {stage1_3[11]},
      {stage2_3[9]}
   );
   gpc1_1 gpc120 (
      {stage1_4[13]},
      {stage2_4[5]}
   );
   gpc1_1 gpc121 (
      {stage1_4[14]},
      {stage2_4[6]}
   );
   gpc1_1 gpc122 (
      {stage1_5[12]},
      {stage2_5[4]}
   );
   gpc1_1 gpc123 (
      {stage1_5[13]},
      {stage2_5[5]}
   );
   gpc1_1 gpc124 (
      {stage1_5[14]},
      {stage2_5[6]}
   );
   gpc1_1 gpc125 (
      {stage1_5[15]},
      {stage2_5[7]}
   );
   gpc1_1 gpc126 (
      {stage1_5[16]},
      {stage2_5[8]}
   );
   gpc1_1 gpc127 (
      {stage1_6[18]},
      {stage2_6[5]}
   );
   gpc1_1 gpc128 (
      {stage1_7[11]},
      {stage2_7[6]}
   );
   gpc1_1 gpc129 (
      {stage1_8[13]},
      {stage2_8[6]}
   );
   gpc1_1 gpc130 (
      {stage1_9[12]},
      {stage2_9[5]}
   );
   gpc1_1 gpc131 (
      {stage1_9[13]},
      {stage2_9[6]}
   );
   gpc1_1 gpc132 (
      {stage1_9[14]},
      {stage2_9[7]}
   );
   gpc1_1 gpc133 (
      {stage1_10[12]},
      {stage2_10[5]}
   );
   gpc1_1 gpc134 (
      {stage1_12[13]},
      {stage2_12[5]}
   );
   gpc1_1 gpc135 (
      {stage1_12[14]},
      {stage2_12[6]}
   );
   gpc1_1 gpc136 (
      {stage1_12[15]},
      {stage2_12[7]}
   );
   gpc1_1 gpc137 (
      {stage1_14[6]},
      {stage2_14[5]}
   );
   gpc1_1 gpc138 (
      {stage1_14[7]},
      {stage2_14[6]}
   );
   gpc1_1 gpc139 (
      {stage1_14[8]},
      {stage2_14[7]}
   );
   gpc1_1 gpc140 (
      {stage1_14[9]},
      {stage2_14[8]}
   );
   gpc1_1 gpc141 (
      {stage1_14[10]},
      {stage2_14[9]}
   );
   gpc1_1 gpc142 (
      {stage1_14[11]},
      {stage2_14[10]}
   );
   gpc1_1 gpc143 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc144 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc145 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc146 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc147 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc148 (
      {stage1_16[0]},
      {stage2_16[3]}
   );
   gpc1_1 gpc149 (
      {stage1_16[1]},
      {stage2_16[4]}
   );
   gpc1_1 gpc150 (
      {stage1_16[2]},
      {stage2_16[5]}
   );
   gpc1_1 gpc151 (
      {stage1_16[3]},
      {stage2_16[6]}
   );
   gpc1_1 gpc152 (
      {stage1_16[4]},
      {stage2_16[7]}
   );
   gpc1_1 gpc153 (
      {stage1_16[5]},
      {stage2_16[8]}
   );
   gpc1_1 gpc154 (
      {stage1_16[6]},
      {stage2_16[9]}
   );
   gpc1_1 gpc155 (
      {stage1_16[7]},
      {stage2_16[10]}
   );
   gpc1_1 gpc156 (
      {stage1_16[8]},
      {stage2_16[11]}
   );
   gpc1_1 gpc157 (
      {stage1_17[0]},
      {stage2_17[2]}
   );
   gpc1_1 gpc158 (
      {stage1_17[1]},
      {stage2_17[3]}
   );
   gpc1_1 gpc159 (
      {stage1_17[2]},
      {stage2_17[4]}
   );
   gpc1_1 gpc160 (
      {stage1_17[3]},
      {stage2_17[5]}
   );
   gpc1_1 gpc161 (
      {stage1_17[4]},
      {stage2_17[6]}
   );
   gpc1163_5 gpc162 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc163 (
      {stage2_0[3], stage2_0[4], 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc164 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2]}
   );
   gpc606_5 gpc165 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc615_5 gpc166 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[2]}
   );
   gpc615_5 gpc167 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc168 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], 1'b0},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[2]}
   );
   gpc606_5 gpc169 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[2]}
   );
   gpc606_5 gpc170 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[2],stage3_14[2]}
   );
   gpc1163_5 gpc171 (
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage2_17[0]},
      {1'b0},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[3]}
   );
   gpc1_1 gpc172 (
      {stage2_3[7]},
      {stage3_3[3]}
   );
   gpc1_1 gpc173 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc174 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc175 (
      {stage2_5[6]},
      {stage3_5[2]}
   );
   gpc1_1 gpc176 (
      {stage2_5[7]},
      {stage3_5[3]}
   );
   gpc1_1 gpc177 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc178 (
      {stage2_7[5]},
      {stage3_7[3]}
   );
   gpc1_1 gpc179 (
      {stage2_7[6]},
      {stage3_7[4]}
   );
   gpc1_1 gpc180 (
      {stage2_8[6]},
      {stage3_8[3]}
   );
   gpc1_1 gpc181 (
      {stage2_9[7]},
      {stage3_9[2]}
   );
   gpc1_1 gpc182 (
      {stage2_12[6]},
      {stage3_12[3]}
   );
   gpc1_1 gpc183 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc184 (
      {stage2_14[12]},
      {stage3_14[3]}
   );
   gpc1_1 gpc185 (
      {stage2_14[13]},
      {stage3_14[4]}
   );
   gpc1_1 gpc186 (
      {stage2_14[14]},
      {stage3_14[5]}
   );
   gpc1_1 gpc187 (
      {stage2_14[15]},
      {stage3_14[6]}
   );
   gpc1_1 gpc188 (
      {stage2_15[3]},
      {stage3_15[4]}
   );
   gpc1_1 gpc189 (
      {stage2_17[1]},
      {stage3_17[2]}
   );
   gpc1_1 gpc190 (
      {stage2_17[2]},
      {stage3_17[3]}
   );
   gpc1_1 gpc191 (
      {stage2_17[3]},
      {stage3_17[4]}
   );
   gpc1_1 gpc192 (
      {stage2_17[4]},
      {stage3_17[5]}
   );
   gpc1_1 gpc193 (
      {stage2_17[5]},
      {stage3_17[6]}
   );
   gpc1_1 gpc194 (
      {stage2_17[6]},
      {stage3_17[7]}
   );
   gpc2135_5 gpc195 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc606_5 gpc196 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], 1'b0, 1'b0},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], 1'b0},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc2135_5 gpc197 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], 1'b0},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc615_5 gpc198 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc2135_5 gpc199 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc117_4 gpc200 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc201 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc202 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc203 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc204 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc205 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc206 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc207 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc208 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc209 (
      {stage3_10[1]},
      {stage4_10[1]}
   );
   gpc1_1 gpc210 (
      {stage3_11[2]},
      {stage4_11[1]}
   );
   gpc1_1 gpc211 (
      {stage3_13[1]},
      {stage4_13[1]}
   );
   gpc1_1 gpc212 (
      {stage3_14[6]},
      {stage4_14[1]}
   );
endmodule
module rowadder2_1_21(input [20:0] src0, input [20:0] src1, output [21:0] dst0);
    wire [20:0] gene;
    wire [20:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[20:20]}),
        .S({3'h0, prop[20:20]})
    );
    assign dst0 = {carryout[20], out[20:0]};
endmodule


module comp2_1test_32_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [20:0] exp;
    wire [20:0] dst;
    assign test = dst == exp;
    compressor2_1_32_16 compressor2_1_32_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, dst, exp, test);
        src0 <= 16'hb0e1;
        src1 <= 16'h880c;
        src2 <= 16'hca77;
        src3 <= 16'h96e2;
        src4 <= 16'he5ca;
        src5 <= 16'hfe6a;
        src6 <= 16'hc84f;
        src7 <= 16'h5c89;
        src8 <= 16'h65b2;
        src9 <= 16'ha122;
        src10 <= 16'h3c2a;
        src11 <= 16'heb56;
        src12 <= 16'h14cd;
        src13 <= 16'h93c;
        src14 <= 16'h5fe;
        src15 <= 16'hde61;
        src16 <= 16'hbf30;
        src17 <= 16'habc3;
        src18 <= 16'he1a5;
        src19 <= 16'h3c8;
        src20 <= 16'h4721;
        src21 <= 16'he601;
        src22 <= 16'h3be;
        src23 <= 16'h20b4;
        src24 <= 16'h2824;
        src25 <= 16'h8759;
        src26 <= 16'hfe89;
        src27 <= 16'h6161;
        src28 <= 16'h8612;
        src29 <= 16'h7dcf;
        src30 <= 16'ha57b;
        src31 <= 16'h580d;
        exp <= 21'h1086d2;
        #1
        src0 <= 16'hd206;
        src1 <= 16'h52dc;
        src2 <= 16'h897d;
        src3 <= 16'hb4cf;
        src4 <= 16'h32a8;
        src5 <= 16'ha719;
        src6 <= 16'h10a1;
        src7 <= 16'h69fc;
        src8 <= 16'h2894;
        src9 <= 16'h1644;
        src10 <= 16'h1281;
        src11 <= 16'h80a1;
        src12 <= 16'ha3d1;
        src13 <= 16'hb705;
        src14 <= 16'h6a09;
        src15 <= 16'hb839;
        src16 <= 16'hfc96;
        src17 <= 16'hd564;
        src18 <= 16'heccd;
        src19 <= 16'h5f4f;
        src20 <= 16'h13e2;
        src21 <= 16'h81ed;
        src22 <= 16'h192b;
        src23 <= 16'h5609;
        src24 <= 16'h89ad;
        src25 <= 16'h1552;
        src26 <= 16'h667;
        src27 <= 16'heb33;
        src28 <= 16'hbec8;
        src29 <= 16'h12a1;
        src30 <= 16'h95c2;
        src31 <= 16'he99c;
        exp <= 21'hf0b17;
        #1
        src0 <= 16'h83ab;
        src1 <= 16'h49d4;
        src2 <= 16'h3a00;
        src3 <= 16'h469d;
        src4 <= 16'hd80d;
        src5 <= 16'h5eea;
        src6 <= 16'h656e;
        src7 <= 16'h54bb;
        src8 <= 16'he466;
        src9 <= 16'h9513;
        src10 <= 16'habf1;
        src11 <= 16'h7f53;
        src12 <= 16'h63d2;
        src13 <= 16'h2d52;
        src14 <= 16'h5814;
        src15 <= 16'ha26c;
        src16 <= 16'h40ef;
        src17 <= 16'h5ab;
        src18 <= 16'h5ddd;
        src19 <= 16'h4ce8;
        src20 <= 16'ha79f;
        src21 <= 16'h507;
        src22 <= 16'h716e;
        src23 <= 16'h16ec;
        src24 <= 16'h3e35;
        src25 <= 16'he445;
        src26 <= 16'hdd7c;
        src27 <= 16'hfdfa;
        src28 <= 16'he73;
        src29 <= 16'hd51f;
        src30 <= 16'hc964;
        src31 <= 16'hcc3d;
        exp <= 21'hf0d1f;
        #1
        src0 <= 16'h9649;
        src1 <= 16'ha38a;
        src2 <= 16'hdf4e;
        src3 <= 16'h8e9b;
        src4 <= 16'hfe16;
        src5 <= 16'hc889;
        src6 <= 16'h2880;
        src7 <= 16'hd76c;
        src8 <= 16'h6f2f;
        src9 <= 16'h74f8;
        src10 <= 16'h761d;
        src11 <= 16'h954a;
        src12 <= 16'hf11a;
        src13 <= 16'h4fb8;
        src14 <= 16'h9ac1;
        src15 <= 16'he243;
        src16 <= 16'hbdea;
        src17 <= 16'h6e5a;
        src18 <= 16'h6c9b;
        src19 <= 16'he1f2;
        src20 <= 16'h22dd;
        src21 <= 16'h1a43;
        src22 <= 16'hef86;
        src23 <= 16'had4;
        src24 <= 16'h9081;
        src25 <= 16'h7809;
        src26 <= 16'hf8e;
        src27 <= 16'h75bc;
        src28 <= 16'hd0bb;
        src29 <= 16'h6bc3;
        src30 <= 16'h2484;
        src31 <= 16'h9f10;
        exp <= 21'h115bdc;
        #1
        src0 <= 16'ha30e;
        src1 <= 16'h5488;
        src2 <= 16'h4226;
        src3 <= 16'h3fa7;
        src4 <= 16'h2f2d;
        src5 <= 16'h5784;
        src6 <= 16'h8071;
        src7 <= 16'h91c3;
        src8 <= 16'hfd76;
        src9 <= 16'h2eed;
        src10 <= 16'h4d9d;
        src11 <= 16'h31f0;
        src12 <= 16'h6333;
        src13 <= 16'hefd8;
        src14 <= 16'h2571;
        src15 <= 16'h38c;
        src16 <= 16'h5f0a;
        src17 <= 16'ha53;
        src18 <= 16'h7bc9;
        src19 <= 16'h7fe1;
        src20 <= 16'h3ec;
        src21 <= 16'h9d6a;
        src22 <= 16'hfcf8;
        src23 <= 16'h9c20;
        src24 <= 16'h4193;
        src25 <= 16'ha6fd;
        src26 <= 16'he04b;
        src27 <= 16'hf980;
        src28 <= 16'h811f;
        src29 <= 16'he247;
        src30 <= 16'h2400;
        src31 <= 16'had86;
        exp <= 21'hed0fc;
        #1
        src0 <= 16'h6fd8;
        src1 <= 16'h9776;
        src2 <= 16'ha77c;
        src3 <= 16'h2443;
        src4 <= 16'hb7a3;
        src5 <= 16'hea59;
        src6 <= 16'ha655;
        src7 <= 16'hf76e;
        src8 <= 16'hf435;
        src9 <= 16'h86d6;
        src10 <= 16'h3f31;
        src11 <= 16'he7e;
        src12 <= 16'h7dd7;
        src13 <= 16'ha932;
        src14 <= 16'h9150;
        src15 <= 16'hf40b;
        src16 <= 16'h1234;
        src17 <= 16'h4f91;
        src18 <= 16'h54b6;
        src19 <= 16'head8;
        src20 <= 16'hf6cd;
        src21 <= 16'h79b1;
        src22 <= 16'hd07a;
        src23 <= 16'h1252;
        src24 <= 16'h3e7c;
        src25 <= 16'h1195;
        src26 <= 16'h5382;
        src27 <= 16'h94d5;
        src28 <= 16'hd1fe;
        src29 <= 16'he625;
        src30 <= 16'hf6d9;
        src31 <= 16'h8a7;
        exp <= 21'h116c92;
        #1
        src0 <= 16'hc5db;
        src1 <= 16'haf3d;
        src2 <= 16'h906e;
        src3 <= 16'h6496;
        src4 <= 16'he92a;
        src5 <= 16'h6749;
        src6 <= 16'h3333;
        src7 <= 16'h39e1;
        src8 <= 16'h645e;
        src9 <= 16'h4c5;
        src10 <= 16'h1af;
        src11 <= 16'h9d6c;
        src12 <= 16'he95a;
        src13 <= 16'hc575;
        src14 <= 16'h1aaf;
        src15 <= 16'hc792;
        src16 <= 16'hb4f3;
        src17 <= 16'h54b9;
        src18 <= 16'hea20;
        src19 <= 16'h3bfe;
        src20 <= 16'ha681;
        src21 <= 16'h38e4;
        src22 <= 16'h9cd6;
        src23 <= 16'hf36a;
        src24 <= 16'he671;
        src25 <= 16'h7a23;
        src26 <= 16'h9f55;
        src27 <= 16'hb312;
        src28 <= 16'h653e;
        src29 <= 16'hb612;
        src30 <= 16'haa8d;
        src31 <= 16'h749;
        exp <= 21'h10e081;
        #1
        src0 <= 16'hbf50;
        src1 <= 16'h17f1;
        src2 <= 16'hf530;
        src3 <= 16'hd494;
        src4 <= 16'h5009;
        src5 <= 16'h80af;
        src6 <= 16'hf84a;
        src7 <= 16'h3053;
        src8 <= 16'h1640;
        src9 <= 16'hdefd;
        src10 <= 16'hb29d;
        src11 <= 16'hd93d;
        src12 <= 16'h5354;
        src13 <= 16'h3819;
        src14 <= 16'hd7f;
        src15 <= 16'h77cf;
        src16 <= 16'h2ae0;
        src17 <= 16'h2c08;
        src18 <= 16'h2303;
        src19 <= 16'hd412;
        src20 <= 16'h8e5e;
        src21 <= 16'h5e54;
        src22 <= 16'he909;
        src23 <= 16'he1e2;
        src24 <= 16'h53f1;
        src25 <= 16'h97dd;
        src26 <= 16'h858b;
        src27 <= 16'h7f69;
        src28 <= 16'hab38;
        src29 <= 16'h3421;
        src30 <= 16'ha3c7;
        src31 <= 16'hb29;
        exp <= 21'hfb0d1;
        #1
        src0 <= 16'h4a05;
        src1 <= 16'h1dee;
        src2 <= 16'ha8c5;
        src3 <= 16'h296c;
        src4 <= 16'h52cb;
        src5 <= 16'hb66f;
        src6 <= 16'hd1fd;
        src7 <= 16'hc29c;
        src8 <= 16'ha31f;
        src9 <= 16'h2fdd;
        src10 <= 16'h6faa;
        src11 <= 16'h63c;
        src12 <= 16'h28f1;
        src13 <= 16'hd8bf;
        src14 <= 16'h3d5;
        src15 <= 16'h7d2a;
        src16 <= 16'h9814;
        src17 <= 16'h1a68;
        src18 <= 16'hcf47;
        src19 <= 16'hd6f0;
        src20 <= 16'h1c62;
        src21 <= 16'hf0e0;
        src22 <= 16'hca98;
        src23 <= 16'h9e73;
        src24 <= 16'habc5;
        src25 <= 16'h3277;
        src26 <= 16'hd9e8;
        src27 <= 16'h11f3;
        src28 <= 16'hf452;
        src29 <= 16'hd08f;
        src30 <= 16'h9b65;
        src31 <= 16'hdbbd;
        exp <= 21'h1078a2;
        #1
        src0 <= 16'h31be;
        src1 <= 16'hdfd9;
        src2 <= 16'hdd10;
        src3 <= 16'heb17;
        src4 <= 16'h390;
        src5 <= 16'h5c28;
        src6 <= 16'h5e46;
        src7 <= 16'h65e3;
        src8 <= 16'hd15e;
        src9 <= 16'h3163;
        src10 <= 16'hf39a;
        src11 <= 16'h6ca1;
        src12 <= 16'haf66;
        src13 <= 16'hb8a9;
        src14 <= 16'h273f;
        src15 <= 16'hd2f2;
        src16 <= 16'ha8c6;
        src17 <= 16'h9004;
        src18 <= 16'h5642;
        src19 <= 16'h483c;
        src20 <= 16'hc99c;
        src21 <= 16'h7bfe;
        src22 <= 16'hd0ee;
        src23 <= 16'hd771;
        src24 <= 16'hda2c;
        src25 <= 16'h19ba;
        src26 <= 16'hb439;
        src27 <= 16'h6f6b;
        src28 <= 16'h10e6;
        src29 <= 16'h869;
        src30 <= 16'h57ce;
        src31 <= 16'h2708;
        exp <= 21'h1037cb;
        #1
        src0 <= 16'h8044;
        src1 <= 16'hd8be;
        src2 <= 16'hbb7e;
        src3 <= 16'h5d20;
        src4 <= 16'h3dd;
        src5 <= 16'h734f;
        src6 <= 16'h7393;
        src7 <= 16'h88dc;
        src8 <= 16'hccc2;
        src9 <= 16'h20d0;
        src10 <= 16'hd2e7;
        src11 <= 16'h7c89;
        src12 <= 16'hcbfc;
        src13 <= 16'h7ed6;
        src14 <= 16'hd521;
        src15 <= 16'hcd1d;
        src16 <= 16'h7dba;
        src17 <= 16'hce24;
        src18 <= 16'hb4ce;
        src19 <= 16'h927e;
        src20 <= 16'hd81b;
        src21 <= 16'h86ce;
        src22 <= 16'hdea9;
        src23 <= 16'h8a7;
        src24 <= 16'heb9f;
        src25 <= 16'h73c9;
        src26 <= 16'habc9;
        src27 <= 16'h269d;
        src28 <= 16'h2c10;
        src29 <= 16'h53e9;
        src30 <= 16'h1b64;
        src31 <= 16'hec01;
        exp <= 21'h11a1dc;
        #1
        src0 <= 16'h37c4;
        src1 <= 16'h1704;
        src2 <= 16'h1b87;
        src3 <= 16'h815c;
        src4 <= 16'hb9b4;
        src5 <= 16'h1623;
        src6 <= 16'h3962;
        src7 <= 16'h98e4;
        src8 <= 16'h6078;
        src9 <= 16'ha6d4;
        src10 <= 16'h830e;
        src11 <= 16'hf952;
        src12 <= 16'hcb76;
        src13 <= 16'ha731;
        src14 <= 16'h9374;
        src15 <= 16'h61db;
        src16 <= 16'hff43;
        src17 <= 16'h51b4;
        src18 <= 16'hc3b9;
        src19 <= 16'h21d5;
        src20 <= 16'he2be;
        src21 <= 16'h35d;
        src22 <= 16'hb318;
        src23 <= 16'h9c70;
        src24 <= 16'h9952;
        src25 <= 16'h4f07;
        src26 <= 16'hf9ef;
        src27 <= 16'h880c;
        src28 <= 16'hbf05;
        src29 <= 16'hded7;
        src30 <= 16'hd3c4;
        src31 <= 16'h7b74;
        exp <= 21'h113cfa;
        #1
        src0 <= 16'hfa0b;
        src1 <= 16'hc07c;
        src2 <= 16'h6ccb;
        src3 <= 16'he6a6;
        src4 <= 16'hec1f;
        src5 <= 16'h3b10;
        src6 <= 16'hde30;
        src7 <= 16'h711;
        src8 <= 16'hcb5;
        src9 <= 16'hf1c9;
        src10 <= 16'hc54c;
        src11 <= 16'hd061;
        src12 <= 16'ha791;
        src13 <= 16'ha732;
        src14 <= 16'h8720;
        src15 <= 16'h8d1c;
        src16 <= 16'h3cfc;
        src17 <= 16'h2366;
        src18 <= 16'h46c3;
        src19 <= 16'hb61f;
        src20 <= 16'h8752;
        src21 <= 16'haf5d;
        src22 <= 16'h191e;
        src23 <= 16'h4f51;
        src24 <= 16'ha968;
        src25 <= 16'h5f72;
        src26 <= 16'he675;
        src27 <= 16'h5277;
        src28 <= 16'h2cc9;
        src29 <= 16'he15d;
        src30 <= 16'h3068;
        src31 <= 16'hff8c;
        exp <= 21'h118dd4;
        #1
        src0 <= 16'h8db;
        src1 <= 16'h947c;
        src2 <= 16'habf0;
        src3 <= 16'h6bd4;
        src4 <= 16'hcb33;
        src5 <= 16'h8811;
        src6 <= 16'h7f60;
        src7 <= 16'h3338;
        src8 <= 16'h5426;
        src9 <= 16'h9a6b;
        src10 <= 16'h4f99;
        src11 <= 16'h2ed3;
        src12 <= 16'hc64b;
        src13 <= 16'hb90e;
        src14 <= 16'h5309;
        src15 <= 16'h8f90;
        src16 <= 16'h3652;
        src17 <= 16'h133f;
        src18 <= 16'habe;
        src19 <= 16'hb245;
        src20 <= 16'h4878;
        src21 <= 16'h5b9f;
        src22 <= 16'hfc31;
        src23 <= 16'h5a7a;
        src24 <= 16'h9a48;
        src25 <= 16'h7df2;
        src26 <= 16'hd603;
        src27 <= 16'h29e5;
        src28 <= 16'h3e9;
        src29 <= 16'h73ac;
        src30 <= 16'he0be;
        src31 <= 16'h30a8;
        exp <= 21'he2c59;
        #1
        src0 <= 16'h2083;
        src1 <= 16'h51b;
        src2 <= 16'ha839;
        src3 <= 16'hd0ec;
        src4 <= 16'hf8bc;
        src5 <= 16'hd19e;
        src6 <= 16'h7ff;
        src7 <= 16'h96c1;
        src8 <= 16'hd1d;
        src9 <= 16'haafa;
        src10 <= 16'h661b;
        src11 <= 16'hc4a;
        src12 <= 16'h941e;
        src13 <= 16'hd68c;
        src14 <= 16'he2;
        src15 <= 16'h9eef;
        src16 <= 16'h927d;
        src17 <= 16'h740a;
        src18 <= 16'h133e;
        src19 <= 16'h3773;
        src20 <= 16'h8c9d;
        src21 <= 16'h2137;
        src22 <= 16'ha715;
        src23 <= 16'h9b5f;
        src24 <= 16'hb9b5;
        src25 <= 16'ha9da;
        src26 <= 16'h78d0;
        src27 <= 16'h9fff;
        src28 <= 16'h3eba;
        src29 <= 16'h3fa4;
        src30 <= 16'h7b57;
        src31 <= 16'h52bd;
        exp <= 21'he4724;
        #1
        src0 <= 16'hae4e;
        src1 <= 16'hc807;
        src2 <= 16'h21a4;
        src3 <= 16'hf6c2;
        src4 <= 16'h5304;
        src5 <= 16'hdd3b;
        src6 <= 16'h232c;
        src7 <= 16'h8c4a;
        src8 <= 16'h5769;
        src9 <= 16'h4a99;
        src10 <= 16'h9831;
        src11 <= 16'h80a4;
        src12 <= 16'h6644;
        src13 <= 16'hc803;
        src14 <= 16'h5acc;
        src15 <= 16'he1fb;
        src16 <= 16'h218e;
        src17 <= 16'h35c;
        src18 <= 16'h7c33;
        src19 <= 16'h7f2f;
        src20 <= 16'hc407;
        src21 <= 16'h9464;
        src22 <= 16'h7dc8;
        src23 <= 16'h6c9a;
        src24 <= 16'hadca;
        src25 <= 16'hd045;
        src26 <= 16'hc4c2;
        src27 <= 16'hb290;
        src28 <= 16'h9d5b;
        src29 <= 16'h8e;
        src30 <= 16'h965a;
        src31 <= 16'h8a54;
        exp <= 21'h10ab66;
        #1
        src0 <= 16'h310e;
        src1 <= 16'h8afa;
        src2 <= 16'hd3;
        src3 <= 16'h18c2;
        src4 <= 16'h1503;
        src5 <= 16'h65ab;
        src6 <= 16'hdb;
        src7 <= 16'h46ff;
        src8 <= 16'hb4f8;
        src9 <= 16'h2d06;
        src10 <= 16'h87ab;
        src11 <= 16'ha3b7;
        src12 <= 16'h5926;
        src13 <= 16'he324;
        src14 <= 16'he9a5;
        src15 <= 16'h65ad;
        src16 <= 16'h4580;
        src17 <= 16'hd8ff;
        src18 <= 16'h2c19;
        src19 <= 16'h5117;
        src20 <= 16'h7345;
        src21 <= 16'hd860;
        src22 <= 16'h85c1;
        src23 <= 16'hd5da;
        src24 <= 16'hbaa;
        src25 <= 16'h2c8a;
        src26 <= 16'h20f1;
        src27 <= 16'h142d;
        src28 <= 16'h663b;
        src29 <= 16'h8f9c;
        src30 <= 16'ha77;
        src31 <= 16'h4db2;
        exp <= 21'hc2f62;
        #1
        src0 <= 16'hbc12;
        src1 <= 16'h23a0;
        src2 <= 16'h7038;
        src3 <= 16'h709c;
        src4 <= 16'h3cf9;
        src5 <= 16'h2fbf;
        src6 <= 16'he74;
        src7 <= 16'hae4f;
        src8 <= 16'ha768;
        src9 <= 16'h48ee;
        src10 <= 16'h7d8e;
        src11 <= 16'hf936;
        src12 <= 16'hee85;
        src13 <= 16'hd146;
        src14 <= 16'hac08;
        src15 <= 16'h56bd;
        src16 <= 16'hcefb;
        src17 <= 16'h9726;
        src18 <= 16'h9ad4;
        src19 <= 16'h12a6;
        src20 <= 16'h4939;
        src21 <= 16'h3b35;
        src22 <= 16'hfed5;
        src23 <= 16'h106d;
        src24 <= 16'hd83b;
        src25 <= 16'h695d;
        src26 <= 16'h4322;
        src27 <= 16'h68c4;
        src28 <= 16'had2c;
        src29 <= 16'h8006;
        src30 <= 16'hcf96;
        src31 <= 16'hc4f1;
        exp <= 21'h106a2d;
        #1
        src0 <= 16'h9d16;
        src1 <= 16'h9e58;
        src2 <= 16'h4573;
        src3 <= 16'h1a69;
        src4 <= 16'h30e7;
        src5 <= 16'h72ea;
        src6 <= 16'h6c7e;
        src7 <= 16'hc0f9;
        src8 <= 16'hd44d;
        src9 <= 16'hb539;
        src10 <= 16'hb4a6;
        src11 <= 16'hc5c4;
        src12 <= 16'hdf60;
        src13 <= 16'hfd24;
        src14 <= 16'h1273;
        src15 <= 16'hf188;
        src16 <= 16'h8e0;
        src17 <= 16'h10e9;
        src18 <= 16'h3403;
        src19 <= 16'hdf16;
        src20 <= 16'h6773;
        src21 <= 16'hda42;
        src22 <= 16'he49d;
        src23 <= 16'h1dc0;
        src24 <= 16'hfb8a;
        src25 <= 16'h36a2;
        src26 <= 16'hec17;
        src27 <= 16'hce01;
        src28 <= 16'h2f1e;
        src29 <= 16'h343a;
        src30 <= 16'h2012;
        src31 <= 16'h33f6;
        exp <= 21'h106599;
        #1
        src0 <= 16'h4270;
        src1 <= 16'he94c;
        src2 <= 16'ha0d0;
        src3 <= 16'h299;
        src4 <= 16'hb5c0;
        src5 <= 16'h23f0;
        src6 <= 16'hc73d;
        src7 <= 16'h47c8;
        src8 <= 16'h6c62;
        src9 <= 16'h473f;
        src10 <= 16'h2a18;
        src11 <= 16'he7f0;
        src12 <= 16'h3e;
        src13 <= 16'h5ecf;
        src14 <= 16'h2b37;
        src15 <= 16'h209b;
        src16 <= 16'h905c;
        src17 <= 16'hc479;
        src18 <= 16'h1a39;
        src19 <= 16'h6db0;
        src20 <= 16'h544c;
        src21 <= 16'h1a68;
        src22 <= 16'hbf06;
        src23 <= 16'hc3ab;
        src24 <= 16'h9fd6;
        src25 <= 16'hbdf0;
        src26 <= 16'h914b;
        src27 <= 16'h33da;
        src28 <= 16'h9129;
        src29 <= 16'h9d9;
        src30 <= 16'ha5b7;
        src31 <= 16'h8913;
        exp <= 21'hde33c;
        #1
        src0 <= 16'h7ead;
        src1 <= 16'ha1bf;
        src2 <= 16'hfe27;
        src3 <= 16'h9af4;
        src4 <= 16'h670a;
        src5 <= 16'hddbb;
        src6 <= 16'hb0e4;
        src7 <= 16'ha8b2;
        src8 <= 16'hbdc2;
        src9 <= 16'h171b;
        src10 <= 16'h5327;
        src11 <= 16'hdd7d;
        src12 <= 16'h2b7a;
        src13 <= 16'hd770;
        src14 <= 16'h66cb;
        src15 <= 16'hb551;
        src16 <= 16'h8733;
        src17 <= 16'h93a2;
        src18 <= 16'h3aa;
        src19 <= 16'h7eb1;
        src20 <= 16'hdbdc;
        src21 <= 16'h5c6d;
        src22 <= 16'heb9;
        src23 <= 16'h2f08;
        src24 <= 16'hedc9;
        src25 <= 16'hef31;
        src26 <= 16'h58da;
        src27 <= 16'h9be5;
        src28 <= 16'hbcf2;
        src29 <= 16'h9ad6;
        src30 <= 16'h14f7;
        src31 <= 16'hfe49;
        exp <= 21'h11cc64;
        #1
        src0 <= 16'hc2bd;
        src1 <= 16'ha402;
        src2 <= 16'h3f66;
        src3 <= 16'h217d;
        src4 <= 16'hac27;
        src5 <= 16'hd7b5;
        src6 <= 16'h2dd7;
        src7 <= 16'h3bb5;
        src8 <= 16'h7c0c;
        src9 <= 16'h1c77;
        src10 <= 16'hf82f;
        src11 <= 16'h6a2f;
        src12 <= 16'h2237;
        src13 <= 16'ha9b4;
        src14 <= 16'h6696;
        src15 <= 16'haa88;
        src16 <= 16'h518a;
        src17 <= 16'h4eff;
        src18 <= 16'h74c5;
        src19 <= 16'h1d67;
        src20 <= 16'h3715;
        src21 <= 16'ha5a9;
        src22 <= 16'h5f76;
        src23 <= 16'h3e69;
        src24 <= 16'ha49e;
        src25 <= 16'hb797;
        src26 <= 16'hbadb;
        src27 <= 16'had75;
        src28 <= 16'h2e77;
        src29 <= 16'hd804;
        src30 <= 16'h3920;
        src31 <= 16'hc939;
        exp <= 21'hf079f;
        #1
        src0 <= 16'h82e9;
        src1 <= 16'h2e4f;
        src2 <= 16'h6a68;
        src3 <= 16'hab04;
        src4 <= 16'h90ee;
        src5 <= 16'h6056;
        src6 <= 16'h771d;
        src7 <= 16'hc667;
        src8 <= 16'h14ec;
        src9 <= 16'h9774;
        src10 <= 16'h7f89;
        src11 <= 16'ha5af;
        src12 <= 16'hed5c;
        src13 <= 16'h7cea;
        src14 <= 16'h1205;
        src15 <= 16'h2036;
        src16 <= 16'h95ae;
        src17 <= 16'haa63;
        src18 <= 16'h4f80;
        src19 <= 16'hf0c;
        src20 <= 16'h9ff;
        src21 <= 16'h9f5e;
        src22 <= 16'h476e;
        src23 <= 16'h6c7;
        src24 <= 16'hb9b3;
        src25 <= 16'hb21d;
        src26 <= 16'ha2ff;
        src27 <= 16'h51ff;
        src28 <= 16'hb9d4;
        src29 <= 16'h21e9;
        src30 <= 16'he175;
        src31 <= 16'h4bd5;
        exp <= 21'he6389;
        #1
        src0 <= 16'h5adc;
        src1 <= 16'h8849;
        src2 <= 16'h76d6;
        src3 <= 16'h874;
        src4 <= 16'hc355;
        src5 <= 16'hd897;
        src6 <= 16'h289e;
        src7 <= 16'h668d;
        src8 <= 16'h126e;
        src9 <= 16'hd402;
        src10 <= 16'h2b0f;
        src11 <= 16'h1543;
        src12 <= 16'hc81;
        src13 <= 16'h8334;
        src14 <= 16'hc2de;
        src15 <= 16'h2173;
        src16 <= 16'h76fd;
        src17 <= 16'h3231;
        src18 <= 16'hdd2e;
        src19 <= 16'h3b80;
        src20 <= 16'haa9e;
        src21 <= 16'h71da;
        src22 <= 16'h732f;
        src23 <= 16'hc347;
        src24 <= 16'h5a86;
        src25 <= 16'hae7f;
        src26 <= 16'h3081;
        src27 <= 16'h397e;
        src28 <= 16'ha415;
        src29 <= 16'h3f47;
        src30 <= 16'h80ea;
        src31 <= 16'ha003;
        exp <= 21'hdb465;
        #1
        src0 <= 16'he08;
        src1 <= 16'h7226;
        src2 <= 16'h2b46;
        src3 <= 16'hd76e;
        src4 <= 16'hce7b;
        src5 <= 16'h6b09;
        src6 <= 16'h17e;
        src7 <= 16'h8270;
        src8 <= 16'hc141;
        src9 <= 16'h5121;
        src10 <= 16'h8dc;
        src11 <= 16'hb580;
        src12 <= 16'hc393;
        src13 <= 16'hf6d4;
        src14 <= 16'h5d05;
        src15 <= 16'h8c6a;
        src16 <= 16'h6941;
        src17 <= 16'hcf2;
        src18 <= 16'h76c2;
        src19 <= 16'h6051;
        src20 <= 16'hc9bb;
        src21 <= 16'h6f9c;
        src22 <= 16'ha4a0;
        src23 <= 16'h2d2c;
        src24 <= 16'h6a67;
        src25 <= 16'h8b67;
        src26 <= 16'h346;
        src27 <= 16'h39eb;
        src28 <= 16'h99a6;
        src29 <= 16'h2116;
        src30 <= 16'hed19;
        src31 <= 16'h15c2;
        exp <= 21'hdfde7;
        #1
        src0 <= 16'hdce1;
        src1 <= 16'ha2c8;
        src2 <= 16'h7d6b;
        src3 <= 16'h5e41;
        src4 <= 16'hef32;
        src5 <= 16'h7e3a;
        src6 <= 16'h8af9;
        src7 <= 16'h4039;
        src8 <= 16'hc779;
        src9 <= 16'h7953;
        src10 <= 16'h634b;
        src11 <= 16'h90a3;
        src12 <= 16'h5e48;
        src13 <= 16'h89c1;
        src14 <= 16'hfc7c;
        src15 <= 16'h647b;
        src16 <= 16'h4503;
        src17 <= 16'h4494;
        src18 <= 16'h2113;
        src19 <= 16'h6660;
        src20 <= 16'h8df7;
        src21 <= 16'h81b7;
        src22 <= 16'h9909;
        src23 <= 16'h6f23;
        src24 <= 16'h527e;
        src25 <= 16'h314b;
        src26 <= 16'h7d22;
        src27 <= 16'h2bf1;
        src28 <= 16'heef5;
        src29 <= 16'h37db;
        src30 <= 16'h6b33;
        src31 <= 16'h7233;
        exp <= 21'hf6ba3;
        #1
        src0 <= 16'h7832;
        src1 <= 16'hcba2;
        src2 <= 16'he571;
        src3 <= 16'h216c;
        src4 <= 16'h5b1d;
        src5 <= 16'he043;
        src6 <= 16'h8dcd;
        src7 <= 16'h8007;
        src8 <= 16'hc839;
        src9 <= 16'h364b;
        src10 <= 16'h124;
        src11 <= 16'ha71a;
        src12 <= 16'hd0f;
        src13 <= 16'h655e;
        src14 <= 16'h92c0;
        src15 <= 16'h4e21;
        src16 <= 16'h2778;
        src17 <= 16'hd0b8;
        src18 <= 16'h986c;
        src19 <= 16'hcc04;
        src20 <= 16'h958;
        src21 <= 16'h1cf8;
        src22 <= 16'h5e44;
        src23 <= 16'h17d;
        src24 <= 16'h2d4e;
        src25 <= 16'he066;
        src26 <= 16'hdae8;
        src27 <= 16'hf56c;
        src28 <= 16'hc997;
        src29 <= 16'hb30e;
        src30 <= 16'h7a5c;
        src31 <= 16'hc569;
        exp <= 21'h100b18;
        #1
        src0 <= 16'h4020;
        src1 <= 16'h86c7;
        src2 <= 16'h1f9d;
        src3 <= 16'h3978;
        src4 <= 16'hdfef;
        src5 <= 16'h9639;
        src6 <= 16'ha045;
        src7 <= 16'h45b2;
        src8 <= 16'hc3d7;
        src9 <= 16'hf6dc;
        src10 <= 16'he0fc;
        src11 <= 16'h81f8;
        src12 <= 16'h809f;
        src13 <= 16'h19af;
        src14 <= 16'h6c3a;
        src15 <= 16'hb720;
        src16 <= 16'h10d6;
        src17 <= 16'hc769;
        src18 <= 16'h84e2;
        src19 <= 16'h4524;
        src20 <= 16'h9443;
        src21 <= 16'h1382;
        src22 <= 16'h1383;
        src23 <= 16'hf1ce;
        src24 <= 16'h3cd5;
        src25 <= 16'h21ee;
        src26 <= 16'hb23d;
        src27 <= 16'h307a;
        src28 <= 16'h404e;
        src29 <= 16'hde09;
        src30 <= 16'h4c50;
        src31 <= 16'h7203;
        exp <= 21'hec4e9;
        #1
        src0 <= 16'h71c2;
        src1 <= 16'he9d0;
        src2 <= 16'h66fd;
        src3 <= 16'ha6eb;
        src4 <= 16'h70c9;
        src5 <= 16'h4e3e;
        src6 <= 16'h46e2;
        src7 <= 16'hcc25;
        src8 <= 16'hda39;
        src9 <= 16'h4a5d;
        src10 <= 16'h8590;
        src11 <= 16'h92fb;
        src12 <= 16'hdd2;
        src13 <= 16'h8574;
        src14 <= 16'hde89;
        src15 <= 16'hbc02;
        src16 <= 16'hc922;
        src17 <= 16'h7dcf;
        src18 <= 16'hea8d;
        src19 <= 16'hcad0;
        src20 <= 16'hb4e2;
        src21 <= 16'ha03a;
        src22 <= 16'h9fe7;
        src23 <= 16'hb477;
        src24 <= 16'h689e;
        src25 <= 16'h80e9;
        src26 <= 16'h2f3f;
        src27 <= 16'hb3cd;
        src28 <= 16'h8df1;
        src29 <= 16'h63ae;
        src30 <= 16'h6bde;
        src31 <= 16'h3196;
        exp <= 21'h11a7e8;
        #1
        src0 <= 16'hb089;
        src1 <= 16'hb5a5;
        src2 <= 16'h2af6;
        src3 <= 16'heb98;
        src4 <= 16'h3b86;
        src5 <= 16'hb36b;
        src6 <= 16'h9421;
        src7 <= 16'hf61b;
        src8 <= 16'hf8e1;
        src9 <= 16'h7d21;
        src10 <= 16'h68a1;
        src11 <= 16'ha44d;
        src12 <= 16'h8c16;
        src13 <= 16'h8590;
        src14 <= 16'h53ac;
        src15 <= 16'h9e83;
        src16 <= 16'h1172;
        src17 <= 16'h1840;
        src18 <= 16'ha0fb;
        src19 <= 16'h4a91;
        src20 <= 16'h685c;
        src21 <= 16'h2ec;
        src22 <= 16'h2a8a;
        src23 <= 16'he22b;
        src24 <= 16'hc6d3;
        src25 <= 16'h4e53;
        src26 <= 16'hbd8c;
        src27 <= 16'h115f;
        src28 <= 16'h15cd;
        src29 <= 16'h2acf;
        src30 <= 16'h3d54;
        src31 <= 16'h13a4;
        exp <= 21'he7f8e;
        #1
        src0 <= 16'hab26;
        src1 <= 16'he4c9;
        src2 <= 16'hfbe8;
        src3 <= 16'hdb35;
        src4 <= 16'h4f11;
        src5 <= 16'haf70;
        src6 <= 16'h6e5a;
        src7 <= 16'h591b;
        src8 <= 16'h7d7c;
        src9 <= 16'hc9c7;
        src10 <= 16'h1a3b;
        src11 <= 16'h5486;
        src12 <= 16'habb7;
        src13 <= 16'hf749;
        src14 <= 16'h7786;
        src15 <= 16'h7135;
        src16 <= 16'h4f0c;
        src17 <= 16'hb60c;
        src18 <= 16'h8ba7;
        src19 <= 16'hf81c;
        src20 <= 16'h55e9;
        src21 <= 16'h71ac;
        src22 <= 16'h3fdc;
        src23 <= 16'hd06e;
        src24 <= 16'hb1d9;
        src25 <= 16'hfda5;
        src26 <= 16'h3588;
        src27 <= 16'hd52a;
        src28 <= 16'h34aa;
        src29 <= 16'hab03;
        src30 <= 16'h4960;
        src31 <= 16'had41;
        exp <= 21'h125ff9;
        #1
        src0 <= 16'h9122;
        src1 <= 16'h9b56;
        src2 <= 16'hbe52;
        src3 <= 16'h7aa8;
        src4 <= 16'h6a71;
        src5 <= 16'h36dc;
        src6 <= 16'hb67c;
        src7 <= 16'hba03;
        src8 <= 16'h7d22;
        src9 <= 16'h1273;
        src10 <= 16'h83b5;
        src11 <= 16'hcefb;
        src12 <= 16'h5216;
        src13 <= 16'h5553;
        src14 <= 16'he933;
        src15 <= 16'hd267;
        src16 <= 16'h1fc7;
        src17 <= 16'hbe7b;
        src18 <= 16'haea4;
        src19 <= 16'h39ec;
        src20 <= 16'h1700;
        src21 <= 16'h473a;
        src22 <= 16'he306;
        src23 <= 16'h900d;
        src24 <= 16'h70b4;
        src25 <= 16'hcefd;
        src26 <= 16'hc140;
        src27 <= 16'hec82;
        src28 <= 16'h2f90;
        src29 <= 16'h9ebf;
        src30 <= 16'h18ae;
        src31 <= 16'h562a;
        exp <= 21'h107f3f;
        #1
        src0 <= 16'h771a;
        src1 <= 16'h3fb2;
        src2 <= 16'h6453;
        src3 <= 16'hde8f;
        src4 <= 16'hf0a1;
        src5 <= 16'h1826;
        src6 <= 16'hae21;
        src7 <= 16'hd1c1;
        src8 <= 16'h8929;
        src9 <= 16'hc1f1;
        src10 <= 16'h5a4;
        src11 <= 16'h3e66;
        src12 <= 16'hf2ea;
        src13 <= 16'h45a;
        src14 <= 16'hff65;
        src15 <= 16'h95b9;
        src16 <= 16'hccb2;
        src17 <= 16'hc4ae;
        src18 <= 16'hf687;
        src19 <= 16'h1e0;
        src20 <= 16'h584c;
        src21 <= 16'h48ae;
        src22 <= 16'h37b9;
        src23 <= 16'hb8ed;
        src24 <= 16'h52fc;
        src25 <= 16'h8ca1;
        src26 <= 16'h38e7;
        src27 <= 16'h9755;
        src28 <= 16'h445a;
        src29 <= 16'hcb65;
        src30 <= 16'hfa15;
        src31 <= 16'h9463;
        exp <= 21'h110754;
        #1
        src0 <= 16'hb289;
        src1 <= 16'hf9f6;
        src2 <= 16'ha5e7;
        src3 <= 16'hb385;
        src4 <= 16'hbd52;
        src5 <= 16'hc331;
        src6 <= 16'h1b98;
        src7 <= 16'ha84f;
        src8 <= 16'h9daf;
        src9 <= 16'h753d;
        src10 <= 16'hafba;
        src11 <= 16'hc4f0;
        src12 <= 16'h44cd;
        src13 <= 16'haf19;
        src14 <= 16'hb08b;
        src15 <= 16'h76c7;
        src16 <= 16'h34d9;
        src17 <= 16'he9f0;
        src18 <= 16'h692f;
        src19 <= 16'hc2ff;
        src20 <= 16'h417e;
        src21 <= 16'hae43;
        src22 <= 16'h453d;
        src23 <= 16'h8154;
        src24 <= 16'h20e4;
        src25 <= 16'he6f9;
        src26 <= 16'h91f3;
        src27 <= 16'h7a03;
        src28 <= 16'h8cd6;
        src29 <= 16'he237;
        src30 <= 16'hece;
        src31 <= 16'hf8a5;
        exp <= 21'h1278bf;
        #1
        src0 <= 16'h1d69;
        src1 <= 16'h697b;
        src2 <= 16'h592f;
        src3 <= 16'h5fd0;
        src4 <= 16'h801d;
        src5 <= 16'h57fd;
        src6 <= 16'he2ca;
        src7 <= 16'hcec1;
        src8 <= 16'h6728;
        src9 <= 16'hd887;
        src10 <= 16'h8632;
        src11 <= 16'h8b07;
        src12 <= 16'h1ff2;
        src13 <= 16'h7963;
        src14 <= 16'h8cea;
        src15 <= 16'h9a23;
        src16 <= 16'ha6e0;
        src17 <= 16'h8169;
        src18 <= 16'h1e42;
        src19 <= 16'h9569;
        src20 <= 16'h1f23;
        src21 <= 16'hddbc;
        src22 <= 16'hfa1f;
        src23 <= 16'h351b;
        src24 <= 16'hb365;
        src25 <= 16'h68b0;
        src26 <= 16'h6b4;
        src27 <= 16'hcb70;
        src28 <= 16'h1059;
        src29 <= 16'hd3e2;
        src30 <= 16'hb1ca;
        src31 <= 16'h8caf;
        exp <= 21'hff3cc;
        #1
        src0 <= 16'hb191;
        src1 <= 16'hc384;
        src2 <= 16'hdae0;
        src3 <= 16'h9bab;
        src4 <= 16'h4d50;
        src5 <= 16'h2064;
        src6 <= 16'h8144;
        src7 <= 16'hf3b1;
        src8 <= 16'h3e3d;
        src9 <= 16'hf341;
        src10 <= 16'h7577;
        src11 <= 16'h4bc6;
        src12 <= 16'h75e1;
        src13 <= 16'h4f62;
        src14 <= 16'hdca1;
        src15 <= 16'hf049;
        src16 <= 16'heaf0;
        src17 <= 16'h5785;
        src18 <= 16'h8ad8;
        src19 <= 16'h4e6a;
        src20 <= 16'h86ef;
        src21 <= 16'h6135;
        src22 <= 16'hdf28;
        src23 <= 16'hefd0;
        src24 <= 16'h1c2f;
        src25 <= 16'hd271;
        src26 <= 16'hc89d;
        src27 <= 16'hf171;
        src28 <= 16'hdd53;
        src29 <= 16'h2adb;
        src30 <= 16'h7d27;
        src31 <= 16'hdb15;
        exp <= 21'h132f1c;
        #1
        src0 <= 16'h8752;
        src1 <= 16'h22ce;
        src2 <= 16'hc98f;
        src3 <= 16'h9a94;
        src4 <= 16'h1e09;
        src5 <= 16'hc352;
        src6 <= 16'h66d2;
        src7 <= 16'h49c4;
        src8 <= 16'h50a7;
        src9 <= 16'hac4f;
        src10 <= 16'ha6d8;
        src11 <= 16'hcc15;
        src12 <= 16'hfceb;
        src13 <= 16'h6aeb;
        src14 <= 16'h452c;
        src15 <= 16'h1c0c;
        src16 <= 16'h6e6e;
        src17 <= 16'hf312;
        src18 <= 16'h9872;
        src19 <= 16'hc695;
        src20 <= 16'he78b;
        src21 <= 16'h1f8;
        src22 <= 16'h8228;
        src23 <= 16'h6e44;
        src24 <= 16'h40ab;
        src25 <= 16'hf02;
        src26 <= 16'h6d5b;
        src27 <= 16'hf973;
        src28 <= 16'h4822;
        src29 <= 16'h28ca;
        src30 <= 16'h25c2;
        src31 <= 16'h9c11;
        exp <= 21'hf5cd5;
        #1
        src0 <= 16'ha988;
        src1 <= 16'hf006;
        src2 <= 16'h149e;
        src3 <= 16'h74c1;
        src4 <= 16'hdd21;
        src5 <= 16'hce72;
        src6 <= 16'h8620;
        src7 <= 16'h34d1;
        src8 <= 16'hc17f;
        src9 <= 16'h48d3;
        src10 <= 16'he765;
        src11 <= 16'h351b;
        src12 <= 16'hc4ed;
        src13 <= 16'hb22b;
        src14 <= 16'h2be3;
        src15 <= 16'h9004;
        src16 <= 16'hb96d;
        src17 <= 16'h63b6;
        src18 <= 16'h79f1;
        src19 <= 16'h7a73;
        src20 <= 16'h86cd;
        src21 <= 16'hf3ef;
        src22 <= 16'hd491;
        src23 <= 16'hd40d;
        src24 <= 16'h705f;
        src25 <= 16'hb7d0;
        src26 <= 16'h6dce;
        src27 <= 16'hf7fe;
        src28 <= 16'h16fd;
        src29 <= 16'h403f;
        src30 <= 16'hd859;
        src31 <= 16'hb355;
        exp <= 21'h128908;
        #1
        src0 <= 16'h22b0;
        src1 <= 16'hf469;
        src2 <= 16'h5187;
        src3 <= 16'hf6fe;
        src4 <= 16'h4216;
        src5 <= 16'ha36c;
        src6 <= 16'hd810;
        src7 <= 16'h3883;
        src8 <= 16'ha03c;
        src9 <= 16'h7a46;
        src10 <= 16'hd00c;
        src11 <= 16'h3359;
        src12 <= 16'hb5b8;
        src13 <= 16'h1b86;
        src14 <= 16'h53ed;
        src15 <= 16'h1e8b;
        src16 <= 16'h449d;
        src17 <= 16'h589d;
        src18 <= 16'h187b;
        src19 <= 16'h6b75;
        src20 <= 16'h45fb;
        src21 <= 16'h5ab0;
        src22 <= 16'h1cc3;
        src23 <= 16'h423e;
        src24 <= 16'h1865;
        src25 <= 16'h9e84;
        src26 <= 16'he390;
        src27 <= 16'h3ffc;
        src28 <= 16'hc477;
        src29 <= 16'had03;
        src30 <= 16'hc325;
        src31 <= 16'h57ae;
        exp <= 21'he3ee8;
        #1
        src0 <= 16'h33dc;
        src1 <= 16'h17a0;
        src2 <= 16'h7;
        src3 <= 16'hecb0;
        src4 <= 16'h77ae;
        src5 <= 16'hbd21;
        src6 <= 16'hfabc;
        src7 <= 16'h697f;
        src8 <= 16'h3e61;
        src9 <= 16'h320c;
        src10 <= 16'hf285;
        src11 <= 16'h9288;
        src12 <= 16'h3463;
        src13 <= 16'ha386;
        src14 <= 16'hb26c;
        src15 <= 16'h37c;
        src16 <= 16'h3222;
        src17 <= 16'h4a72;
        src18 <= 16'ha44b;
        src19 <= 16'hd7e3;
        src20 <= 16'h789e;
        src21 <= 16'h5e65;
        src22 <= 16'hb588;
        src23 <= 16'hcd60;
        src24 <= 16'h3eed;
        src25 <= 16'h6be5;
        src26 <= 16'h169a;
        src27 <= 16'hfab7;
        src28 <= 16'h4c01;
        src29 <= 16'hb4ab;
        src30 <= 16'h10e6;
        src31 <= 16'h96d;
        exp <= 21'he7e57;
        #1
        src0 <= 16'h7435;
        src1 <= 16'h926c;
        src2 <= 16'h85c8;
        src3 <= 16'hacaa;
        src4 <= 16'h41dd;
        src5 <= 16'hcca1;
        src6 <= 16'h1e6c;
        src7 <= 16'hc9ca;
        src8 <= 16'h9889;
        src9 <= 16'h2f9a;
        src10 <= 16'h46a4;
        src11 <= 16'hb989;
        src12 <= 16'h2e67;
        src13 <= 16'hdd39;
        src14 <= 16'h2525;
        src15 <= 16'h180;
        src16 <= 16'hc16a;
        src17 <= 16'h9669;
        src18 <= 16'hd12a;
        src19 <= 16'h9b27;
        src20 <= 16'h415a;
        src21 <= 16'hd27c;
        src22 <= 16'hbf76;
        src23 <= 16'h62eb;
        src24 <= 16'h1af6;
        src25 <= 16'h7253;
        src26 <= 16'h292e;
        src27 <= 16'h4e19;
        src28 <= 16'hcf8f;
        src29 <= 16'h98cc;
        src30 <= 16'hf752;
        src31 <= 16'hc5da;
        exp <= 21'h104ece;
        #1
        src0 <= 16'h6a4d;
        src1 <= 16'h10b6;
        src2 <= 16'h87a7;
        src3 <= 16'h9fae;
        src4 <= 16'ha2a0;
        src5 <= 16'h1c;
        src6 <= 16'h45ca;
        src7 <= 16'hd4;
        src8 <= 16'ha044;
        src9 <= 16'h93ea;
        src10 <= 16'had96;
        src11 <= 16'hb5a6;
        src12 <= 16'hbe85;
        src13 <= 16'h76ca;
        src14 <= 16'h6d40;
        src15 <= 16'h9926;
        src16 <= 16'h830;
        src17 <= 16'h1d0c;
        src18 <= 16'hdd69;
        src19 <= 16'hf467;
        src20 <= 16'ha162;
        src21 <= 16'ha261;
        src22 <= 16'h205a;
        src23 <= 16'h7726;
        src24 <= 16'h5349;
        src25 <= 16'hed8a;
        src26 <= 16'h9ef7;
        src27 <= 16'h81dd;
        src28 <= 16'h7e4f;
        src29 <= 16'h8eca;
        src30 <= 16'h2e14;
        src31 <= 16'h6491;
        exp <= 21'hf3285;
        #1
        src0 <= 16'h5f33;
        src1 <= 16'hcf81;
        src2 <= 16'h1d9d;
        src3 <= 16'h92d1;
        src4 <= 16'h1f17;
        src5 <= 16'h4cbe;
        src6 <= 16'h7e27;
        src7 <= 16'h3ff1;
        src8 <= 16'h68ac;
        src9 <= 16'h45ec;
        src10 <= 16'he5e5;
        src11 <= 16'h9aba;
        src12 <= 16'h7475;
        src13 <= 16'h563a;
        src14 <= 16'hcd8b;
        src15 <= 16'h2d7f;
        src16 <= 16'h8856;
        src17 <= 16'h14da;
        src18 <= 16'h135b;
        src19 <= 16'h914e;
        src20 <= 16'h8f33;
        src21 <= 16'h74d0;
        src22 <= 16'hccfa;
        src23 <= 16'h7dac;
        src24 <= 16'he221;
        src25 <= 16'hecc0;
        src26 <= 16'h17d7;
        src27 <= 16'ha53f;
        src28 <= 16'hf6bc;
        src29 <= 16'h37af;
        src30 <= 16'h867;
        src31 <= 16'hbae8;
        exp <= 21'hf0c32;
        #1
        src0 <= 16'h68c8;
        src1 <= 16'hf352;
        src2 <= 16'hbadd;
        src3 <= 16'h3410;
        src4 <= 16'h3fb3;
        src5 <= 16'h17fd;
        src6 <= 16'h8174;
        src7 <= 16'h46ec;
        src8 <= 16'hf885;
        src9 <= 16'h18b7;
        src10 <= 16'h87dc;
        src11 <= 16'hc87b;
        src12 <= 16'he84f;
        src13 <= 16'h322b;
        src14 <= 16'hc1a5;
        src15 <= 16'hbe1a;
        src16 <= 16'h83d1;
        src17 <= 16'hb704;
        src18 <= 16'h4620;
        src19 <= 16'h9acf;
        src20 <= 16'h1280;
        src21 <= 16'had99;
        src22 <= 16'h3e24;
        src23 <= 16'h9c9d;
        src24 <= 16'h70fb;
        src25 <= 16'h9c94;
        src26 <= 16'h9cf;
        src27 <= 16'h7a7f;
        src28 <= 16'he753;
        src29 <= 16'hd80d;
        src30 <= 16'h18e8;
        src31 <= 16'h4096;
        exp <= 21'hfc83c;
        #1
        src0 <= 16'he637;
        src1 <= 16'h58c8;
        src2 <= 16'h38bd;
        src3 <= 16'h21c4;
        src4 <= 16'h5dad;
        src5 <= 16'hcbbe;
        src6 <= 16'h7926;
        src7 <= 16'hffb;
        src8 <= 16'hc7e1;
        src9 <= 16'hd47b;
        src10 <= 16'hd6b3;
        src11 <= 16'hfc84;
        src12 <= 16'h7542;
        src13 <= 16'h8900;
        src14 <= 16'h8fdd;
        src15 <= 16'hcb21;
        src16 <= 16'h9dc9;
        src17 <= 16'h94df;
        src18 <= 16'hd842;
        src19 <= 16'h4b5b;
        src20 <= 16'hf97b;
        src21 <= 16'hef21;
        src22 <= 16'hf783;
        src23 <= 16'h9b3b;
        src24 <= 16'hf68b;
        src25 <= 16'h8574;
        src26 <= 16'h2040;
        src27 <= 16'h3116;
        src28 <= 16'h8e52;
        src29 <= 16'h10d4;
        src30 <= 16'hb838;
        src31 <= 16'h3b62;
        exp <= 21'h124693;
        #1
        src0 <= 16'hefb;
        src1 <= 16'h5c8a;
        src2 <= 16'h33b6;
        src3 <= 16'hae7d;
        src4 <= 16'hdd70;
        src5 <= 16'h5cf6;
        src6 <= 16'h9f6f;
        src7 <= 16'h8302;
        src8 <= 16'h6289;
        src9 <= 16'h9eb4;
        src10 <= 16'he8b5;
        src11 <= 16'h415;
        src12 <= 16'h57ec;
        src13 <= 16'hfd1c;
        src14 <= 16'hccd;
        src15 <= 16'ha771;
        src16 <= 16'hbec5;
        src17 <= 16'hfe7f;
        src18 <= 16'h87d;
        src19 <= 16'h611a;
        src20 <= 16'h4b50;
        src21 <= 16'h321c;
        src22 <= 16'h32a5;
        src23 <= 16'hf15c;
        src24 <= 16'hc667;
        src25 <= 16'h3b4;
        src26 <= 16'hdb91;
        src27 <= 16'ha845;
        src28 <= 16'h2b6d;
        src29 <= 16'he281;
        src30 <= 16'h1b00;
        src31 <= 16'h2e4b;
        exp <= 21'hf0f4e;
        #1
        src0 <= 16'hef7;
        src1 <= 16'h4863;
        src2 <= 16'he734;
        src3 <= 16'h376d;
        src4 <= 16'h8f17;
        src5 <= 16'hec84;
        src6 <= 16'hd23d;
        src7 <= 16'he737;
        src8 <= 16'hf11d;
        src9 <= 16'h4fe6;
        src10 <= 16'he1b1;
        src11 <= 16'h578a;
        src12 <= 16'h547c;
        src13 <= 16'ha5e4;
        src14 <= 16'h1498;
        src15 <= 16'h59ad;
        src16 <= 16'ha644;
        src17 <= 16'hc29d;
        src18 <= 16'hd04d;
        src19 <= 16'h71fe;
        src20 <= 16'he17;
        src21 <= 16'h667e;
        src22 <= 16'haae3;
        src23 <= 16'h21b1;
        src24 <= 16'hccbb;
        src25 <= 16'h2724;
        src26 <= 16'hedd;
        src27 <= 16'h3261;
        src28 <= 16'hffc3;
        src29 <= 16'hb36c;
        src30 <= 16'hcfe1;
        src31 <= 16'hbd72;
        exp <= 21'h10efe1;
        #1
        src0 <= 16'h1306;
        src1 <= 16'h16ab;
        src2 <= 16'h8fe6;
        src3 <= 16'h23cb;
        src4 <= 16'h6d3f;
        src5 <= 16'h8a3d;
        src6 <= 16'h6b95;
        src7 <= 16'hfbfd;
        src8 <= 16'he710;
        src9 <= 16'h196c;
        src10 <= 16'h57a9;
        src11 <= 16'hd492;
        src12 <= 16'h8c0e;
        src13 <= 16'h606a;
        src14 <= 16'hff09;
        src15 <= 16'hbd92;
        src16 <= 16'hebf3;
        src17 <= 16'hcf4f;
        src18 <= 16'h3415;
        src19 <= 16'hcad1;
        src20 <= 16'h6ad7;
        src21 <= 16'hdc0;
        src22 <= 16'hf24a;
        src23 <= 16'hf92c;
        src24 <= 16'h5cb9;
        src25 <= 16'h939b;
        src26 <= 16'h86;
        src27 <= 16'h2e23;
        src28 <= 16'h16b9;
        src29 <= 16'hec80;
        src30 <= 16'h22d0;
        src31 <= 16'hc572;
        exp <= 21'h103ae7;
        #1
        src0 <= 16'h2920;
        src1 <= 16'h1a88;
        src2 <= 16'hd2b6;
        src3 <= 16'hffc4;
        src4 <= 16'hb62a;
        src5 <= 16'h7fb;
        src6 <= 16'h6435;
        src7 <= 16'ha8d;
        src8 <= 16'hf24f;
        src9 <= 16'h20fd;
        src10 <= 16'hd594;
        src11 <= 16'hbf4;
        src12 <= 16'hdc98;
        src13 <= 16'h79ed;
        src14 <= 16'ha34d;
        src15 <= 16'hfbf7;
        src16 <= 16'hb0a6;
        src17 <= 16'h8c21;
        src18 <= 16'hbde7;
        src19 <= 16'hce20;
        src20 <= 16'h782f;
        src21 <= 16'h348c;
        src22 <= 16'h7bea;
        src23 <= 16'ha1cd;
        src24 <= 16'h3d70;
        src25 <= 16'h363;
        src26 <= 16'hda4c;
        src27 <= 16'h655a;
        src28 <= 16'h392b;
        src29 <= 16'h88ca;
        src30 <= 16'h9b7f;
        src31 <= 16'hdaa6;
        exp <= 21'h107979;
        #1
        src0 <= 16'hfe1a;
        src1 <= 16'hf6d6;
        src2 <= 16'h8881;
        src3 <= 16'h5e6d;
        src4 <= 16'hdccc;
        src5 <= 16'hf8ba;
        src6 <= 16'he5a9;
        src7 <= 16'ha95f;
        src8 <= 16'ha2fb;
        src9 <= 16'h50db;
        src10 <= 16'h3ab;
        src11 <= 16'hd914;
        src12 <= 16'hd04f;
        src13 <= 16'haeb8;
        src14 <= 16'ha1eb;
        src15 <= 16'h5c45;
        src16 <= 16'hd043;
        src17 <= 16'he6d5;
        src18 <= 16'h5f9;
        src19 <= 16'hf82;
        src20 <= 16'h1a70;
        src21 <= 16'he15b;
        src22 <= 16'h9b1d;
        src23 <= 16'hb190;
        src24 <= 16'haa7f;
        src25 <= 16'hd08;
        src26 <= 16'h649;
        src27 <= 16'hc0ac;
        src28 <= 16'h3b92;
        src29 <= 16'h3af2;
        src30 <= 16'hc809;
        src31 <= 16'h91c2;
        exp <= 21'h11f20e;
        #1
        src0 <= 16'hb135;
        src1 <= 16'hd9a1;
        src2 <= 16'h895b;
        src3 <= 16'h7589;
        src4 <= 16'h25c3;
        src5 <= 16'hf09c;
        src6 <= 16'h2e6d;
        src7 <= 16'h272c;
        src8 <= 16'hadf8;
        src9 <= 16'h863a;
        src10 <= 16'hcd03;
        src11 <= 16'h903;
        src12 <= 16'h2841;
        src13 <= 16'hca17;
        src14 <= 16'h2337;
        src15 <= 16'hc96d;
        src16 <= 16'ha304;
        src17 <= 16'h1eb2;
        src18 <= 16'h55be;
        src19 <= 16'he561;
        src20 <= 16'h9b92;
        src21 <= 16'h5ba5;
        src22 <= 16'hbe13;
        src23 <= 16'he588;
        src24 <= 16'hc2a4;
        src25 <= 16'h7a04;
        src26 <= 16'hc98e;
        src27 <= 16'hcdea;
        src28 <= 16'h172f;
        src29 <= 16'h6957;
        src30 <= 16'hb31;
        src31 <= 16'h23f0;
        exp <= 21'hffa54;
        #1
        src0 <= 16'ha853;
        src1 <= 16'h3ec5;
        src2 <= 16'h8107;
        src3 <= 16'hea77;
        src4 <= 16'hb166;
        src5 <= 16'h188;
        src6 <= 16'h771f;
        src7 <= 16'h3cb6;
        src8 <= 16'had42;
        src9 <= 16'h4a69;
        src10 <= 16'h27d3;
        src11 <= 16'hc470;
        src12 <= 16'hbbcd;
        src13 <= 16'h98b;
        src14 <= 16'h448d;
        src15 <= 16'ha39d;
        src16 <= 16'h8e9d;
        src17 <= 16'hef51;
        src18 <= 16'h70ef;
        src19 <= 16'h79e0;
        src20 <= 16'hda59;
        src21 <= 16'h82a3;
        src22 <= 16'h8317;
        src23 <= 16'h4187;
        src24 <= 16'h5be6;
        src25 <= 16'h1351;
        src26 <= 16'h2805;
        src27 <= 16'h1515;
        src28 <= 16'hf8f4;
        src29 <= 16'h9e2b;
        src30 <= 16'h62a8;
        src31 <= 16'h7f74;
        exp <= 21'hefaac;
        #1
        src0 <= 16'h49d9;
        src1 <= 16'hc399;
        src2 <= 16'h338e;
        src3 <= 16'h80f1;
        src4 <= 16'h3e2c;
        src5 <= 16'h15ad;
        src6 <= 16'h5d84;
        src7 <= 16'hfd04;
        src8 <= 16'h73d7;
        src9 <= 16'hd88b;
        src10 <= 16'hb9fe;
        src11 <= 16'h8fef;
        src12 <= 16'hf0a5;
        src13 <= 16'h460;
        src14 <= 16'h719d;
        src15 <= 16'habcf;
        src16 <= 16'ha2cb;
        src17 <= 16'h5b09;
        src18 <= 16'h5d1;
        src19 <= 16'h14a1;
        src20 <= 16'hdee;
        src21 <= 16'h9b06;
        src22 <= 16'hf7d3;
        src23 <= 16'h72a8;
        src24 <= 16'haa68;
        src25 <= 16'h725f;
        src26 <= 16'h28aa;
        src27 <= 16'h3663;
        src28 <= 16'he60c;
        src29 <= 16'hd68a;
        src30 <= 16'ha25c;
        src31 <= 16'h2b36;
        exp <= 21'hf4ac3;
        #1
        src0 <= 16'ha45e;
        src1 <= 16'hc140;
        src2 <= 16'h71d0;
        src3 <= 16'hd5c3;
        src4 <= 16'h54d2;
        src5 <= 16'h74d;
        src6 <= 16'hafd1;
        src7 <= 16'hce52;
        src8 <= 16'hbd8;
        src9 <= 16'ha669;
        src10 <= 16'hf7f;
        src11 <= 16'h63a7;
        src12 <= 16'h484c;
        src13 <= 16'hf6bd;
        src14 <= 16'ha3cb;
        src15 <= 16'h7629;
        src16 <= 16'hd083;
        src17 <= 16'h5e7e;
        src18 <= 16'hf52;
        src19 <= 16'hb32;
        src20 <= 16'h4f64;
        src21 <= 16'hd70d;
        src22 <= 16'h7cdd;
        src23 <= 16'h1781;
        src24 <= 16'h16b8;
        src25 <= 16'h1d5b;
        src26 <= 16'hb7d4;
        src27 <= 16'h1457;
        src28 <= 16'ha9b8;
        src29 <= 16'h20b2;
        src30 <= 16'h6136;
        src31 <= 16'h9487;
        exp <= 21'hdca90;
        #1
        src0 <= 16'he74e;
        src1 <= 16'h553f;
        src2 <= 16'h6205;
        src3 <= 16'he895;
        src4 <= 16'h25ec;
        src5 <= 16'hf397;
        src6 <= 16'h5eea;
        src7 <= 16'h3646;
        src8 <= 16'h2b75;
        src9 <= 16'h8a88;
        src10 <= 16'hddf7;
        src11 <= 16'h7a44;
        src12 <= 16'h284a;
        src13 <= 16'h8e7a;
        src14 <= 16'hbf4e;
        src15 <= 16'h1d7a;
        src16 <= 16'h5883;
        src17 <= 16'hf1fe;
        src18 <= 16'h1ea5;
        src19 <= 16'h88a6;
        src20 <= 16'hdaef;
        src21 <= 16'h3f6a;
        src22 <= 16'h5522;
        src23 <= 16'hd7f8;
        src24 <= 16'hab15;
        src25 <= 16'hd0e8;
        src26 <= 16'hf59a;
        src27 <= 16'hda08;
        src28 <= 16'hecb7;
        src29 <= 16'he7a9;
        src30 <= 16'he63a;
        src31 <= 16'h9938;
        exp <= 21'h12b04e;
        #1
        src0 <= 16'h2486;
        src1 <= 16'h74f6;
        src2 <= 16'h9b9a;
        src3 <= 16'h74de;
        src4 <= 16'h3bd0;
        src5 <= 16'hdac6;
        src6 <= 16'h3178;
        src7 <= 16'h1d14;
        src8 <= 16'h4b8d;
        src9 <= 16'h5fa6;
        src10 <= 16'h7b01;
        src11 <= 16'h866d;
        src12 <= 16'h4867;
        src13 <= 16'hace1;
        src14 <= 16'h1c53;
        src15 <= 16'hecc9;
        src16 <= 16'hfa23;
        src17 <= 16'he6f2;
        src18 <= 16'hb86a;
        src19 <= 16'hf94d;
        src20 <= 16'hd6d8;
        src21 <= 16'h91fe;
        src22 <= 16'h3b0d;
        src23 <= 16'he0c0;
        src24 <= 16'h8755;
        src25 <= 16'h69f6;
        src26 <= 16'hac0;
        src27 <= 16'ha3da;
        src28 <= 16'h1560;
        src29 <= 16'hcef7;
        src30 <= 16'h4fde;
        src31 <= 16'h4162;
        exp <= 21'hfe706;
        #1
        src0 <= 16'h6f29;
        src1 <= 16'h1545;
        src2 <= 16'h725f;
        src3 <= 16'h8913;
        src4 <= 16'h9809;
        src5 <= 16'hb31b;
        src6 <= 16'h5164;
        src7 <= 16'h5f46;
        src8 <= 16'h18b3;
        src9 <= 16'h8480;
        src10 <= 16'h1a26;
        src11 <= 16'h5280;
        src12 <= 16'hc89d;
        src13 <= 16'h7ec1;
        src14 <= 16'hf424;
        src15 <= 16'h7f43;
        src16 <= 16'h87ce;
        src17 <= 16'h7db3;
        src18 <= 16'h51a;
        src19 <= 16'hb2d2;
        src20 <= 16'hf6fc;
        src21 <= 16'h4124;
        src22 <= 16'haeaa;
        src23 <= 16'hba33;
        src24 <= 16'h63c6;
        src25 <= 16'h318f;
        src26 <= 16'h68e2;
        src27 <= 16'h6e84;
        src28 <= 16'h12ab;
        src29 <= 16'hba39;
        src30 <= 16'h8a5c;
        src31 <= 16'h26b7;
        exp <= 21'he8968;
        #1
        src0 <= 16'h4554;
        src1 <= 16'he138;
        src2 <= 16'hd133;
        src3 <= 16'h17b5;
        src4 <= 16'he4af;
        src5 <= 16'hc07f;
        src6 <= 16'h2328;
        src7 <= 16'hc83d;
        src8 <= 16'h92;
        src9 <= 16'hc422;
        src10 <= 16'h2441;
        src11 <= 16'h1c7e;
        src12 <= 16'hc8ab;
        src13 <= 16'h99cc;
        src14 <= 16'h6b27;
        src15 <= 16'h5468;
        src16 <= 16'h9547;
        src17 <= 16'h2655;
        src18 <= 16'h80b8;
        src19 <= 16'hda4;
        src20 <= 16'h7129;
        src21 <= 16'h20eb;
        src22 <= 16'h2def;
        src23 <= 16'h9912;
        src24 <= 16'h2003;
        src25 <= 16'hfe39;
        src26 <= 16'h78a2;
        src27 <= 16'h6408;
        src28 <= 16'hb69;
        src29 <= 16'h1dd7;
        src30 <= 16'hf285;
        src31 <= 16'h6b6e;
        exp <= 21'hdeca6;
        #1
        src0 <= 16'hd994;
        src1 <= 16'h6395;
        src2 <= 16'hcc0;
        src3 <= 16'h6505;
        src4 <= 16'hda7d;
        src5 <= 16'h4b97;
        src6 <= 16'h3c;
        src7 <= 16'h3301;
        src8 <= 16'ha365;
        src9 <= 16'h5353;
        src10 <= 16'h3f2;
        src11 <= 16'hc25d;
        src12 <= 16'hfa33;
        src13 <= 16'h9c75;
        src14 <= 16'h9e74;
        src15 <= 16'h553e;
        src16 <= 16'h21a7;
        src17 <= 16'ha0bd;
        src18 <= 16'h5e3a;
        src19 <= 16'h372f;
        src20 <= 16'he2a3;
        src21 <= 16'he06;
        src22 <= 16'h851b;
        src23 <= 16'h29c6;
        src24 <= 16'h75fa;
        src25 <= 16'hf3cf;
        src26 <= 16'h544a;
        src27 <= 16'h2320;
        src28 <= 16'hbffc;
        src29 <= 16'h64ba;
        src30 <= 16'he997;
        src31 <= 16'hc1ec;
        exp <= 21'hef863;
        #1
        src0 <= 16'ha5d8;
        src1 <= 16'h95e1;
        src2 <= 16'h4945;
        src3 <= 16'h2573;
        src4 <= 16'h3d31;
        src5 <= 16'h3636;
        src6 <= 16'hba61;
        src7 <= 16'h260d;
        src8 <= 16'h213a;
        src9 <= 16'hc679;
        src10 <= 16'h94d2;
        src11 <= 16'h965c;
        src12 <= 16'hf07e;
        src13 <= 16'h7922;
        src14 <= 16'h1a1c;
        src15 <= 16'h9273;
        src16 <= 16'h2777;
        src17 <= 16'hf3aa;
        src18 <= 16'he1cc;
        src19 <= 16'hbe1b;
        src20 <= 16'h3af6;
        src21 <= 16'ha239;
        src22 <= 16'h820;
        src23 <= 16'h2bff;
        src24 <= 16'hca13;
        src25 <= 16'ha22d;
        src26 <= 16'hbd87;
        src27 <= 16'h65a2;
        src28 <= 16'h2ae1;
        src29 <= 16'he256;
        src30 <= 16'hb204;
        src31 <= 16'hf42;
        exp <= 21'hf5192;
        #1
        src0 <= 16'h6be9;
        src1 <= 16'hcaab;
        src2 <= 16'h78e1;
        src3 <= 16'he991;
        src4 <= 16'he87c;
        src5 <= 16'hb954;
        src6 <= 16'hd556;
        src7 <= 16'h240e;
        src8 <= 16'h8562;
        src9 <= 16'hc0bd;
        src10 <= 16'hc0f6;
        src11 <= 16'hec75;
        src12 <= 16'h49d5;
        src13 <= 16'heebb;
        src14 <= 16'h6cf0;
        src15 <= 16'he242;
        src16 <= 16'h7e4c;
        src17 <= 16'hfb65;
        src18 <= 16'ha632;
        src19 <= 16'h30e4;
        src20 <= 16'hd83d;
        src21 <= 16'h7ce3;
        src22 <= 16'hc4f0;
        src23 <= 16'h3d06;
        src24 <= 16'hd790;
        src25 <= 16'h99be;
        src26 <= 16'h8b09;
        src27 <= 16'h9e1d;
        src28 <= 16'hb1bf;
        src29 <= 16'hae2;
        src30 <= 16'h5148;
        src31 <= 16'h5781;
        exp <= 21'h135741;
        #1
        src0 <= 16'ha56e;
        src1 <= 16'h8e70;
        src2 <= 16'hdbb6;
        src3 <= 16'h5719;
        src4 <= 16'ha07f;
        src5 <= 16'hbccd;
        src6 <= 16'hb69a;
        src7 <= 16'h2833;
        src8 <= 16'hfb87;
        src9 <= 16'h7c6a;
        src10 <= 16'h132;
        src11 <= 16'h7c53;
        src12 <= 16'h89ca;
        src13 <= 16'hf2a8;
        src14 <= 16'hce76;
        src15 <= 16'h2ccf;
        src16 <= 16'hcdd8;
        src17 <= 16'h8b1e;
        src18 <= 16'hed85;
        src19 <= 16'h9ba7;
        src20 <= 16'h3c9f;
        src21 <= 16'hb058;
        src22 <= 16'ha725;
        src23 <= 16'hf852;
        src24 <= 16'hbab2;
        src25 <= 16'h4658;
        src26 <= 16'hb280;
        src27 <= 16'h943a;
        src28 <= 16'h8290;
        src29 <= 16'he8f9;
        src30 <= 16'h3f4c;
        src31 <= 16'h2f61;
        exp <= 21'h12a07d;
        #1
        src0 <= 16'h4833;
        src1 <= 16'hb870;
        src2 <= 16'h276b;
        src3 <= 16'h9ca3;
        src4 <= 16'h91c4;
        src5 <= 16'h5558;
        src6 <= 16'h3053;
        src7 <= 16'h7326;
        src8 <= 16'h1107;
        src9 <= 16'h1124;
        src10 <= 16'h47fa;
        src11 <= 16'h9855;
        src12 <= 16'h72aa;
        src13 <= 16'h6b74;
        src14 <= 16'h4a0e;
        src15 <= 16'h52dd;
        src16 <= 16'h2593;
        src17 <= 16'h42fe;
        src18 <= 16'h786;
        src19 <= 16'h3efc;
        src20 <= 16'h6006;
        src21 <= 16'h71d7;
        src22 <= 16'hfa7e;
        src23 <= 16'hf6cf;
        src24 <= 16'h30f0;
        src25 <= 16'h9832;
        src26 <= 16'hb824;
        src27 <= 16'h52ce;
        src28 <= 16'h6e7f;
        src29 <= 16'h81d;
        src30 <= 16'h2fec;
        src31 <= 16'h5c67;
        exp <= 21'hc1609;
        #1
        src0 <= 16'h8ab9;
        src1 <= 16'h2ef9;
        src2 <= 16'h4218;
        src3 <= 16'hca8a;
        src4 <= 16'h3c0c;
        src5 <= 16'he4d7;
        src6 <= 16'h74c4;
        src7 <= 16'h25bf;
        src8 <= 16'h5066;
        src9 <= 16'h36a1;
        src10 <= 16'hc1dc;
        src11 <= 16'h7658;
        src12 <= 16'hf6ff;
        src13 <= 16'hc26c;
        src14 <= 16'h5abd;
        src15 <= 16'h33f;
        src16 <= 16'h2c63;
        src17 <= 16'hd91f;
        src18 <= 16'hf0c4;
        src19 <= 16'he6ef;
        src20 <= 16'h2a86;
        src21 <= 16'he32d;
        src22 <= 16'h519a;
        src23 <= 16'ha7f3;
        src24 <= 16'hedd;
        src25 <= 16'h9468;
        src26 <= 16'h30a9;
        src27 <= 16'h80c9;
        src28 <= 16'h1579;
        src29 <= 16'ha210;
        src30 <= 16'h5855;
        src31 <= 16'hec42;
        exp <= 21'hf8da8;
        #1
        src0 <= 16'hb1fc;
        src1 <= 16'h83ff;
        src2 <= 16'hbfe5;
        src3 <= 16'hbfcb;
        src4 <= 16'hc78f;
        src5 <= 16'hd4a8;
        src6 <= 16'h330e;
        src7 <= 16'h4501;
        src8 <= 16'h355b;
        src9 <= 16'h716b;
        src10 <= 16'hef0e;
        src11 <= 16'hec3b;
        src12 <= 16'hf335;
        src13 <= 16'hdc11;
        src14 <= 16'hbf12;
        src15 <= 16'hfe4e;
        src16 <= 16'h2c7c;
        src17 <= 16'hc1bb;
        src18 <= 16'hfd9d;
        src19 <= 16'h15bf;
        src20 <= 16'h785;
        src21 <= 16'h7591;
        src22 <= 16'h5bf6;
        src23 <= 16'hbb05;
        src24 <= 16'hf50f;
        src25 <= 16'h2e90;
        src26 <= 16'h482d;
        src27 <= 16'hc0a2;
        src28 <= 16'hcf42;
        src29 <= 16'h13e3;
        src30 <= 16'h158f;
        src31 <= 16'hf93c;
        exp <= 21'h128ca8;
        #1
        src0 <= 16'h4001;
        src1 <= 16'h7dd2;
        src2 <= 16'hd29b;
        src3 <= 16'h55b5;
        src4 <= 16'hb0e4;
        src5 <= 16'hcd3;
        src6 <= 16'hf9e4;
        src7 <= 16'h20c0;
        src8 <= 16'hc238;
        src9 <= 16'h4c19;
        src10 <= 16'h29c2;
        src11 <= 16'h2807;
        src12 <= 16'h6b69;
        src13 <= 16'hbaee;
        src14 <= 16'h8198;
        src15 <= 16'h70cc;
        src16 <= 16'h22cd;
        src17 <= 16'h54b3;
        src18 <= 16'h7927;
        src19 <= 16'he27b;
        src20 <= 16'h835c;
        src21 <= 16'h4a25;
        src22 <= 16'hc283;
        src23 <= 16'h9b4b;
        src24 <= 16'h7aee;
        src25 <= 16'h90c7;
        src26 <= 16'hc8fb;
        src27 <= 16'hd8be;
        src28 <= 16'h3d0d;
        src29 <= 16'h3fe5;
        src30 <= 16'hb797;
        src31 <= 16'h8439;
        exp <= 21'hf9bf4;
        #1
        src0 <= 16'h2201;
        src1 <= 16'ha3d4;
        src2 <= 16'h900c;
        src3 <= 16'h994e;
        src4 <= 16'h1937;
        src5 <= 16'h8897;
        src6 <= 16'hf331;
        src7 <= 16'h9084;
        src8 <= 16'ha842;
        src9 <= 16'hecc7;
        src10 <= 16'hf7aa;
        src11 <= 16'h403;
        src12 <= 16'hfcbf;
        src13 <= 16'h24c1;
        src14 <= 16'h9571;
        src15 <= 16'h3468;
        src16 <= 16'hcb84;
        src17 <= 16'hb46c;
        src18 <= 16'ha084;
        src19 <= 16'he3b1;
        src20 <= 16'h72cb;
        src21 <= 16'hc5ae;
        src22 <= 16'haf86;
        src23 <= 16'hff6c;
        src24 <= 16'h5fc0;
        src25 <= 16'h8a92;
        src26 <= 16'h6878;
        src27 <= 16'h9604;
        src28 <= 16'h7f08;
        src29 <= 16'hf963;
        src30 <= 16'hd8b8;
        src31 <= 16'h8fd1;
        exp <= 21'h134613;
        #1
        src0 <= 16'hab11;
        src1 <= 16'h9a79;
        src2 <= 16'hb59c;
        src3 <= 16'h3764;
        src4 <= 16'hbe4;
        src5 <= 16'hdac;
        src6 <= 16'hc08d;
        src7 <= 16'h766f;
        src8 <= 16'hc2e3;
        src9 <= 16'hfb0d;
        src10 <= 16'hb137;
        src11 <= 16'h2649;
        src12 <= 16'h3231;
        src13 <= 16'h50e6;
        src14 <= 16'h7ec0;
        src15 <= 16'h7f9;
        src16 <= 16'h8f00;
        src17 <= 16'hb4fe;
        src18 <= 16'hfb10;
        src19 <= 16'h8d9c;
        src20 <= 16'h524a;
        src21 <= 16'h5509;
        src22 <= 16'h8405;
        src23 <= 16'hf651;
        src24 <= 16'h6f0d;
        src25 <= 16'hea3;
        src26 <= 16'h5f10;
        src27 <= 16'h43c0;
        src28 <= 16'h724c;
        src29 <= 16'h149a;
        src30 <= 16'h418a;
        src31 <= 16'h9b0b;
        exp <= 21'he94a4;
        #1
        src0 <= 16'h41ac;
        src1 <= 16'h2992;
        src2 <= 16'haba4;
        src3 <= 16'h19fd;
        src4 <= 16'h8238;
        src5 <= 16'h1f16;
        src6 <= 16'hade0;
        src7 <= 16'h8a1;
        src8 <= 16'h1b6;
        src9 <= 16'h8c9e;
        src10 <= 16'hc9a8;
        src11 <= 16'hf075;
        src12 <= 16'hd8a0;
        src13 <= 16'h918d;
        src14 <= 16'hb1d9;
        src15 <= 16'h3da0;
        src16 <= 16'h7048;
        src17 <= 16'h8a02;
        src18 <= 16'hb423;
        src19 <= 16'h5a34;
        src20 <= 16'h5f88;
        src21 <= 16'hd371;
        src22 <= 16'h8012;
        src23 <= 16'had60;
        src24 <= 16'hca06;
        src25 <= 16'h8530;
        src26 <= 16'h4b18;
        src27 <= 16'h78e3;
        src28 <= 16'h3dab;
        src29 <= 16'he2d2;
        src30 <= 16'he1de;
        src31 <= 16'h57d5;
        exp <= 21'h100132;
        #1
        src0 <= 16'h89b3;
        src1 <= 16'h7f7f;
        src2 <= 16'h8299;
        src3 <= 16'h66a2;
        src4 <= 16'hf125;
        src5 <= 16'h84ec;
        src6 <= 16'h67e8;
        src7 <= 16'h7a04;
        src8 <= 16'ha71;
        src9 <= 16'hc83;
        src10 <= 16'hf48f;
        src11 <= 16'ha12e;
        src12 <= 16'hd8cf;
        src13 <= 16'h4b01;
        src14 <= 16'hbd35;
        src15 <= 16'h6960;
        src16 <= 16'h9ff6;
        src17 <= 16'h461c;
        src18 <= 16'hca2e;
        src19 <= 16'h952b;
        src20 <= 16'h6c02;
        src21 <= 16'h6fa1;
        src22 <= 16'he14d;
        src23 <= 16'h53f9;
        src24 <= 16'h7db8;
        src25 <= 16'h7b9b;
        src26 <= 16'h37aa;
        src27 <= 16'h41e1;
        src28 <= 16'h9185;
        src29 <= 16'ha741;
        src30 <= 16'h266d;
        src31 <= 16'hefba;
        exp <= 21'h10599f;
        #1
        src0 <= 16'h9e3a;
        src1 <= 16'hfd8f;
        src2 <= 16'hb444;
        src3 <= 16'h472d;
        src4 <= 16'h4892;
        src5 <= 16'h3865;
        src6 <= 16'hdc55;
        src7 <= 16'h3fe9;
        src8 <= 16'h6a92;
        src9 <= 16'h7d1a;
        src10 <= 16'h4736;
        src11 <= 16'ha130;
        src12 <= 16'hf9b3;
        src13 <= 16'h4b47;
        src14 <= 16'hd509;
        src15 <= 16'h84ea;
        src16 <= 16'hcd12;
        src17 <= 16'hb962;
        src18 <= 16'h2b22;
        src19 <= 16'hd67a;
        src20 <= 16'h84c1;
        src21 <= 16'hd4db;
        src22 <= 16'h6931;
        src23 <= 16'h217d;
        src24 <= 16'ha911;
        src25 <= 16'hb8a2;
        src26 <= 16'h896f;
        src27 <= 16'hb224;
        src28 <= 16'h2764;
        src29 <= 16'h233a;
        src30 <= 16'hc28b;
        src31 <= 16'hb661;
        exp <= 21'h117098;
        #1
        src0 <= 16'h7f78;
        src1 <= 16'h1b0d;
        src2 <= 16'h83a1;
        src3 <= 16'h255a;
        src4 <= 16'h9c3d;
        src5 <= 16'ha0c7;
        src6 <= 16'h7d1e;
        src7 <= 16'hb724;
        src8 <= 16'heefe;
        src9 <= 16'haa06;
        src10 <= 16'h7da0;
        src11 <= 16'hbf3a;
        src12 <= 16'he41c;
        src13 <= 16'h2b65;
        src14 <= 16'h64f2;
        src15 <= 16'hdf97;
        src16 <= 16'hac3d;
        src17 <= 16'hcf94;
        src18 <= 16'h68f2;
        src19 <= 16'hbb9f;
        src20 <= 16'h71e3;
        src21 <= 16'hfdaa;
        src22 <= 16'h4636;
        src23 <= 16'h4ed6;
        src24 <= 16'hffd7;
        src25 <= 16'hbaa4;
        src26 <= 16'h4f6e;
        src27 <= 16'h96c;
        src28 <= 16'h823f;
        src29 <= 16'h4e3;
        src30 <= 16'h8e15;
        src31 <= 16'hb049;
        exp <= 21'h115c7e;
        #1
        src0 <= 16'h675a;
        src1 <= 16'h2ef;
        src2 <= 16'hc6d5;
        src3 <= 16'h9a96;
        src4 <= 16'h4424;
        src5 <= 16'he3b0;
        src6 <= 16'hca39;
        src7 <= 16'h4cb1;
        src8 <= 16'h616b;
        src9 <= 16'h6538;
        src10 <= 16'h76ed;
        src11 <= 16'hc48c;
        src12 <= 16'hded4;
        src13 <= 16'he14e;
        src14 <= 16'hb3e1;
        src15 <= 16'h3db5;
        src16 <= 16'hb6a1;
        src17 <= 16'hd3ef;
        src18 <= 16'h86c7;
        src19 <= 16'h6959;
        src20 <= 16'hd612;
        src21 <= 16'h3387;
        src22 <= 16'h4566;
        src23 <= 16'hbc7d;
        src24 <= 16'h6be2;
        src25 <= 16'h9874;
        src26 <= 16'ha23d;
        src27 <= 16'hef2b;
        src28 <= 16'h36;
        src29 <= 16'h6121;
        src30 <= 16'ha570;
        src31 <= 16'hc68b;
        exp <= 21'h11a782;
        #1
        src0 <= 16'h2776;
        src1 <= 16'h4cd0;
        src2 <= 16'h9876;
        src3 <= 16'h7d14;
        src4 <= 16'h7271;
        src5 <= 16'h344a;
        src6 <= 16'hbfb8;
        src7 <= 16'he2f6;
        src8 <= 16'h8c66;
        src9 <= 16'hcffe;
        src10 <= 16'hc620;
        src11 <= 16'h78b2;
        src12 <= 16'hf47e;
        src13 <= 16'hbe9;
        src14 <= 16'hf82f;
        src15 <= 16'hbaa4;
        src16 <= 16'h8fc4;
        src17 <= 16'h56a7;
        src18 <= 16'h6745;
        src19 <= 16'h3043;
        src20 <= 16'h9a40;
        src21 <= 16'ha81e;
        src22 <= 16'h395d;
        src23 <= 16'hc7d6;
        src24 <= 16'hb71b;
        src25 <= 16'ha5bb;
        src26 <= 16'hca5d;
        src27 <= 16'h8ae1;
        src28 <= 16'ha45a;
        src29 <= 16'hba11;
        src30 <= 16'h8691;
        src31 <= 16'h8c47;
        exp <= 21'h120684;
        #1
        src0 <= 16'h280d;
        src1 <= 16'h6941;
        src2 <= 16'h5b2;
        src3 <= 16'hc81a;
        src4 <= 16'h71cd;
        src5 <= 16'h69fc;
        src6 <= 16'hcb7b;
        src7 <= 16'hd138;
        src8 <= 16'h35d6;
        src9 <= 16'h311f;
        src10 <= 16'hc9d;
        src11 <= 16'h7988;
        src12 <= 16'hb93c;
        src13 <= 16'h2c79;
        src14 <= 16'h7d1e;
        src15 <= 16'h488;
        src16 <= 16'hcdd2;
        src17 <= 16'ha9c6;
        src18 <= 16'hbab6;
        src19 <= 16'hb610;
        src20 <= 16'he5ba;
        src21 <= 16'h7e82;
        src22 <= 16'h1fb2;
        src23 <= 16'h37d4;
        src24 <= 16'h3d2d;
        src25 <= 16'hb5a1;
        src26 <= 16'h9212;
        src27 <= 16'hf80e;
        src28 <= 16'h4a17;
        src29 <= 16'h32f5;
        src30 <= 16'h1ce8;
        src31 <= 16'hc4c5;
        exp <= 21'heabd2;
        #1
        src0 <= 16'h9d6;
        src1 <= 16'h90fb;
        src2 <= 16'h47bb;
        src3 <= 16'h51d7;
        src4 <= 16'h69d1;
        src5 <= 16'h671d;
        src6 <= 16'h6f48;
        src7 <= 16'hcd3c;
        src8 <= 16'heeab;
        src9 <= 16'hd591;
        src10 <= 16'h7605;
        src11 <= 16'hd47c;
        src12 <= 16'hfd4;
        src13 <= 16'h14a1;
        src14 <= 16'hd322;
        src15 <= 16'h195b;
        src16 <= 16'hd884;
        src17 <= 16'h62c2;
        src18 <= 16'h6684;
        src19 <= 16'h6edf;
        src20 <= 16'h76aa;
        src21 <= 16'h1292;
        src22 <= 16'h4c9c;
        src23 <= 16'h7f3f;
        src24 <= 16'hefd0;
        src25 <= 16'h8ac9;
        src26 <= 16'h30fa;
        src27 <= 16'h2191;
        src28 <= 16'h3642;
        src29 <= 16'h57b8;
        src30 <= 16'ha3bb;
        src31 <= 16'hbb3;
        exp <= 21'hdd1d0;
        #1
        src0 <= 16'h7651;
        src1 <= 16'hed45;
        src2 <= 16'h2329;
        src3 <= 16'hb90a;
        src4 <= 16'h7263;
        src5 <= 16'he896;
        src6 <= 16'h79f;
        src7 <= 16'h6fca;
        src8 <= 16'hfce5;
        src9 <= 16'h5906;
        src10 <= 16'h168b;
        src11 <= 16'h1646;
        src12 <= 16'h28af;
        src13 <= 16'he0e5;
        src14 <= 16'ha95d;
        src15 <= 16'hb203;
        src16 <= 16'haac4;
        src17 <= 16'haa8a;
        src18 <= 16'h4815;
        src19 <= 16'h8c93;
        src20 <= 16'h5db;
        src21 <= 16'h9a3f;
        src22 <= 16'h87a9;
        src23 <= 16'h25ab;
        src24 <= 16'h3de0;
        src25 <= 16'h9b48;
        src26 <= 16'hb66d;
        src27 <= 16'h512a;
        src28 <= 16'h3f40;
        src29 <= 16'he142;
        src30 <= 16'hb94e;
        src31 <= 16'h6879;
        exp <= 21'hf9447;
        #1
        src0 <= 16'hfa34;
        src1 <= 16'he6f5;
        src2 <= 16'h6b24;
        src3 <= 16'h5865;
        src4 <= 16'hd5b1;
        src5 <= 16'hf084;
        src6 <= 16'h627a;
        src7 <= 16'hbd39;
        src8 <= 16'h6f93;
        src9 <= 16'haedf;
        src10 <= 16'h1f8b;
        src11 <= 16'h9ea3;
        src12 <= 16'h821b;
        src13 <= 16'h91dc;
        src14 <= 16'h98fe;
        src15 <= 16'hf3d1;
        src16 <= 16'h3397;
        src17 <= 16'hde4e;
        src18 <= 16'h7bcf;
        src19 <= 16'h807e;
        src20 <= 16'h3b7b;
        src21 <= 16'ha580;
        src22 <= 16'h2af9;
        src23 <= 16'h442d;
        src24 <= 16'h6cd;
        src25 <= 16'h336a;
        src26 <= 16'hbe9;
        src27 <= 16'hd09e;
        src28 <= 16'h14a6;
        src29 <= 16'hcf9d;
        src30 <= 16'h7e87;
        src31 <= 16'hc2ac;
        exp <= 21'h10a287;
        #1
        src0 <= 16'h55af;
        src1 <= 16'h378f;
        src2 <= 16'h21ef;
        src3 <= 16'h92b0;
        src4 <= 16'h49c7;
        src5 <= 16'hfd0;
        src6 <= 16'hf05b;
        src7 <= 16'h8ed7;
        src8 <= 16'h363;
        src9 <= 16'h96aa;
        src10 <= 16'h1949;
        src11 <= 16'h3ff3;
        src12 <= 16'h15b6;
        src13 <= 16'hfee0;
        src14 <= 16'he545;
        src15 <= 16'hb21d;
        src16 <= 16'h58aa;
        src17 <= 16'h3c6a;
        src18 <= 16'hcbc6;
        src19 <= 16'h8a41;
        src20 <= 16'h46dc;
        src21 <= 16'h319e;
        src22 <= 16'h6efd;
        src23 <= 16'h66a9;
        src24 <= 16'hd24f;
        src25 <= 16'hdf97;
        src26 <= 16'hb1df;
        src27 <= 16'h4cc8;
        src28 <= 16'ha7e9;
        src29 <= 16'h96d8;
        src30 <= 16'hf657;
        src31 <= 16'h2537;
        exp <= 21'hefdfe;
        #1
        src0 <= 16'hc1e5;
        src1 <= 16'h1e78;
        src2 <= 16'h4c81;
        src3 <= 16'he6bc;
        src4 <= 16'h5d30;
        src5 <= 16'he3d4;
        src6 <= 16'h8708;
        src7 <= 16'hedf4;
        src8 <= 16'hf078;
        src9 <= 16'h753;
        src10 <= 16'h72ad;
        src11 <= 16'h5bf3;
        src12 <= 16'hf473;
        src13 <= 16'haa6a;
        src14 <= 16'hf330;
        src15 <= 16'hef43;
        src16 <= 16'hfe9;
        src17 <= 16'ha655;
        src18 <= 16'he0e8;
        src19 <= 16'hb4cc;
        src20 <= 16'h22a7;
        src21 <= 16'h266b;
        src22 <= 16'h983b;
        src23 <= 16'h8e66;
        src24 <= 16'hded2;
        src25 <= 16'h1850;
        src26 <= 16'h4244;
        src27 <= 16'h4f00;
        src28 <= 16'h8a08;
        src29 <= 16'h89e4;
        src30 <= 16'h36cf;
        src31 <= 16'h6d2b;
        exp <= 21'h110d46;
        #1
        src0 <= 16'h1e6c;
        src1 <= 16'h2c77;
        src2 <= 16'h4a68;
        src3 <= 16'h82bf;
        src4 <= 16'hce97;
        src5 <= 16'h5601;
        src6 <= 16'hf6e6;
        src7 <= 16'hde1c;
        src8 <= 16'hbbbc;
        src9 <= 16'h96b9;
        src10 <= 16'hf5a6;
        src11 <= 16'hbc9e;
        src12 <= 16'h96c4;
        src13 <= 16'hd9f3;
        src14 <= 16'h65f;
        src15 <= 16'h626;
        src16 <= 16'hfd1a;
        src17 <= 16'h5aa7;
        src18 <= 16'hde72;
        src19 <= 16'ha1aa;
        src20 <= 16'hf36;
        src21 <= 16'hcd7f;
        src22 <= 16'h6db4;
        src23 <= 16'h5634;
        src24 <= 16'h7f89;
        src25 <= 16'hf84d;
        src26 <= 16'hec9;
        src27 <= 16'hd2f5;
        src28 <= 16'h30e7;
        src29 <= 16'hf48;
        src30 <= 16'hcc09;
        src31 <= 16'h445d;
        exp <= 21'h10b63c;
        #1
        src0 <= 16'h2c58;
        src1 <= 16'h22b9;
        src2 <= 16'h90d4;
        src3 <= 16'h8f92;
        src4 <= 16'h846d;
        src5 <= 16'h9309;
        src6 <= 16'h960a;
        src7 <= 16'hfcba;
        src8 <= 16'ha8c9;
        src9 <= 16'h997e;
        src10 <= 16'h96a6;
        src11 <= 16'h94b5;
        src12 <= 16'hb043;
        src13 <= 16'h1ed8;
        src14 <= 16'h39bb;
        src15 <= 16'h6044;
        src16 <= 16'heaf6;
        src17 <= 16'h3c60;
        src18 <= 16'h8abc;
        src19 <= 16'hb647;
        src20 <= 16'h10b5;
        src21 <= 16'h1c01;
        src22 <= 16'hb446;
        src23 <= 16'hc36d;
        src24 <= 16'h381a;
        src25 <= 16'h96e7;
        src26 <= 16'hde7d;
        src27 <= 16'hf891;
        src28 <= 16'h224;
        src29 <= 16'he5ee;
        src30 <= 16'h386c;
        src31 <= 16'hd110;
        exp <= 21'h1094cc;
        #1
        src0 <= 16'hf1e7;
        src1 <= 16'h1c21;
        src2 <= 16'h85bf;
        src3 <= 16'h7875;
        src4 <= 16'h3def;
        src5 <= 16'he95;
        src6 <= 16'h4a5e;
        src7 <= 16'h463b;
        src8 <= 16'hd294;
        src9 <= 16'hd8c3;
        src10 <= 16'hac8b;
        src11 <= 16'hf8de;
        src12 <= 16'haca1;
        src13 <= 16'h1f11;
        src14 <= 16'h79c2;
        src15 <= 16'h35aa;
        src16 <= 16'he564;
        src17 <= 16'ha02e;
        src18 <= 16'hede1;
        src19 <= 16'h60bb;
        src20 <= 16'hed08;
        src21 <= 16'hdc6c;
        src22 <= 16'h1cb3;
        src23 <= 16'hdac3;
        src24 <= 16'ha91;
        src25 <= 16'ha353;
        src26 <= 16'he1b5;
        src27 <= 16'ha3ca;
        src28 <= 16'hbcb7;
        src29 <= 16'ha3d0;
        src30 <= 16'hd327;
        src31 <= 16'h5040;
        exp <= 21'h1201a0;
        #1
        src0 <= 16'h6e0f;
        src1 <= 16'hb315;
        src2 <= 16'h2cbe;
        src3 <= 16'h67db;
        src4 <= 16'h1d2c;
        src5 <= 16'ha616;
        src6 <= 16'h39b5;
        src7 <= 16'h6c32;
        src8 <= 16'h34df;
        src9 <= 16'hf519;
        src10 <= 16'hfcae;
        src11 <= 16'hd6fc;
        src12 <= 16'h3645;
        src13 <= 16'h1f27;
        src14 <= 16'hd448;
        src15 <= 16'had62;
        src16 <= 16'ha255;
        src17 <= 16'h69e2;
        src18 <= 16'h7744;
        src19 <= 16'h6779;
        src20 <= 16'hdbaf;
        src21 <= 16'heae5;
        src22 <= 16'h1276;
        src23 <= 16'h4032;
        src24 <= 16'h2d90;
        src25 <= 16'haa3e;
        src26 <= 16'hafa1;
        src27 <= 16'h6fa6;
        src28 <= 16'he392;
        src29 <= 16'h9512;
        src30 <= 16'hff14;
        src31 <= 16'h5c55;
        exp <= 21'h10c2f0;
        #1
        src0 <= 16'he4df;
        src1 <= 16'hcd83;
        src2 <= 16'h4702;
        src3 <= 16'h29f8;
        src4 <= 16'he573;
        src5 <= 16'h6c1f;
        src6 <= 16'h1693;
        src7 <= 16'h125f;
        src8 <= 16'h5cf9;
        src9 <= 16'h4cf3;
        src10 <= 16'h4e7a;
        src11 <= 16'hef9a;
        src12 <= 16'hda45;
        src13 <= 16'hf6e1;
        src14 <= 16'h33e;
        src15 <= 16'h63b3;
        src16 <= 16'h42c3;
        src17 <= 16'h39be;
        src18 <= 16'hb3d9;
        src19 <= 16'h7922;
        src20 <= 16'h3dd9;
        src21 <= 16'hb0d8;
        src22 <= 16'h90f1;
        src23 <= 16'hf6f3;
        src24 <= 16'hbe93;
        src25 <= 16'ha811;
        src26 <= 16'h5558;
        src27 <= 16'hf552;
        src28 <= 16'h9a24;
        src29 <= 16'h110f;
        src30 <= 16'hf2a6;
        src31 <= 16'h43d1;
        exp <= 21'h107100;
        #1
        src0 <= 16'h6f16;
        src1 <= 16'h2e16;
        src2 <= 16'h1a07;
        src3 <= 16'hd204;
        src4 <= 16'h690;
        src5 <= 16'h3;
        src6 <= 16'hf7ee;
        src7 <= 16'h23a8;
        src8 <= 16'h1bf7;
        src9 <= 16'h5bf6;
        src10 <= 16'h4708;
        src11 <= 16'h54a0;
        src12 <= 16'hbb92;
        src13 <= 16'hbde2;
        src14 <= 16'h7642;
        src15 <= 16'hdc12;
        src16 <= 16'hc1d1;
        src17 <= 16'h30d5;
        src18 <= 16'hafb2;
        src19 <= 16'h9622;
        src20 <= 16'hbbd8;
        src21 <= 16'hcfa8;
        src22 <= 16'hf14d;
        src23 <= 16'hb407;
        src24 <= 16'h4179;
        src25 <= 16'hd20d;
        src26 <= 16'h3237;
        src27 <= 16'h53f;
        src28 <= 16'h5d9;
        src29 <= 16'h3abc;
        src30 <= 16'h1395;
        src31 <= 16'h750e;
        exp <= 21'he083f;
        #1
        src0 <= 16'h9c2b;
        src1 <= 16'h6dd7;
        src2 <= 16'h3a4b;
        src3 <= 16'hf283;
        src4 <= 16'h7a10;
        src5 <= 16'h106e;
        src6 <= 16'h9486;
        src7 <= 16'h5c58;
        src8 <= 16'ha7c4;
        src9 <= 16'h3cd3;
        src10 <= 16'h41c3;
        src11 <= 16'h530e;
        src12 <= 16'hafc;
        src13 <= 16'h3d0a;
        src14 <= 16'h8f74;
        src15 <= 16'hc49c;
        src16 <= 16'hc034;
        src17 <= 16'h517;
        src18 <= 16'hde65;
        src19 <= 16'hffb9;
        src20 <= 16'h1b9e;
        src21 <= 16'h8c55;
        src22 <= 16'hec60;
        src23 <= 16'hcd0;
        src24 <= 16'h6fa;
        src25 <= 16'h108b;
        src26 <= 16'hbb91;
        src27 <= 16'h27a2;
        src28 <= 16'h8381;
        src29 <= 16'ha739;
        src30 <= 16'h5707;
        src31 <= 16'h4b9c;
        exp <= 21'hdd44b;
        #1
        src0 <= 16'he673;
        src1 <= 16'hcfe;
        src2 <= 16'h85d5;
        src3 <= 16'h120;
        src4 <= 16'h715d;
        src5 <= 16'h757e;
        src6 <= 16'he5d0;
        src7 <= 16'hda8d;
        src8 <= 16'hc1f0;
        src9 <= 16'hc8c6;
        src10 <= 16'hd374;
        src11 <= 16'h58ee;
        src12 <= 16'h7636;
        src13 <= 16'h1251;
        src14 <= 16'h4bb;
        src15 <= 16'h4710;
        src16 <= 16'h19b5;
        src17 <= 16'ha853;
        src18 <= 16'h1d82;
        src19 <= 16'h7589;
        src20 <= 16'hc3be;
        src21 <= 16'hfae9;
        src22 <= 16'hf68c;
        src23 <= 16'hed69;
        src24 <= 16'h61ea;
        src25 <= 16'heebc;
        src26 <= 16'h919;
        src27 <= 16'h5e76;
        src28 <= 16'h3fe0;
        src29 <= 16'hc0a8;
        src30 <= 16'hbd68;
        src31 <= 16'ha300;
        exp <= 21'h10bddc;
        #1
        src0 <= 16'h4e96;
        src1 <= 16'h5602;
        src2 <= 16'h271c;
        src3 <= 16'h2dc2;
        src4 <= 16'h738a;
        src5 <= 16'hd638;
        src6 <= 16'hae3d;
        src7 <= 16'h4b51;
        src8 <= 16'h729e;
        src9 <= 16'h402a;
        src10 <= 16'hdff0;
        src11 <= 16'hb576;
        src12 <= 16'ha606;
        src13 <= 16'h2ed7;
        src14 <= 16'h6ae0;
        src15 <= 16'h340e;
        src16 <= 16'hf083;
        src17 <= 16'h61cf;
        src18 <= 16'h6b80;
        src19 <= 16'hed62;
        src20 <= 16'h97e1;
        src21 <= 16'hc81e;
        src22 <= 16'he910;
        src23 <= 16'h5fc2;
        src24 <= 16'h9b;
        src25 <= 16'h189d;
        src26 <= 16'h7833;
        src27 <= 16'h2710;
        src28 <= 16'h1b6e;
        src29 <= 16'h3f96;
        src30 <= 16'he70e;
        src31 <= 16'h1186;
        exp <= 21'he58d7;
        #1
        src0 <= 16'h4faf;
        src1 <= 16'hd1f5;
        src2 <= 16'hf580;
        src3 <= 16'ha6a8;
        src4 <= 16'h2897;
        src5 <= 16'h9719;
        src6 <= 16'h298f;
        src7 <= 16'h59d7;
        src8 <= 16'h1783;
        src9 <= 16'hc0fb;
        src10 <= 16'h7134;
        src11 <= 16'haeff;
        src12 <= 16'h47f8;
        src13 <= 16'he2c9;
        src14 <= 16'hafd1;
        src15 <= 16'h894a;
        src16 <= 16'ha716;
        src17 <= 16'h5264;
        src18 <= 16'h67c9;
        src19 <= 16'h6048;
        src20 <= 16'h8795;
        src21 <= 16'h7b2a;
        src22 <= 16'hf68c;
        src23 <= 16'hb9b8;
        src24 <= 16'h14fa;
        src25 <= 16'h271d;
        src26 <= 16'hd839;
        src27 <= 16'h2178;
        src28 <= 16'h3de;
        src29 <= 16'ha4e4;
        src30 <= 16'hab7;
        src31 <= 16'hb052;
        exp <= 21'hf6b90;
        #1
        src0 <= 16'h1fa1;
        src1 <= 16'h710b;
        src2 <= 16'hd51d;
        src3 <= 16'h4a07;
        src4 <= 16'h1be9;
        src5 <= 16'h8660;
        src6 <= 16'h238c;
        src7 <= 16'h9c5d;
        src8 <= 16'h6a80;
        src9 <= 16'h1728;
        src10 <= 16'h9f03;
        src11 <= 16'hfee2;
        src12 <= 16'h8b52;
        src13 <= 16'hff7a;
        src14 <= 16'hf724;
        src15 <= 16'h5a91;
        src16 <= 16'h11cd;
        src17 <= 16'h8448;
        src18 <= 16'hcd;
        src19 <= 16'h897b;
        src20 <= 16'hfc0;
        src21 <= 16'he3c8;
        src22 <= 16'h3921;
        src23 <= 16'hd459;
        src24 <= 16'hca6f;
        src25 <= 16'h26d;
        src26 <= 16'h7890;
        src27 <= 16'ha66f;
        src28 <= 16'he103;
        src29 <= 16'h12d4;
        src30 <= 16'h8213;
        src31 <= 16'h823b;
        exp <= 21'hf136f;
        #1
        src0 <= 16'hf28b;
        src1 <= 16'h40a;
        src2 <= 16'hc8e4;
        src3 <= 16'h28d6;
        src4 <= 16'h5105;
        src5 <= 16'hde91;
        src6 <= 16'h8f09;
        src7 <= 16'h25c1;
        src8 <= 16'hf1bb;
        src9 <= 16'h74c5;
        src10 <= 16'h5eb4;
        src11 <= 16'h122b;
        src12 <= 16'hc8b1;
        src13 <= 16'ha83d;
        src14 <= 16'h784;
        src15 <= 16'h8760;
        src16 <= 16'h7a60;
        src17 <= 16'ha729;
        src18 <= 16'h34a1;
        src19 <= 16'hbf41;
        src20 <= 16'hfd0e;
        src21 <= 16'h8763;
        src22 <= 16'h178b;
        src23 <= 16'h23ac;
        src24 <= 16'h519e;
        src25 <= 16'h83f2;
        src26 <= 16'ha7a;
        src27 <= 16'hc06a;
        src28 <= 16'h2be7;
        src29 <= 16'h59da;
        src30 <= 16'h6079;
        src31 <= 16'h3ed7;
        exp <= 21'he3e78;
        #1
        src0 <= 16'he61;
        src1 <= 16'h4f13;
        src2 <= 16'h59c0;
        src3 <= 16'h872f;
        src4 <= 16'h650;
        src5 <= 16'h1aa;
        src6 <= 16'h7570;
        src7 <= 16'h9435;
        src8 <= 16'h56fb;
        src9 <= 16'hbd9;
        src10 <= 16'hd0c4;
        src11 <= 16'h22f4;
        src12 <= 16'h4d96;
        src13 <= 16'h78b6;
        src14 <= 16'h8454;
        src15 <= 16'hd4a8;
        src16 <= 16'hfd9;
        src17 <= 16'h5737;
        src18 <= 16'h7b81;
        src19 <= 16'h1067;
        src20 <= 16'h6734;
        src21 <= 16'h5134;
        src22 <= 16'h65f1;
        src23 <= 16'h90e5;
        src24 <= 16'h149f;
        src25 <= 16'h492d;
        src26 <= 16'hbc15;
        src27 <= 16'h644;
        src28 <= 16'h3720;
        src29 <= 16'hc562;
        src30 <= 16'h922c;
        src31 <= 16'hc2e8;
        exp <= 21'hbd9c7;
        #1
        src0 <= 16'hd42e;
        src1 <= 16'h854d;
        src2 <= 16'hb7ac;
        src3 <= 16'h2fff;
        src4 <= 16'hcb52;
        src5 <= 16'h5b82;
        src6 <= 16'haa47;
        src7 <= 16'hc517;
        src8 <= 16'h3c8b;
        src9 <= 16'hc0fd;
        src10 <= 16'hae53;
        src11 <= 16'he1fa;
        src12 <= 16'hfb74;
        src13 <= 16'hd178;
        src14 <= 16'ha278;
        src15 <= 16'h6d6f;
        src16 <= 16'h4b97;
        src17 <= 16'h94d0;
        src18 <= 16'h56d2;
        src19 <= 16'h5d8b;
        src20 <= 16'h390a;
        src21 <= 16'hfe9b;
        src22 <= 16'h5970;
        src23 <= 16'ha5a5;
        src24 <= 16'h4ad5;
        src25 <= 16'hdcf6;
        src26 <= 16'h7b00;
        src27 <= 16'h114;
        src28 <= 16'hc48c;
        src29 <= 16'h7414;
        src30 <= 16'h5e40;
        src31 <= 16'he6a6;
        exp <= 21'h122ee3;
        #1
        src0 <= 16'h4c9;
        src1 <= 16'h4b91;
        src2 <= 16'he1f1;
        src3 <= 16'h422d;
        src4 <= 16'hda92;
        src5 <= 16'hbf67;
        src6 <= 16'hd673;
        src7 <= 16'hdf10;
        src8 <= 16'h17e4;
        src9 <= 16'hebd8;
        src10 <= 16'h822e;
        src11 <= 16'hbf7e;
        src12 <= 16'he66b;
        src13 <= 16'h8148;
        src14 <= 16'hbdd8;
        src15 <= 16'h9971;
        src16 <= 16'hbe6e;
        src17 <= 16'h53e3;
        src18 <= 16'h81bc;
        src19 <= 16'hdc3b;
        src20 <= 16'h5f3f;
        src21 <= 16'h7ed2;
        src22 <= 16'ha6ab;
        src23 <= 16'hcb9a;
        src24 <= 16'h49a8;
        src25 <= 16'he16f;
        src26 <= 16'h993a;
        src27 <= 16'he6d9;
        src28 <= 16'hf103;
        src29 <= 16'hbc31;
        src30 <= 16'h57a6;
        src31 <= 16'h2fa8;
        exp <= 21'h1368a2;
        #1
        src0 <= 16'hc204;
        src1 <= 16'hd414;
        src2 <= 16'h7154;
        src3 <= 16'he649;
        src4 <= 16'h6783;
        src5 <= 16'h9261;
        src6 <= 16'h3516;
        src7 <= 16'h35c4;
        src8 <= 16'hd6bd;
        src9 <= 16'hb3a3;
        src10 <= 16'he1ca;
        src11 <= 16'h5e72;
        src12 <= 16'h74d3;
        src13 <= 16'h815;
        src14 <= 16'hd5c5;
        src15 <= 16'h9735;
        src16 <= 16'hcf22;
        src17 <= 16'hbb35;
        src18 <= 16'h4294;
        src19 <= 16'h4622;
        src20 <= 16'h4e53;
        src21 <= 16'h8406;
        src22 <= 16'h9473;
        src23 <= 16'h78e9;
        src24 <= 16'h34e9;
        src25 <= 16'h33f1;
        src26 <= 16'h837d;
        src27 <= 16'h7715;
        src28 <= 16'h6003;
        src29 <= 16'h8e13;
        src30 <= 16'he521;
        src31 <= 16'h22b1;
        exp <= 21'h105307;
        #1
        src0 <= 16'hc249;
        src1 <= 16'h2fc7;
        src2 <= 16'h63b;
        src3 <= 16'hdee3;
        src4 <= 16'hbac6;
        src5 <= 16'hf6a4;
        src6 <= 16'he185;
        src7 <= 16'h500a;
        src8 <= 16'h8cb8;
        src9 <= 16'hcc8e;
        src10 <= 16'h233c;
        src11 <= 16'hf76b;
        src12 <= 16'h1901;
        src13 <= 16'h7834;
        src14 <= 16'hf9bb;
        src15 <= 16'h6d10;
        src16 <= 16'h2d3b;
        src17 <= 16'h3341;
        src18 <= 16'hd055;
        src19 <= 16'h1396;
        src20 <= 16'had4a;
        src21 <= 16'hd0aa;
        src22 <= 16'h48d6;
        src23 <= 16'hf2aa;
        src24 <= 16'hdd5;
        src25 <= 16'h275e;
        src26 <= 16'h322a;
        src27 <= 16'hb4fa;
        src28 <= 16'h1e9a;
        src29 <= 16'h8b40;
        src30 <= 16'h1c0b;
        src31 <= 16'he443;
        exp <= 21'hfea6e;
        #1
        src0 <= 16'h2e45;
        src1 <= 16'hbb9a;
        src2 <= 16'hf392;
        src3 <= 16'h359;
        src4 <= 16'h2343;
        src5 <= 16'hba49;
        src6 <= 16'h2f62;
        src7 <= 16'hf58f;
        src8 <= 16'hc3c;
        src9 <= 16'h249d;
        src10 <= 16'h4b4a;
        src11 <= 16'hc4b3;
        src12 <= 16'hbb63;
        src13 <= 16'h2f95;
        src14 <= 16'h4141;
        src15 <= 16'hf8e0;
        src16 <= 16'h23a5;
        src17 <= 16'h75dc;
        src18 <= 16'ha0c5;
        src19 <= 16'h630f;
        src20 <= 16'h1bbf;
        src21 <= 16'h9a06;
        src22 <= 16'hd0ce;
        src23 <= 16'hd1e;
        src24 <= 16'hf670;
        src25 <= 16'h537b;
        src26 <= 16'hc101;
        src27 <= 16'h9b42;
        src28 <= 16'hf956;
        src29 <= 16'he454;
        src30 <= 16'h5539;
        src31 <= 16'h91a2;
        exp <= 21'hfe4ef;
        #1
        src0 <= 16'hfbd3;
        src1 <= 16'h845e;
        src2 <= 16'h34cd;
        src3 <= 16'h8506;
        src4 <= 16'h7330;
        src5 <= 16'he6ce;
        src6 <= 16'h1c0a;
        src7 <= 16'hff67;
        src8 <= 16'h2ad8;
        src9 <= 16'heb4f;
        src10 <= 16'h7ce1;
        src11 <= 16'hb672;
        src12 <= 16'h8385;
        src13 <= 16'h2235;
        src14 <= 16'hccc7;
        src15 <= 16'h2ce0;
        src16 <= 16'h70a2;
        src17 <= 16'h83db;
        src18 <= 16'h412b;
        src19 <= 16'h474b;
        src20 <= 16'h73df;
        src21 <= 16'hc588;
        src22 <= 16'hd724;
        src23 <= 16'h44d2;
        src24 <= 16'h57fc;
        src25 <= 16'hae05;
        src26 <= 16'h2bcd;
        src27 <= 16'hb039;
        src28 <= 16'hf23a;
        src29 <= 16'hd988;
        src30 <= 16'ha6b;
        src31 <= 16'hed1c;
        exp <= 21'h110fee;
        #1
        src0 <= 16'h866c;
        src1 <= 16'hc80c;
        src2 <= 16'h11d8;
        src3 <= 16'h6a50;
        src4 <= 16'h75b6;
        src5 <= 16'hdefd;
        src6 <= 16'ha34f;
        src7 <= 16'hfbc2;
        src8 <= 16'h9662;
        src9 <= 16'h3b12;
        src10 <= 16'h137;
        src11 <= 16'h25b8;
        src12 <= 16'h4585;
        src13 <= 16'hb509;
        src14 <= 16'h9d42;
        src15 <= 16'h3d20;
        src16 <= 16'h847d;
        src17 <= 16'h9a3b;
        src18 <= 16'hb1d8;
        src19 <= 16'hdd80;
        src20 <= 16'hd94c;
        src21 <= 16'hacf8;
        src22 <= 16'hbc50;
        src23 <= 16'h2676;
        src24 <= 16'h6dc6;
        src25 <= 16'h9c53;
        src26 <= 16'h2cc7;
        src27 <= 16'h9755;
        src28 <= 16'h9963;
        src29 <= 16'hc7b2;
        src30 <= 16'hee62;
        src31 <= 16'hd7e6;
        exp <= 21'h119863;
        #1
        $finish;
    end
endmodule

