module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    compressor_CLA64_64 compressor_CLA64_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
        src16 <= 64'h0;
        src17 <= 64'h0;
        src18 <= 64'h0;
        src19 <= 64'h0;
        src20 <= 64'h0;
        src21 <= 64'h0;
        src22 <= 64'h0;
        src23 <= 64'h0;
        src24 <= 64'h0;
        src25 <= 64'h0;
        src26 <= 64'h0;
        src27 <= 64'h0;
        src28 <= 64'h0;
        src29 <= 64'h0;
        src30 <= 64'h0;
        src31 <= 64'h0;
        src32 <= 64'h0;
        src33 <= 64'h0;
        src34 <= 64'h0;
        src35 <= 64'h0;
        src36 <= 64'h0;
        src37 <= 64'h0;
        src38 <= 64'h0;
        src39 <= 64'h0;
        src40 <= 64'h0;
        src41 <= 64'h0;
        src42 <= 64'h0;
        src43 <= 64'h0;
        src44 <= 64'h0;
        src45 <= 64'h0;
        src46 <= 64'h0;
        src47 <= 64'h0;
        src48 <= 64'h0;
        src49 <= 64'h0;
        src50 <= 64'h0;
        src51 <= 64'h0;
        src52 <= 64'h0;
        src53 <= 64'h0;
        src54 <= 64'h0;
        src55 <= 64'h0;
        src56 <= 64'h0;
        src57 <= 64'h0;
        src58 <= 64'h0;
        src59 <= 64'h0;
        src60 <= 64'h0;
        src61 <= 64'h0;
        src62 <= 64'h0;
        src63 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA64_64(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    input [63:0]src16,
    input [63:0]src17,
    input [63:0]src18,
    input [63:0]src19,
    input [63:0]src20,
    input [63:0]src21,
    input [63:0]src22,
    input [63:0]src23,
    input [63:0]src24,
    input [63:0]src25,
    input [63:0]src26,
    input [63:0]src27,
    input [63:0]src28,
    input [63:0]src29,
    input [63:0]src30,
    input [63:0]src31,
    input [63:0]src32,
    input [63:0]src33,
    input [63:0]src34,
    input [63:0]src35,
    input [63:0]src36,
    input [63:0]src37,
    input [63:0]src38,
    input [63:0]src39,
    input [63:0]src40,
    input [63:0]src41,
    input [63:0]src42,
    input [63:0]src43,
    input [63:0]src44,
    input [63:0]src45,
    input [63:0]src46,
    input [63:0]src47,
    input [63:0]src48,
    input [63:0]src49,
    input [63:0]src50,
    input [63:0]src51,
    input [63:0]src52,
    input [63:0]src53,
    input [63:0]src54,
    input [63:0]src55,
    input [63:0]src56,
    input [63:0]src57,
    input [63:0]src58,
    input [63:0]src59,
    input [63:0]src60,
    input [63:0]src61,
    input [63:0]src62,
    input [63:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [0:0] comp_out67;
    wire [1:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out68[1], 1'h0, comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      input wire [63:0] src32,
      input wire [63:0] src33,
      input wire [63:0] src34,
      input wire [63:0] src35,
      input wire [63:0] src36,
      input wire [63:0] src37,
      input wire [63:0] src38,
      input wire [63:0] src39,
      input wire [63:0] src40,
      input wire [63:0] src41,
      input wire [63:0] src42,
      input wire [63:0] src43,
      input wire [63:0] src44,
      input wire [63:0] src45,
      input wire [63:0] src46,
      input wire [63:0] src47,
      input wire [63:0] src48,
      input wire [63:0] src49,
      input wire [63:0] src50,
      input wire [63:0] src51,
      input wire [63:0] src52,
      input wire [63:0] src53,
      input wire [63:0] src54,
      input wire [63:0] src55,
      input wire [63:0] src56,
      input wire [63:0] src57,
      input wire [63:0] src58,
      input wire [63:0] src59,
      input wire [63:0] src60,
      input wire [63:0] src61,
      input wire [63:0] src62,
      input wire [63:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [0:0] dst67,
      output wire [1:0] dst68,
      output wire [0:0] dst69);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [63:0] stage0_16;
   wire [63:0] stage0_17;
   wire [63:0] stage0_18;
   wire [63:0] stage0_19;
   wire [63:0] stage0_20;
   wire [63:0] stage0_21;
   wire [63:0] stage0_22;
   wire [63:0] stage0_23;
   wire [63:0] stage0_24;
   wire [63:0] stage0_25;
   wire [63:0] stage0_26;
   wire [63:0] stage0_27;
   wire [63:0] stage0_28;
   wire [63:0] stage0_29;
   wire [63:0] stage0_30;
   wire [63:0] stage0_31;
   wire [63:0] stage0_32;
   wire [63:0] stage0_33;
   wire [63:0] stage0_34;
   wire [63:0] stage0_35;
   wire [63:0] stage0_36;
   wire [63:0] stage0_37;
   wire [63:0] stage0_38;
   wire [63:0] stage0_39;
   wire [63:0] stage0_40;
   wire [63:0] stage0_41;
   wire [63:0] stage0_42;
   wire [63:0] stage0_43;
   wire [63:0] stage0_44;
   wire [63:0] stage0_45;
   wire [63:0] stage0_46;
   wire [63:0] stage0_47;
   wire [63:0] stage0_48;
   wire [63:0] stage0_49;
   wire [63:0] stage0_50;
   wire [63:0] stage0_51;
   wire [63:0] stage0_52;
   wire [63:0] stage0_53;
   wire [63:0] stage0_54;
   wire [63:0] stage0_55;
   wire [63:0] stage0_56;
   wire [63:0] stage0_57;
   wire [63:0] stage0_58;
   wire [63:0] stage0_59;
   wire [63:0] stage0_60;
   wire [63:0] stage0_61;
   wire [63:0] stage0_62;
   wire [63:0] stage0_63;
   wire [18:0] stage1_0;
   wire [47:0] stage1_1;
   wire [23:0] stage1_2;
   wire [27:0] stage1_3;
   wire [37:0] stage1_4;
   wire [26:0] stage1_5;
   wire [21:0] stage1_6;
   wire [35:0] stage1_7;
   wire [26:0] stage1_8;
   wire [28:0] stage1_9;
   wire [33:0] stage1_10;
   wire [32:0] stage1_11;
   wire [26:0] stage1_12;
   wire [30:0] stage1_13;
   wire [24:0] stage1_14;
   wire [44:0] stage1_15;
   wire [30:0] stage1_16;
   wire [44:0] stage1_17;
   wire [22:0] stage1_18;
   wire [28:0] stage1_19;
   wire [40:0] stage1_20;
   wire [32:0] stage1_21;
   wire [30:0] stage1_22;
   wire [34:0] stage1_23;
   wire [26:0] stage1_24;
   wire [44:0] stage1_25;
   wire [28:0] stage1_26;
   wire [40:0] stage1_27;
   wire [26:0] stage1_28;
   wire [28:0] stage1_29;
   wire [25:0] stage1_30;
   wire [22:0] stage1_31;
   wire [30:0] stage1_32;
   wire [37:0] stage1_33;
   wire [23:0] stage1_34;
   wire [29:0] stage1_35;
   wire [43:0] stage1_36;
   wire [23:0] stage1_37;
   wire [41:0] stage1_38;
   wire [22:0] stage1_39;
   wire [26:0] stage1_40;
   wire [35:0] stage1_41;
   wire [28:0] stage1_42;
   wire [35:0] stage1_43;
   wire [32:0] stage1_44;
   wire [47:0] stage1_45;
   wire [16:0] stage1_46;
   wire [40:0] stage1_47;
   wire [31:0] stage1_48;
   wire [24:0] stage1_49;
   wire [24:0] stage1_50;
   wire [31:0] stage1_51;
   wire [42:0] stage1_52;
   wire [26:0] stage1_53;
   wire [32:0] stage1_54;
   wire [24:0] stage1_55;
   wire [25:0] stage1_56;
   wire [25:0] stage1_57;
   wire [40:0] stage1_58;
   wire [41:0] stage1_59;
   wire [32:0] stage1_60;
   wire [30:0] stage1_61;
   wire [32:0] stage1_62;
   wire [27:0] stage1_63;
   wire [15:0] stage1_64;
   wire [8:0] stage1_65;
   wire [5:0] stage2_0;
   wire [8:0] stage2_1;
   wire [11:0] stage2_2;
   wire [11:0] stage2_3;
   wire [25:0] stage2_4;
   wire [21:0] stage2_5;
   wire [13:0] stage2_6;
   wire [19:0] stage2_7;
   wire [19:0] stage2_8;
   wire [10:0] stage2_9;
   wire [30:0] stage2_10;
   wire [15:0] stage2_11;
   wire [18:0] stage2_12;
   wire [8:0] stage2_13;
   wire [15:0] stage2_14;
   wire [20:0] stage2_15;
   wire [15:0] stage2_16;
   wire [21:0] stage2_17;
   wire [18:0] stage2_18;
   wire [14:0] stage2_19;
   wire [23:0] stage2_20;
   wire [12:0] stage2_21;
   wire [10:0] stage2_22;
   wire [16:0] stage2_23;
   wire [13:0] stage2_24;
   wire [13:0] stage2_25;
   wire [19:0] stage2_26;
   wire [25:0] stage2_27;
   wire [15:0] stage2_28;
   wire [9:0] stage2_29;
   wire [19:0] stage2_30;
   wire [12:0] stage2_31;
   wire [18:0] stage2_32;
   wire [22:0] stage2_33;
   wire [12:0] stage2_34;
   wire [12:0] stage2_35;
   wire [17:0] stage2_36;
   wire [17:0] stage2_37;
   wire [23:0] stage2_38;
   wire [12:0] stage2_39;
   wire [11:0] stage2_40;
   wire [19:0] stage2_41;
   wire [14:0] stage2_42;
   wire [12:0] stage2_43;
   wire [17:0] stage2_44;
   wire [13:0] stage2_45;
   wire [11:0] stage2_46;
   wire [18:0] stage2_47;
   wire [16:0] stage2_48;
   wire [10:0] stage2_49;
   wire [11:0] stage2_50;
   wire [15:0] stage2_51;
   wire [11:0] stage2_52;
   wire [17:0] stage2_53;
   wire [14:0] stage2_54;
   wire [16:0] stage2_55;
   wire [9:0] stage2_56;
   wire [13:0] stage2_57;
   wire [17:0] stage2_58;
   wire [19:0] stage2_59;
   wire [13:0] stage2_60;
   wire [14:0] stage2_61;
   wire [12:0] stage2_62;
   wire [12:0] stage2_63;
   wire [10:0] stage2_64;
   wire [7:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage2_67;
   wire [5:0] stage3_0;
   wire [3:0] stage3_1;
   wire [2:0] stage3_2;
   wire [4:0] stage3_3;
   wire [6:0] stage3_4;
   wire [8:0] stage3_5;
   wire [7:0] stage3_6;
   wire [10:0] stage3_7;
   wire [8:0] stage3_8;
   wire [11:0] stage3_9;
   wire [6:0] stage3_10;
   wire [8:0] stage3_11;
   wire [7:0] stage3_12;
   wire [8:0] stage3_13;
   wire [6:0] stage3_14;
   wire [8:0] stage3_15;
   wire [7:0] stage3_16;
   wire [6:0] stage3_17;
   wire [12:0] stage3_18;
   wire [6:0] stage3_19;
   wire [5:0] stage3_20;
   wire [8:0] stage3_21;
   wire [6:0] stage3_22;
   wire [7:0] stage3_23;
   wire [6:0] stage3_24;
   wire [7:0] stage3_25;
   wire [6:0] stage3_26;
   wire [6:0] stage3_27;
   wire [8:0] stage3_28;
   wire [8:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [6:0] stage3_32;
   wire [16:0] stage3_33;
   wire [6:0] stage3_34;
   wire [5:0] stage3_35;
   wire [9:0] stage3_36;
   wire [5:0] stage3_37;
   wire [10:0] stage3_38;
   wire [6:0] stage3_39;
   wire [5:0] stage3_40;
   wire [13:0] stage3_41;
   wire [3:0] stage3_42;
   wire [5:0] stage3_43;
   wire [16:0] stage3_44;
   wire [4:0] stage3_45;
   wire [6:0] stage3_46;
   wire [8:0] stage3_47;
   wire [5:0] stage3_48;
   wire [5:0] stage3_49;
   wire [6:0] stage3_50;
   wire [8:0] stage3_51;
   wire [6:0] stage3_52;
   wire [5:0] stage3_53;
   wire [5:0] stage3_54;
   wire [9:0] stage3_55;
   wire [5:0] stage3_56;
   wire [7:0] stage3_57;
   wire [7:0] stage3_58;
   wire [7:0] stage3_59;
   wire [13:0] stage3_60;
   wire [6:0] stage3_61;
   wire [4:0] stage3_62;
   wire [5:0] stage3_63;
   wire [4:0] stage3_64;
   wire [5:0] stage3_65;
   wire [2:0] stage3_66;
   wire [2:0] stage3_67;
   wire [0:0] stage3_68;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [2:0] stage4_2;
   wire [1:0] stage4_3;
   wire [3:0] stage4_4;
   wire [1:0] stage4_5;
   wire [2:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [4:0] stage4_11;
   wire [2:0] stage4_12;
   wire [3:0] stage4_13;
   wire [3:0] stage4_14;
   wire [3:0] stage4_15;
   wire [4:0] stage4_16;
   wire [2:0] stage4_17;
   wire [3:0] stage4_18;
   wire [2:0] stage4_19;
   wire [3:0] stage4_20;
   wire [7:0] stage4_21;
   wire [1:0] stage4_22;
   wire [3:0] stage4_23;
   wire [3:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [3:0] stage4_27;
   wire [3:0] stage4_28;
   wire [3:0] stage4_29;
   wire [2:0] stage4_30;
   wire [2:0] stage4_31;
   wire [3:0] stage4_32;
   wire [5:0] stage4_33;
   wire [4:0] stage4_34;
   wire [2:0] stage4_35;
   wire [3:0] stage4_36;
   wire [4:0] stage4_37;
   wire [2:0] stage4_38;
   wire [2:0] stage4_39;
   wire [2:0] stage4_40;
   wire [3:0] stage4_41;
   wire [3:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [2:0] stage4_45;
   wire [3:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [3:0] stage4_49;
   wire [3:0] stage4_50;
   wire [5:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [2:0] stage4_54;
   wire [6:0] stage4_55;
   wire [1:0] stage4_56;
   wire [3:0] stage4_57;
   wire [5:0] stage4_58;
   wire [2:0] stage4_59;
   wire [5:0] stage4_60;
   wire [4:0] stage4_61;
   wire [2:0] stage4_62;
   wire [1:0] stage4_63;
   wire [6:0] stage4_64;
   wire [2:0] stage4_65;
   wire [1:0] stage4_66;
   wire [0:0] stage4_67;
   wire [0:0] stage4_68;
   wire [0:0] stage4_69;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [0:0] stage5_67;
   wire [1:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc615_5 gpc14 (
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[5],stage1_4[14],stage1_3[14]}
   );
   gpc615_5 gpc15 (
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[6],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[7],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[8],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc18 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[5],stage1_5[10],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[6],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[7],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[8],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[9],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[10],stage1_5[15],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[11],stage1_5[16],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[12],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[13],stage1_6[13],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[14],stage1_6[14],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[15],stage1_6[15],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[16],stage1_6[16],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[17],stage1_6[17],stage1_5[22]}
   );
   gpc615_5 gpc32 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[30]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[5],stage1_8[13],stage1_7[18],stage1_6[18]}
   );
   gpc615_5 gpc33 (
      {stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_7[31]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[6],stage1_8[14],stage1_7[19],stage1_6[19]}
   );
   gpc615_5 gpc34 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62]},
      {stage0_7[32]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[7],stage1_8[15],stage1_7[20],stage1_6[20]}
   );
   gpc615_5 gpc35 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[8],stage1_8[16],stage1_7[21]}
   );
   gpc615_5 gpc36 (
      {stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42]},
      {stage0_8[19]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[9],stage1_8[17],stage1_7[22]}
   );
   gpc615_5 gpc37 (
      {stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage0_8[20]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[10],stage1_8[18],stage1_7[23]}
   );
   gpc615_5 gpc38 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52]},
      {stage0_8[21]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[11],stage1_8[19],stage1_7[24]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[4],stage1_10[7],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[5],stage1_10[8],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[6],stage1_10[9],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc42 (
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[7],stage1_10[10],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc43 (
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[8],stage1_10[11],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc44 (
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[9],stage1_10[12],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc45 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[10],stage1_10[13],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc46 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[11],stage1_10[14],stage1_9[19]}
   );
   gpc606_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[12],stage1_10[15],stage1_9[20]}
   );
   gpc606_5 gpc48 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[13],stage1_10[16],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[14],stage1_10[17],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[15],stage1_10[18],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[16],stage1_10[19],stage1_9[24]}
   );
   gpc615_5 gpc52 (
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46]},
      {stage0_11[36]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[6],stage1_12[13],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc53 (
      {stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51]},
      {stage0_11[37]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[7],stage1_12[14],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc54 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[8],stage1_12[15],stage1_11[19]}
   );
   gpc615_5 gpc55 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[9],stage1_12[16],stage1_11[20]}
   );
   gpc615_5 gpc56 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52]},
      {stage0_12[14]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[4],stage1_13[10],stage1_12[17],stage1_11[21]}
   );
   gpc606_5 gpc57 (
      {stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[3],stage1_14[5],stage1_13[11],stage1_12[18]}
   );
   gpc606_5 gpc58 (
      {stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[4],stage1_14[6],stage1_13[12],stage1_12[19]}
   );
   gpc606_5 gpc59 (
      {stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[5],stage1_14[7],stage1_13[13],stage1_12[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[6],stage1_14[8],stage1_13[14],stage1_12[21]}
   );
   gpc606_5 gpc61 (
      {stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[7],stage1_14[9],stage1_13[15],stage1_12[22]}
   );
   gpc606_5 gpc62 (
      {stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[8],stage1_14[10],stage1_13[16],stage1_12[23]}
   );
   gpc606_5 gpc63 (
      {stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[9],stage1_14[11],stage1_13[17],stage1_12[24]}
   );
   gpc606_5 gpc64 (
      {stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[10],stage1_14[12],stage1_13[18],stage1_12[25]}
   );
   gpc2135_5 gpc65 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22]},
      {stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[0]},
      {stage0_16[0], stage0_16[1]},
      {stage1_17[0],stage1_16[8],stage1_15[11],stage1_14[13],stage1_13[19]}
   );
   gpc606_5 gpc66 (
      {stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[1],stage1_16[9],stage1_15[12],stage1_14[14],stage1_13[20]}
   );
   gpc606_5 gpc67 (
      {stage0_13[29], stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[2],stage1_16[10],stage1_15[13],stage1_14[15],stage1_13[21]}
   );
   gpc606_5 gpc68 (
      {stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[3],stage1_16[11],stage1_15[14],stage1_14[16],stage1_13[22]}
   );
   gpc606_5 gpc69 (
      {stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage1_17[4],stage1_16[12],stage1_15[15],stage1_14[17],stage1_13[23]}
   );
   gpc606_5 gpc70 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52]},
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30]},
      {stage1_17[5],stage1_16[13],stage1_15[16],stage1_14[18],stage1_13[24]}
   );
   gpc606_5 gpc71 (
      {stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58]},
      {stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36]},
      {stage1_17[6],stage1_16[14],stage1_15[17],stage1_14[19],stage1_13[25]}
   );
   gpc615_5 gpc72 (
      {stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage0_15[37]},
      {stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7]},
      {stage1_18[0],stage1_17[7],stage1_16[15],stage1_15[18],stage1_14[20]}
   );
   gpc615_5 gpc73 (
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage0_15[38]},
      {stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13]},
      {stage1_18[1],stage1_17[8],stage1_16[16],stage1_15[19],stage1_14[21]}
   );
   gpc606_5 gpc74 (
      {stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[9],stage1_16[17]}
   );
   gpc606_5 gpc75 (
      {stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[10],stage1_16[18]}
   );
   gpc606_5 gpc76 (
      {stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[2],stage1_18[4],stage1_17[11],stage1_16[19]}
   );
   gpc606_5 gpc77 (
      {stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[3],stage1_18[5],stage1_17[12],stage1_16[20]}
   );
   gpc615_5 gpc78 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_17[0]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[4],stage1_18[6],stage1_17[13],stage1_16[21]}
   );
   gpc615_5 gpc79 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage0_17[1]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[5],stage1_18[7],stage1_17[14],stage1_16[22]}
   );
   gpc615_5 gpc80 (
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52]},
      {stage0_17[2]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[6],stage1_18[8],stage1_17[15],stage1_16[23]}
   );
   gpc615_5 gpc81 (
      {stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage0_17[3]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[7],stage1_18[9],stage1_17[16],stage1_16[24]}
   );
   gpc606_5 gpc82 (
      {stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[8],stage1_19[8],stage1_18[10],stage1_17[17]}
   );
   gpc606_5 gpc83 (
      {stage0_17[10], stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[9],stage1_19[9],stage1_18[11],stage1_17[18]}
   );
   gpc606_5 gpc84 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[10],stage1_19[10],stage1_18[12],stage1_17[19]}
   );
   gpc606_5 gpc85 (
      {stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[11],stage1_19[11],stage1_18[13],stage1_17[20]}
   );
   gpc606_5 gpc86 (
      {stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[12],stage1_19[12],stage1_18[14],stage1_17[21]}
   );
   gpc606_5 gpc87 (
      {stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[13],stage1_19[13],stage1_18[15],stage1_17[22]}
   );
   gpc623_5 gpc88 (
      {stage0_17[40], stage0_17[41], stage0_17[42]},
      {stage0_18[48], stage0_18[49]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[14],stage1_19[14],stage1_18[16],stage1_17[23]}
   );
   gpc615_5 gpc89 (
      {stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53], stage0_18[54]},
      {stage0_19[42]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[7],stage1_20[15],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc90 (
      {stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage0_19[43]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[8],stage1_20[16],stage1_19[16],stage1_18[18]}
   );
   gpc615_5 gpc91 (
      {stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[9],stage1_20[17],stage1_19[17]}
   );
   gpc615_5 gpc92 (
      {stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage0_20[13]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[3],stage1_21[10],stage1_20[18],stage1_19[18]}
   );
   gpc615_5 gpc93 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[4],stage1_21[11],stage1_20[19]}
   );
   gpc615_5 gpc94 (
      {stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[5],stage1_21[12],stage1_20[20]}
   );
   gpc615_5 gpc95 (
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[6],stage1_21[13],stage1_20[21]}
   );
   gpc615_5 gpc96 (
      {stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[7],stage1_21[14],stage1_20[22]}
   );
   gpc615_5 gpc97 (
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[8],stage1_21[15],stage1_20[23]}
   );
   gpc615_5 gpc98 (
      {stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[9],stage1_21[16],stage1_20[24]}
   );
   gpc615_5 gpc99 (
      {stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47], stage0_20[48]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[10],stage1_21[17],stage1_20[25]}
   );
   gpc606_5 gpc100 (
      {stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[7],stage1_23[9],stage1_22[11],stage1_21[18]}
   );
   gpc606_5 gpc101 (
      {stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[8],stage1_23[10],stage1_22[12],stage1_21[19]}
   );
   gpc606_5 gpc102 (
      {stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[9],stage1_23[11],stage1_22[13],stage1_21[20]}
   );
   gpc606_5 gpc103 (
      {stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[10],stage1_23[12],stage1_22[14],stage1_21[21]}
   );
   gpc606_5 gpc104 (
      {stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[11],stage1_23[13],stage1_22[15],stage1_21[22]}
   );
   gpc606_5 gpc105 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[12],stage1_23[14],stage1_22[16],stage1_21[23]}
   );
   gpc615_5 gpc106 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46]},
      {stage0_23[36]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[6],stage1_24[13],stage1_23[15],stage1_22[17]}
   );
   gpc615_5 gpc107 (
      {stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51]},
      {stage0_23[37]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[7],stage1_24[14],stage1_23[16],stage1_22[18]}
   );
   gpc615_5 gpc108 (
      {stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage0_24[12]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[2],stage1_25[8],stage1_24[15],stage1_23[17]}
   );
   gpc615_5 gpc109 (
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage0_24[13]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[3],stage1_25[9],stage1_24[16],stage1_23[18]}
   );
   gpc606_5 gpc110 (
      {stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18], stage0_24[19]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[4],stage1_25[10],stage1_24[17]}
   );
   gpc606_5 gpc111 (
      {stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24], stage0_24[25]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[5],stage1_25[11],stage1_24[18]}
   );
   gpc606_5 gpc112 (
      {stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[6],stage1_25[12],stage1_24[19]}
   );
   gpc606_5 gpc113 (
      {stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36], stage0_24[37]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[7],stage1_25[13],stage1_24[20]}
   );
   gpc606_5 gpc114 (
      {stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42], stage0_24[43]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[8],stage1_25[14],stage1_24[21]}
   );
   gpc606_5 gpc115 (
      {stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47], stage0_24[48], stage0_24[49]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[9],stage1_25[15],stage1_24[22]}
   );
   gpc606_5 gpc116 (
      {stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53], stage0_24[54], stage0_24[55]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[10],stage1_25[16],stage1_24[23]}
   );
   gpc606_5 gpc117 (
      {stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59], stage0_24[60], stage0_24[61]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[11],stage1_25[17],stage1_24[24]}
   );
   gpc606_5 gpc118 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[10],stage1_26[12],stage1_25[18]}
   );
   gpc606_5 gpc119 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[11],stage1_26[13],stage1_25[19]}
   );
   gpc606_5 gpc120 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[12],stage1_26[14],stage1_25[20]}
   );
   gpc606_5 gpc121 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[13],stage1_26[15],stage1_25[21]}
   );
   gpc606_5 gpc122 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[14],stage1_26[16],stage1_25[22]}
   );
   gpc615_5 gpc123 (
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52]},
      {stage0_27[30]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[5],stage1_28[13],stage1_27[15],stage1_26[17]}
   );
   gpc615_5 gpc124 (
      {stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage0_28[6]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[6],stage1_28[14],stage1_27[16]}
   );
   gpc615_5 gpc125 (
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40]},
      {stage0_28[7]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[2],stage1_29[7],stage1_28[15],stage1_27[17]}
   );
   gpc606_5 gpc126 (
      {stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[3],stage1_29[8],stage1_28[16]}
   );
   gpc606_5 gpc127 (
      {stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[3],stage1_30[4],stage1_29[9],stage1_28[17]}
   );
   gpc606_5 gpc128 (
      {stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[4],stage1_30[5],stage1_29[10],stage1_28[18]}
   );
   gpc606_5 gpc129 (
      {stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[5],stage1_30[6],stage1_29[11],stage1_28[19]}
   );
   gpc606_5 gpc130 (
      {stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36], stage0_28[37]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[6],stage1_30[7],stage1_29[12],stage1_28[20]}
   );
   gpc606_5 gpc131 (
      {stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42], stage0_28[43]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[7],stage1_30[8],stage1_29[13],stage1_28[21]}
   );
   gpc606_5 gpc132 (
      {stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48], stage0_28[49]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[8],stage1_30[9],stage1_29[14],stage1_28[22]}
   );
   gpc606_5 gpc133 (
      {stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], stage0_28[54], stage0_28[55]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[9],stage1_30[10],stage1_29[15],stage1_28[23]}
   );
   gpc606_5 gpc134 (
      {stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59], stage0_28[60], stage0_28[61]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[10],stage1_30[11],stage1_29[16],stage1_28[24]}
   );
   gpc606_5 gpc135 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[11],stage1_30[12],stage1_29[17]}
   );
   gpc606_5 gpc136 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[12],stage1_30[13],stage1_29[18]}
   );
   gpc606_5 gpc137 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[13],stage1_30[14],stage1_29[19]}
   );
   gpc606_5 gpc138 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[14],stage1_30[15],stage1_29[20]}
   );
   gpc606_5 gpc139 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[15],stage1_30[16],stage1_29[21]}
   );
   gpc606_5 gpc140 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[16],stage1_30[17],stage1_29[22]}
   );
   gpc606_5 gpc141 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[17],stage1_30[18],stage1_29[23]}
   );
   gpc606_5 gpc142 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[18],stage1_30[19],stage1_29[24]}
   );
   gpc615_5 gpc143 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58]},
      {stage0_31[48]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[8],stage1_32[17],stage1_31[19],stage1_30[20]}
   );
   gpc615_5 gpc144 (
      {stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage0_32[6]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[1],stage1_33[9],stage1_32[18],stage1_31[20]}
   );
   gpc615_5 gpc145 (
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58]},
      {stage0_32[7]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[2],stage1_33[10],stage1_32[19],stage1_31[21]}
   );
   gpc615_5 gpc146 (
      {stage0_31[59], stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63]},
      {stage0_32[8]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[3],stage1_33[11],stage1_32[20],stage1_31[22]}
   );
   gpc606_5 gpc147 (
      {stage0_32[9], stage0_32[10], stage0_32[11], stage0_32[12], stage0_32[13], stage0_32[14]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[3],stage1_34[4],stage1_33[12],stage1_32[21]}
   );
   gpc606_5 gpc148 (
      {stage0_32[15], stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[4],stage1_34[5],stage1_33[13],stage1_32[22]}
   );
   gpc606_5 gpc149 (
      {stage0_32[21], stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[5],stage1_34[6],stage1_33[14],stage1_32[23]}
   );
   gpc606_5 gpc150 (
      {stage0_32[27], stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[6],stage1_34[7],stage1_33[15],stage1_32[24]}
   );
   gpc606_5 gpc151 (
      {stage0_32[33], stage0_32[34], stage0_32[35], stage0_32[36], stage0_32[37], stage0_32[38]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[7],stage1_34[8],stage1_33[16],stage1_32[25]}
   );
   gpc606_5 gpc152 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[8],stage1_34[9],stage1_33[17],stage1_32[26]}
   );
   gpc606_5 gpc153 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[9],stage1_34[10],stage1_33[18],stage1_32[27]}
   );
   gpc606_5 gpc154 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[10],stage1_34[11],stage1_33[19],stage1_32[28]}
   );
   gpc606_5 gpc155 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[11],stage1_34[12],stage1_33[20],stage1_32[29]}
   );
   gpc606_5 gpc156 (
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[9],stage1_35[12],stage1_34[13],stage1_33[21]}
   );
   gpc606_5 gpc157 (
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[10],stage1_35[13],stage1_34[14],stage1_33[22]}
   );
   gpc606_5 gpc158 (
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[11],stage1_35[14],stage1_34[15],stage1_33[23]}
   );
   gpc606_5 gpc159 (
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[12],stage1_35[15],stage1_34[16],stage1_33[24]}
   );
   gpc606_5 gpc160 (
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[13],stage1_35[16],stage1_34[17],stage1_33[25]}
   );
   gpc615_5 gpc161 (
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52]},
      {stage0_34[54]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[14],stage1_35[17],stage1_34[18],stage1_33[26]}
   );
   gpc615_5 gpc162 (
      {stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage0_35[36]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[6],stage1_36[15],stage1_35[18],stage1_34[19]}
   );
   gpc615_5 gpc163 (
      {stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage0_36[6]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[1],stage1_37[7],stage1_36[16],stage1_35[19]}
   );
   gpc615_5 gpc164 (
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46]},
      {stage0_36[7]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[2],stage1_37[8],stage1_36[17],stage1_35[20]}
   );
   gpc615_5 gpc165 (
      {stage0_35[47], stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51]},
      {stage0_36[8]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[3],stage1_37[9],stage1_36[18],stage1_35[21]}
   );
   gpc615_5 gpc166 (
      {stage0_35[52], stage0_35[53], stage0_35[54], stage0_35[55], stage0_35[56]},
      {stage0_36[9]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[4],stage1_37[10],stage1_36[19],stage1_35[22]}
   );
   gpc606_5 gpc167 (
      {stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[4],stage1_38[5],stage1_37[11],stage1_36[20]}
   );
   gpc606_5 gpc168 (
      {stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[5],stage1_38[6],stage1_37[12],stage1_36[21]}
   );
   gpc606_5 gpc169 (
      {stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[6],stage1_38[7],stage1_37[13],stage1_36[22]}
   );
   gpc606_5 gpc170 (
      {stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[7],stage1_38[8],stage1_37[14],stage1_36[23]}
   );
   gpc606_5 gpc171 (
      {stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[8],stage1_38[9],stage1_37[15],stage1_36[24]}
   );
   gpc606_5 gpc172 (
      {stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[9],stage1_38[10],stage1_37[16],stage1_36[25]}
   );
   gpc606_5 gpc173 (
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[10],stage1_38[11],stage1_37[17]}
   );
   gpc606_5 gpc174 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[11],stage1_38[12],stage1_37[18]}
   );
   gpc606_5 gpc175 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[12],stage1_38[13],stage1_37[19]}
   );
   gpc606_5 gpc176 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[9],stage1_39[13],stage1_38[14],stage1_37[20]}
   );
   gpc606_5 gpc177 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[10],stage1_39[14],stage1_38[15],stage1_37[21]}
   );
   gpc606_5 gpc178 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[11],stage1_39[15],stage1_38[16],stage1_37[22]}
   );
   gpc606_5 gpc179 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], 1'b0, 1'b0},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[12],stage1_39[16],stage1_38[17],stage1_37[23]}
   );
   gpc615_5 gpc180 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[13],stage1_39[17],stage1_38[18]}
   );
   gpc615_5 gpc181 (
      {stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage0_40[6]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[8],stage1_40[14],stage1_39[18]}
   );
   gpc615_5 gpc182 (
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52]},
      {stage0_40[7]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[2],stage1_41[9],stage1_40[15],stage1_39[19]}
   );
   gpc615_5 gpc183 (
      {stage0_39[53], stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57]},
      {stage0_40[8]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[3],stage1_41[10],stage1_40[16],stage1_39[20]}
   );
   gpc615_5 gpc184 (
      {stage0_39[58], stage0_39[59], stage0_39[60], stage0_39[61], stage0_39[62]},
      {stage0_40[9]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[4],stage1_41[11],stage1_40[17],stage1_39[21]}
   );
   gpc606_5 gpc185 (
      {stage0_40[10], stage0_40[11], stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[4],stage1_42[5],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc186 (
      {stage0_40[16], stage0_40[17], stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[5],stage1_42[6],stage1_41[13],stage1_40[19]}
   );
   gpc606_5 gpc187 (
      {stage0_40[22], stage0_40[23], stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[6],stage1_42[7],stage1_41[14],stage1_40[20]}
   );
   gpc606_5 gpc188 (
      {stage0_40[28], stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[7],stage1_42[8],stage1_41[15],stage1_40[21]}
   );
   gpc606_5 gpc189 (
      {stage0_40[34], stage0_40[35], stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[8],stage1_42[9],stage1_41[16],stage1_40[22]}
   );
   gpc606_5 gpc190 (
      {stage0_40[40], stage0_40[41], stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[9],stage1_42[10],stage1_41[17],stage1_40[23]}
   );
   gpc606_5 gpc191 (
      {stage0_40[46], stage0_40[47], stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[10],stage1_42[11],stage1_41[18],stage1_40[24]}
   );
   gpc606_5 gpc192 (
      {stage0_40[52], stage0_40[53], stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[11],stage1_42[12],stage1_41[19],stage1_40[25]}
   );
   gpc606_5 gpc193 (
      {stage0_40[58], stage0_40[59], stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[12],stage1_42[13],stage1_41[20],stage1_40[26]}
   );
   gpc606_5 gpc194 (
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[9],stage1_43[13],stage1_42[14],stage1_41[21]}
   );
   gpc606_5 gpc195 (
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[10],stage1_43[14],stage1_42[15],stage1_41[22]}
   );
   gpc606_5 gpc196 (
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[11],stage1_43[15],stage1_42[16],stage1_41[23]}
   );
   gpc606_5 gpc197 (
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[12],stage1_43[16],stage1_42[17],stage1_41[24]}
   );
   gpc606_5 gpc198 (
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[13],stage1_43[17],stage1_42[18],stage1_41[25]}
   );
   gpc615_5 gpc199 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[0]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[0],stage1_45[5],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc200 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[1]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[1],stage1_45[6],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc201 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[2]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[2],stage1_45[7],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc202 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[3]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[3],stage1_45[8],stage1_44[17],stage1_43[21]}
   );
   gpc606_5 gpc203 (
      {stage0_44[4], stage0_44[5], stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[4],stage1_46[4],stage1_45[9],stage1_44[18]}
   );
   gpc606_5 gpc204 (
      {stage0_44[10], stage0_44[11], stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[5],stage1_46[5],stage1_45[10],stage1_44[19]}
   );
   gpc606_5 gpc205 (
      {stage0_44[16], stage0_44[17], stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[6],stage1_46[6],stage1_45[11],stage1_44[20]}
   );
   gpc606_5 gpc206 (
      {stage0_44[22], stage0_44[23], stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[7],stage1_46[7],stage1_45[12],stage1_44[21]}
   );
   gpc606_5 gpc207 (
      {stage0_44[28], stage0_44[29], stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[8],stage1_46[8],stage1_45[13],stage1_44[22]}
   );
   gpc606_5 gpc208 (
      {stage0_44[34], stage0_44[35], stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[9],stage1_46[9],stage1_45[14],stage1_44[23]}
   );
   gpc606_5 gpc209 (
      {stage0_44[40], stage0_44[41], stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[10],stage1_46[10],stage1_45[15],stage1_44[24]}
   );
   gpc606_5 gpc210 (
      {stage0_44[46], stage0_44[47], stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[11],stage1_46[11],stage1_45[16],stage1_44[25]}
   );
   gpc606_5 gpc211 (
      {stage0_44[52], stage0_44[53], stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[12],stage1_46[12],stage1_45[17],stage1_44[26]}
   );
   gpc606_5 gpc212 (
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[9],stage1_47[13],stage1_46[13],stage1_45[18]}
   );
   gpc606_5 gpc213 (
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[10],stage1_47[14],stage1_46[14],stage1_45[19]}
   );
   gpc615_5 gpc214 (
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58]},
      {stage0_47[12]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[2],stage1_48[11],stage1_47[15],stage1_46[15]}
   );
   gpc615_5 gpc215 (
      {stage0_46[59], stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63]},
      {stage0_47[13]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[3],stage1_48[12],stage1_47[16],stage1_46[16]}
   );
   gpc606_5 gpc216 (
      {stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[2],stage1_49[4],stage1_48[13],stage1_47[17]}
   );
   gpc606_5 gpc217 (
      {stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[3],stage1_49[5],stage1_48[14],stage1_47[18]}
   );
   gpc615_5 gpc218 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[12]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[4],stage1_49[6],stage1_48[15],stage1_47[19]}
   );
   gpc615_5 gpc219 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[13]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[5],stage1_49[7],stage1_48[16],stage1_47[20]}
   );
   gpc615_5 gpc220 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[14]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[6],stage1_49[8],stage1_48[17],stage1_47[21]}
   );
   gpc615_5 gpc221 (
      {stage0_47[41], stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45]},
      {stage0_48[15]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[7],stage1_49[9],stage1_48[18],stage1_47[22]}
   );
   gpc606_5 gpc222 (
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[8],stage1_49[10],stage1_48[19]}
   );
   gpc606_5 gpc223 (
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[9],stage1_49[11],stage1_48[20]}
   );
   gpc606_5 gpc224 (
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[10],stage1_49[12],stage1_48[21]}
   );
   gpc606_5 gpc225 (
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[9],stage1_50[11],stage1_49[13],stage1_48[22]}
   );
   gpc606_5 gpc226 (
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[10],stage1_50[12],stage1_49[14],stage1_48[23]}
   );
   gpc606_5 gpc227 (
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[11],stage1_50[13],stage1_49[15],stage1_48[24]}
   );
   gpc606_5 gpc228 (
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[12],stage1_50[14],stage1_49[16],stage1_48[25]}
   );
   gpc606_5 gpc229 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[7],stage1_51[13],stage1_50[15],stage1_49[17]}
   );
   gpc606_5 gpc230 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[8],stage1_51[14],stage1_50[16],stage1_49[18]}
   );
   gpc606_5 gpc231 (
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[9],stage1_51[15],stage1_50[17],stage1_49[19]}
   );
   gpc606_5 gpc232 (
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[10],stage1_51[16],stage1_50[18],stage1_49[20]}
   );
   gpc615_5 gpc233 (
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46]},
      {stage0_51[24]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[4],stage1_52[11],stage1_51[17],stage1_50[19]}
   );
   gpc615_5 gpc234 (
      {stage0_50[47], stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51]},
      {stage0_51[25]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[5],stage1_52[12],stage1_51[18],stage1_50[20]}
   );
   gpc615_5 gpc235 (
      {stage0_50[52], stage0_50[53], stage0_50[54], stage0_50[55], stage0_50[56]},
      {stage0_51[26]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[6],stage1_52[13],stage1_51[19],stage1_50[21]}
   );
   gpc615_5 gpc236 (
      {stage0_50[57], stage0_50[58], stage0_50[59], stage0_50[60], stage0_50[61]},
      {stage0_51[27]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[7],stage1_52[14],stage1_51[20],stage1_50[22]}
   );
   gpc606_5 gpc237 (
      {stage0_51[28], stage0_51[29], stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[8],stage1_52[15],stage1_51[21]}
   );
   gpc615_5 gpc238 (
      {stage0_51[34], stage0_51[35], stage0_51[36], stage0_51[37], stage0_51[38]},
      {stage0_52[24]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[9],stage1_52[16],stage1_51[22]}
   );
   gpc615_5 gpc239 (
      {stage0_51[39], stage0_51[40], stage0_51[41], stage0_51[42], stage0_51[43]},
      {stage0_52[25]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[10],stage1_52[17],stage1_51[23]}
   );
   gpc615_5 gpc240 (
      {stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47], stage0_51[48]},
      {stage0_52[26]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[11],stage1_52[18],stage1_51[24]}
   );
   gpc615_5 gpc241 (
      {stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage0_52[27]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[12],stage1_52[19],stage1_51[25]}
   );
   gpc615_5 gpc242 (
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58]},
      {stage0_52[28]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[13],stage1_52[20],stage1_51[26]}
   );
   gpc606_5 gpc243 (
      {stage0_52[29], stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[6],stage1_54[10],stage1_53[14],stage1_52[21]}
   );
   gpc615_5 gpc244 (
      {stage0_52[35], stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39]},
      {stage0_53[36]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[7],stage1_54[11],stage1_53[15],stage1_52[22]}
   );
   gpc615_5 gpc245 (
      {stage0_52[40], stage0_52[41], stage0_52[42], stage0_52[43], stage0_52[44]},
      {stage0_53[37]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[8],stage1_54[12],stage1_53[16],stage1_52[23]}
   );
   gpc615_5 gpc246 (
      {stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41], stage0_53[42]},
      {stage0_54[18]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[3],stage1_55[9],stage1_54[13],stage1_53[17]}
   );
   gpc615_5 gpc247 (
      {stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage0_54[19]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[4],stage1_55[10],stage1_54[14],stage1_53[18]}
   );
   gpc615_5 gpc248 (
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52]},
      {stage0_54[20]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[5],stage1_55[11],stage1_54[15],stage1_53[19]}
   );
   gpc615_5 gpc249 (
      {stage0_53[53], stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57]},
      {stage0_54[21]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[6],stage1_55[12],stage1_54[16],stage1_53[20]}
   );
   gpc606_5 gpc250 (
      {stage0_54[22], stage0_54[23], stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[4],stage1_56[7],stage1_55[13],stage1_54[17]}
   );
   gpc606_5 gpc251 (
      {stage0_54[28], stage0_54[29], stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[5],stage1_56[8],stage1_55[14],stage1_54[18]}
   );
   gpc615_5 gpc252 (
      {stage0_54[34], stage0_54[35], stage0_54[36], stage0_54[37], stage0_54[38]},
      {stage0_55[24]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[6],stage1_56[9],stage1_55[15],stage1_54[19]}
   );
   gpc615_5 gpc253 (
      {stage0_54[39], stage0_54[40], stage0_54[41], stage0_54[42], stage0_54[43]},
      {stage0_55[25]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[7],stage1_56[10],stage1_55[16],stage1_54[20]}
   );
   gpc615_5 gpc254 (
      {stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48]},
      {stage0_55[26]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[8],stage1_56[11],stage1_55[17],stage1_54[21]}
   );
   gpc615_5 gpc255 (
      {stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage0_55[27]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[9],stage1_56[12],stage1_55[18],stage1_54[22]}
   );
   gpc606_5 gpc256 (
      {stage0_55[28], stage0_55[29], stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[10],stage1_56[13],stage1_55[19]}
   );
   gpc606_5 gpc257 (
      {stage0_55[34], stage0_55[35], stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[11],stage1_56[14],stage1_55[20]}
   );
   gpc606_5 gpc258 (
      {stage0_55[40], stage0_55[41], stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[12],stage1_56[15],stage1_55[21]}
   );
   gpc606_5 gpc259 (
      {stage0_55[46], stage0_55[47], stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[13],stage1_56[16],stage1_55[22]}
   );
   gpc606_5 gpc260 (
      {stage0_55[52], stage0_55[53], stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[10],stage1_57[14],stage1_56[17],stage1_55[23]}
   );
   gpc606_5 gpc261 (
      {stage0_55[58], stage0_55[59], stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[11],stage1_57[15],stage1_56[18],stage1_55[24]}
   );
   gpc606_5 gpc262 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[6],stage1_58[12],stage1_57[16],stage1_56[19]}
   );
   gpc615_5 gpc263 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46]},
      {stage0_57[36]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[7],stage1_58[13],stage1_57[17],stage1_56[20]}
   );
   gpc615_5 gpc264 (
      {stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_57[37]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[8],stage1_58[14],stage1_57[18],stage1_56[21]}
   );
   gpc615_5 gpc265 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56]},
      {stage0_57[38]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[9],stage1_58[15],stage1_57[19],stage1_56[22]}
   );
   gpc615_5 gpc266 (
      {stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_57[39]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[10],stage1_58[16],stage1_57[20],stage1_56[23]}
   );
   gpc615_5 gpc267 (
      {stage0_57[40], stage0_57[41], stage0_57[42], stage0_57[43], stage0_57[44]},
      {stage0_58[30]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[5],stage1_59[11],stage1_58[17],stage1_57[21]}
   );
   gpc615_5 gpc268 (
      {stage0_57[45], stage0_57[46], stage0_57[47], stage0_57[48], stage0_57[49]},
      {stage0_58[31]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[6],stage1_59[12],stage1_58[18],stage1_57[22]}
   );
   gpc615_5 gpc269 (
      {stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53], stage0_57[54]},
      {stage0_58[32]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[7],stage1_59[13],stage1_58[19],stage1_57[23]}
   );
   gpc615_5 gpc270 (
      {stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_58[33]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[8],stage1_59[14],stage1_58[20],stage1_57[24]}
   );
   gpc615_5 gpc271 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], 1'b0},
      {stage0_58[34]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[9],stage1_59[15],stage1_58[21],stage1_57[25]}
   );
   gpc1406_5 gpc272 (
      {stage0_58[35], stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3]},
      {stage0_61[0]},
      {stage1_62[0],stage1_61[5],stage1_60[10],stage1_59[16],stage1_58[22]}
   );
   gpc606_5 gpc273 (
      {stage0_58[41], stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46]},
      {stage0_60[4], stage0_60[5], stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9]},
      {stage1_62[1],stage1_61[6],stage1_60[11],stage1_59[17],stage1_58[23]}
   );
   gpc606_5 gpc274 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5], stage0_61[6]},
      {stage1_63[0],stage1_62[2],stage1_61[7],stage1_60[12],stage1_59[18]}
   );
   gpc606_5 gpc275 (
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11], stage0_61[12]},
      {stage1_63[1],stage1_62[3],stage1_61[8],stage1_60[13],stage1_59[19]}
   );
   gpc606_5 gpc276 (
      {stage0_60[10], stage0_60[11], stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[2],stage1_62[4],stage1_61[9],stage1_60[14]}
   );
   gpc606_5 gpc277 (
      {stage0_60[16], stage0_60[17], stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[3],stage1_62[5],stage1_61[10],stage1_60[15]}
   );
   gpc606_5 gpc278 (
      {stage0_60[22], stage0_60[23], stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[4],stage1_62[6],stage1_61[11],stage1_60[16]}
   );
   gpc606_5 gpc279 (
      {stage0_60[28], stage0_60[29], stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[5],stage1_62[7],stage1_61[12],stage1_60[17]}
   );
   gpc606_5 gpc280 (
      {stage0_60[34], stage0_60[35], stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[6],stage1_62[8],stage1_61[13],stage1_60[18]}
   );
   gpc606_5 gpc281 (
      {stage0_60[40], stage0_60[41], stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[7],stage1_62[9],stage1_61[14],stage1_60[19]}
   );
   gpc606_5 gpc282 (
      {stage0_60[46], stage0_60[47], stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[8],stage1_62[10],stage1_61[15],stage1_60[20]}
   );
   gpc615_5 gpc283 (
      {stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_62[42]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[7],stage1_63[9],stage1_62[11],stage1_61[16]}
   );
   gpc615_5 gpc284 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22]},
      {stage0_62[43]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[8],stage1_63[10],stage1_62[12],stage1_61[17]}
   );
   gpc615_5 gpc285 (
      {stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27]},
      {stage0_62[44]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[9],stage1_63[11],stage1_62[13],stage1_61[18]}
   );
   gpc615_5 gpc286 (
      {stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage0_62[45]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[10],stage1_63[12],stage1_62[14],stage1_61[19]}
   );
   gpc615_5 gpc287 (
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37]},
      {stage0_62[46]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[11],stage1_63[13],stage1_62[15],stage1_61[20]}
   );
   gpc615_5 gpc288 (
      {stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42]},
      {stage0_62[47]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[12],stage1_63[14],stage1_62[16],stage1_61[21]}
   );
   gpc615_5 gpc289 (
      {stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_62[48]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[13],stage1_63[15],stage1_62[17],stage1_61[22]}
   );
   gpc615_5 gpc290 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52]},
      {stage0_62[49]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[14],stage1_63[16],stage1_62[18],stage1_61[23]}
   );
   gpc615_5 gpc291 (
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57]},
      {stage0_62[50]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[15],stage1_63[17],stage1_62[19],stage1_61[24]}
   );
   gpc1_1 gpc292 (
      {stage0_0[54]},
      {stage1_0[9]}
   );
   gpc1_1 gpc293 (
      {stage0_0[55]},
      {stage1_0[10]}
   );
   gpc1_1 gpc294 (
      {stage0_0[56]},
      {stage1_0[11]}
   );
   gpc1_1 gpc295 (
      {stage0_0[57]},
      {stage1_0[12]}
   );
   gpc1_1 gpc296 (
      {stage0_0[58]},
      {stage1_0[13]}
   );
   gpc1_1 gpc297 (
      {stage0_0[59]},
      {stage1_0[14]}
   );
   gpc1_1 gpc298 (
      {stage0_0[60]},
      {stage1_0[15]}
   );
   gpc1_1 gpc299 (
      {stage0_0[61]},
      {stage1_0[16]}
   );
   gpc1_1 gpc300 (
      {stage0_0[62]},
      {stage1_0[17]}
   );
   gpc1_1 gpc301 (
      {stage0_0[63]},
      {stage1_0[18]}
   );
   gpc1_1 gpc302 (
      {stage0_1[30]},
      {stage1_1[14]}
   );
   gpc1_1 gpc303 (
      {stage0_1[31]},
      {stage1_1[15]}
   );
   gpc1_1 gpc304 (
      {stage0_1[32]},
      {stage1_1[16]}
   );
   gpc1_1 gpc305 (
      {stage0_1[33]},
      {stage1_1[17]}
   );
   gpc1_1 gpc306 (
      {stage0_1[34]},
      {stage1_1[18]}
   );
   gpc1_1 gpc307 (
      {stage0_1[35]},
      {stage1_1[19]}
   );
   gpc1_1 gpc308 (
      {stage0_1[36]},
      {stage1_1[20]}
   );
   gpc1_1 gpc309 (
      {stage0_1[37]},
      {stage1_1[21]}
   );
   gpc1_1 gpc310 (
      {stage0_1[38]},
      {stage1_1[22]}
   );
   gpc1_1 gpc311 (
      {stage0_1[39]},
      {stage1_1[23]}
   );
   gpc1_1 gpc312 (
      {stage0_1[40]},
      {stage1_1[24]}
   );
   gpc1_1 gpc313 (
      {stage0_1[41]},
      {stage1_1[25]}
   );
   gpc1_1 gpc314 (
      {stage0_1[42]},
      {stage1_1[26]}
   );
   gpc1_1 gpc315 (
      {stage0_1[43]},
      {stage1_1[27]}
   );
   gpc1_1 gpc316 (
      {stage0_1[44]},
      {stage1_1[28]}
   );
   gpc1_1 gpc317 (
      {stage0_1[45]},
      {stage1_1[29]}
   );
   gpc1_1 gpc318 (
      {stage0_1[46]},
      {stage1_1[30]}
   );
   gpc1_1 gpc319 (
      {stage0_1[47]},
      {stage1_1[31]}
   );
   gpc1_1 gpc320 (
      {stage0_1[48]},
      {stage1_1[32]}
   );
   gpc1_1 gpc321 (
      {stage0_1[49]},
      {stage1_1[33]}
   );
   gpc1_1 gpc322 (
      {stage0_1[50]},
      {stage1_1[34]}
   );
   gpc1_1 gpc323 (
      {stage0_1[51]},
      {stage1_1[35]}
   );
   gpc1_1 gpc324 (
      {stage0_1[52]},
      {stage1_1[36]}
   );
   gpc1_1 gpc325 (
      {stage0_1[53]},
      {stage1_1[37]}
   );
   gpc1_1 gpc326 (
      {stage0_1[54]},
      {stage1_1[38]}
   );
   gpc1_1 gpc327 (
      {stage0_1[55]},
      {stage1_1[39]}
   );
   gpc1_1 gpc328 (
      {stage0_1[56]},
      {stage1_1[40]}
   );
   gpc1_1 gpc329 (
      {stage0_1[57]},
      {stage1_1[41]}
   );
   gpc1_1 gpc330 (
      {stage0_1[58]},
      {stage1_1[42]}
   );
   gpc1_1 gpc331 (
      {stage0_1[59]},
      {stage1_1[43]}
   );
   gpc1_1 gpc332 (
      {stage0_1[60]},
      {stage1_1[44]}
   );
   gpc1_1 gpc333 (
      {stage0_1[61]},
      {stage1_1[45]}
   );
   gpc1_1 gpc334 (
      {stage0_1[62]},
      {stage1_1[46]}
   );
   gpc1_1 gpc335 (
      {stage0_1[63]},
      {stage1_1[47]}
   );
   gpc1_1 gpc336 (
      {stage0_2[54]},
      {stage1_2[14]}
   );
   gpc1_1 gpc337 (
      {stage0_2[55]},
      {stage1_2[15]}
   );
   gpc1_1 gpc338 (
      {stage0_2[56]},
      {stage1_2[16]}
   );
   gpc1_1 gpc339 (
      {stage0_2[57]},
      {stage1_2[17]}
   );
   gpc1_1 gpc340 (
      {stage0_2[58]},
      {stage1_2[18]}
   );
   gpc1_1 gpc341 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc342 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc343 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc344 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc345 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc346 (
      {stage0_3[55]},
      {stage1_3[19]}
   );
   gpc1_1 gpc347 (
      {stage0_3[56]},
      {stage1_3[20]}
   );
   gpc1_1 gpc348 (
      {stage0_3[57]},
      {stage1_3[21]}
   );
   gpc1_1 gpc349 (
      {stage0_3[58]},
      {stage1_3[22]}
   );
   gpc1_1 gpc350 (
      {stage0_3[59]},
      {stage1_3[23]}
   );
   gpc1_1 gpc351 (
      {stage0_3[60]},
      {stage1_3[24]}
   );
   gpc1_1 gpc352 (
      {stage0_3[61]},
      {stage1_3[25]}
   );
   gpc1_1 gpc353 (
      {stage0_3[62]},
      {stage1_3[26]}
   );
   gpc1_1 gpc354 (
      {stage0_3[63]},
      {stage1_3[27]}
   );
   gpc1_1 gpc355 (
      {stage0_4[53]},
      {stage1_4[27]}
   );
   gpc1_1 gpc356 (
      {stage0_4[54]},
      {stage1_4[28]}
   );
   gpc1_1 gpc357 (
      {stage0_4[55]},
      {stage1_4[29]}
   );
   gpc1_1 gpc358 (
      {stage0_4[56]},
      {stage1_4[30]}
   );
   gpc1_1 gpc359 (
      {stage0_4[57]},
      {stage1_4[31]}
   );
   gpc1_1 gpc360 (
      {stage0_4[58]},
      {stage1_4[32]}
   );
   gpc1_1 gpc361 (
      {stage0_4[59]},
      {stage1_4[33]}
   );
   gpc1_1 gpc362 (
      {stage0_4[60]},
      {stage1_4[34]}
   );
   gpc1_1 gpc363 (
      {stage0_4[61]},
      {stage1_4[35]}
   );
   gpc1_1 gpc364 (
      {stage0_4[62]},
      {stage1_4[36]}
   );
   gpc1_1 gpc365 (
      {stage0_4[63]},
      {stage1_4[37]}
   );
   gpc1_1 gpc366 (
      {stage0_5[60]},
      {stage1_5[23]}
   );
   gpc1_1 gpc367 (
      {stage0_5[61]},
      {stage1_5[24]}
   );
   gpc1_1 gpc368 (
      {stage0_5[62]},
      {stage1_5[25]}
   );
   gpc1_1 gpc369 (
      {stage0_5[63]},
      {stage1_5[26]}
   );
   gpc1_1 gpc370 (
      {stage0_6[63]},
      {stage1_6[21]}
   );
   gpc1_1 gpc371 (
      {stage0_7[53]},
      {stage1_7[25]}
   );
   gpc1_1 gpc372 (
      {stage0_7[54]},
      {stage1_7[26]}
   );
   gpc1_1 gpc373 (
      {stage0_7[55]},
      {stage1_7[27]}
   );
   gpc1_1 gpc374 (
      {stage0_7[56]},
      {stage1_7[28]}
   );
   gpc1_1 gpc375 (
      {stage0_7[57]},
      {stage1_7[29]}
   );
   gpc1_1 gpc376 (
      {stage0_7[58]},
      {stage1_7[30]}
   );
   gpc1_1 gpc377 (
      {stage0_7[59]},
      {stage1_7[31]}
   );
   gpc1_1 gpc378 (
      {stage0_7[60]},
      {stage1_7[32]}
   );
   gpc1_1 gpc379 (
      {stage0_7[61]},
      {stage1_7[33]}
   );
   gpc1_1 gpc380 (
      {stage0_7[62]},
      {stage1_7[34]}
   );
   gpc1_1 gpc381 (
      {stage0_7[63]},
      {stage1_7[35]}
   );
   gpc1_1 gpc382 (
      {stage0_9[60]},
      {stage1_9[25]}
   );
   gpc1_1 gpc383 (
      {stage0_9[61]},
      {stage1_9[26]}
   );
   gpc1_1 gpc384 (
      {stage0_9[62]},
      {stage1_9[27]}
   );
   gpc1_1 gpc385 (
      {stage0_9[63]},
      {stage1_9[28]}
   );
   gpc1_1 gpc386 (
      {stage0_10[52]},
      {stage1_10[22]}
   );
   gpc1_1 gpc387 (
      {stage0_10[53]},
      {stage1_10[23]}
   );
   gpc1_1 gpc388 (
      {stage0_10[54]},
      {stage1_10[24]}
   );
   gpc1_1 gpc389 (
      {stage0_10[55]},
      {stage1_10[25]}
   );
   gpc1_1 gpc390 (
      {stage0_10[56]},
      {stage1_10[26]}
   );
   gpc1_1 gpc391 (
      {stage0_10[57]},
      {stage1_10[27]}
   );
   gpc1_1 gpc392 (
      {stage0_10[58]},
      {stage1_10[28]}
   );
   gpc1_1 gpc393 (
      {stage0_10[59]},
      {stage1_10[29]}
   );
   gpc1_1 gpc394 (
      {stage0_10[60]},
      {stage1_10[30]}
   );
   gpc1_1 gpc395 (
      {stage0_10[61]},
      {stage1_10[31]}
   );
   gpc1_1 gpc396 (
      {stage0_10[62]},
      {stage1_10[32]}
   );
   gpc1_1 gpc397 (
      {stage0_10[63]},
      {stage1_10[33]}
   );
   gpc1_1 gpc398 (
      {stage0_11[53]},
      {stage1_11[22]}
   );
   gpc1_1 gpc399 (
      {stage0_11[54]},
      {stage1_11[23]}
   );
   gpc1_1 gpc400 (
      {stage0_11[55]},
      {stage1_11[24]}
   );
   gpc1_1 gpc401 (
      {stage0_11[56]},
      {stage1_11[25]}
   );
   gpc1_1 gpc402 (
      {stage0_11[57]},
      {stage1_11[26]}
   );
   gpc1_1 gpc403 (
      {stage0_11[58]},
      {stage1_11[27]}
   );
   gpc1_1 gpc404 (
      {stage0_11[59]},
      {stage1_11[28]}
   );
   gpc1_1 gpc405 (
      {stage0_11[60]},
      {stage1_11[29]}
   );
   gpc1_1 gpc406 (
      {stage0_11[61]},
      {stage1_11[30]}
   );
   gpc1_1 gpc407 (
      {stage0_11[62]},
      {stage1_11[31]}
   );
   gpc1_1 gpc408 (
      {stage0_11[63]},
      {stage1_11[32]}
   );
   gpc1_1 gpc409 (
      {stage0_12[63]},
      {stage1_12[26]}
   );
   gpc1_1 gpc410 (
      {stage0_13[59]},
      {stage1_13[26]}
   );
   gpc1_1 gpc411 (
      {stage0_13[60]},
      {stage1_13[27]}
   );
   gpc1_1 gpc412 (
      {stage0_13[61]},
      {stage1_13[28]}
   );
   gpc1_1 gpc413 (
      {stage0_13[62]},
      {stage1_13[29]}
   );
   gpc1_1 gpc414 (
      {stage0_13[63]},
      {stage1_13[30]}
   );
   gpc1_1 gpc415 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc416 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc417 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc418 (
      {stage0_15[39]},
      {stage1_15[20]}
   );
   gpc1_1 gpc419 (
      {stage0_15[40]},
      {stage1_15[21]}
   );
   gpc1_1 gpc420 (
      {stage0_15[41]},
      {stage1_15[22]}
   );
   gpc1_1 gpc421 (
      {stage0_15[42]},
      {stage1_15[23]}
   );
   gpc1_1 gpc422 (
      {stage0_15[43]},
      {stage1_15[24]}
   );
   gpc1_1 gpc423 (
      {stage0_15[44]},
      {stage1_15[25]}
   );
   gpc1_1 gpc424 (
      {stage0_15[45]},
      {stage1_15[26]}
   );
   gpc1_1 gpc425 (
      {stage0_15[46]},
      {stage1_15[27]}
   );
   gpc1_1 gpc426 (
      {stage0_15[47]},
      {stage1_15[28]}
   );
   gpc1_1 gpc427 (
      {stage0_15[48]},
      {stage1_15[29]}
   );
   gpc1_1 gpc428 (
      {stage0_15[49]},
      {stage1_15[30]}
   );
   gpc1_1 gpc429 (
      {stage0_15[50]},
      {stage1_15[31]}
   );
   gpc1_1 gpc430 (
      {stage0_15[51]},
      {stage1_15[32]}
   );
   gpc1_1 gpc431 (
      {stage0_15[52]},
      {stage1_15[33]}
   );
   gpc1_1 gpc432 (
      {stage0_15[53]},
      {stage1_15[34]}
   );
   gpc1_1 gpc433 (
      {stage0_15[54]},
      {stage1_15[35]}
   );
   gpc1_1 gpc434 (
      {stage0_15[55]},
      {stage1_15[36]}
   );
   gpc1_1 gpc435 (
      {stage0_15[56]},
      {stage1_15[37]}
   );
   gpc1_1 gpc436 (
      {stage0_15[57]},
      {stage1_15[38]}
   );
   gpc1_1 gpc437 (
      {stage0_15[58]},
      {stage1_15[39]}
   );
   gpc1_1 gpc438 (
      {stage0_15[59]},
      {stage1_15[40]}
   );
   gpc1_1 gpc439 (
      {stage0_15[60]},
      {stage1_15[41]}
   );
   gpc1_1 gpc440 (
      {stage0_15[61]},
      {stage1_15[42]}
   );
   gpc1_1 gpc441 (
      {stage0_15[62]},
      {stage1_15[43]}
   );
   gpc1_1 gpc442 (
      {stage0_15[63]},
      {stage1_15[44]}
   );
   gpc1_1 gpc443 (
      {stage0_16[58]},
      {stage1_16[25]}
   );
   gpc1_1 gpc444 (
      {stage0_16[59]},
      {stage1_16[26]}
   );
   gpc1_1 gpc445 (
      {stage0_16[60]},
      {stage1_16[27]}
   );
   gpc1_1 gpc446 (
      {stage0_16[61]},
      {stage1_16[28]}
   );
   gpc1_1 gpc447 (
      {stage0_16[62]},
      {stage1_16[29]}
   );
   gpc1_1 gpc448 (
      {stage0_16[63]},
      {stage1_16[30]}
   );
   gpc1_1 gpc449 (
      {stage0_17[43]},
      {stage1_17[24]}
   );
   gpc1_1 gpc450 (
      {stage0_17[44]},
      {stage1_17[25]}
   );
   gpc1_1 gpc451 (
      {stage0_17[45]},
      {stage1_17[26]}
   );
   gpc1_1 gpc452 (
      {stage0_17[46]},
      {stage1_17[27]}
   );
   gpc1_1 gpc453 (
      {stage0_17[47]},
      {stage1_17[28]}
   );
   gpc1_1 gpc454 (
      {stage0_17[48]},
      {stage1_17[29]}
   );
   gpc1_1 gpc455 (
      {stage0_17[49]},
      {stage1_17[30]}
   );
   gpc1_1 gpc456 (
      {stage0_17[50]},
      {stage1_17[31]}
   );
   gpc1_1 gpc457 (
      {stage0_17[51]},
      {stage1_17[32]}
   );
   gpc1_1 gpc458 (
      {stage0_17[52]},
      {stage1_17[33]}
   );
   gpc1_1 gpc459 (
      {stage0_17[53]},
      {stage1_17[34]}
   );
   gpc1_1 gpc460 (
      {stage0_17[54]},
      {stage1_17[35]}
   );
   gpc1_1 gpc461 (
      {stage0_17[55]},
      {stage1_17[36]}
   );
   gpc1_1 gpc462 (
      {stage0_17[56]},
      {stage1_17[37]}
   );
   gpc1_1 gpc463 (
      {stage0_17[57]},
      {stage1_17[38]}
   );
   gpc1_1 gpc464 (
      {stage0_17[58]},
      {stage1_17[39]}
   );
   gpc1_1 gpc465 (
      {stage0_17[59]},
      {stage1_17[40]}
   );
   gpc1_1 gpc466 (
      {stage0_17[60]},
      {stage1_17[41]}
   );
   gpc1_1 gpc467 (
      {stage0_17[61]},
      {stage1_17[42]}
   );
   gpc1_1 gpc468 (
      {stage0_17[62]},
      {stage1_17[43]}
   );
   gpc1_1 gpc469 (
      {stage0_17[63]},
      {stage1_17[44]}
   );
   gpc1_1 gpc470 (
      {stage0_18[60]},
      {stage1_18[19]}
   );
   gpc1_1 gpc471 (
      {stage0_18[61]},
      {stage1_18[20]}
   );
   gpc1_1 gpc472 (
      {stage0_18[62]},
      {stage1_18[21]}
   );
   gpc1_1 gpc473 (
      {stage0_18[63]},
      {stage1_18[22]}
   );
   gpc1_1 gpc474 (
      {stage0_19[54]},
      {stage1_19[19]}
   );
   gpc1_1 gpc475 (
      {stage0_19[55]},
      {stage1_19[20]}
   );
   gpc1_1 gpc476 (
      {stage0_19[56]},
      {stage1_19[21]}
   );
   gpc1_1 gpc477 (
      {stage0_19[57]},
      {stage1_19[22]}
   );
   gpc1_1 gpc478 (
      {stage0_19[58]},
      {stage1_19[23]}
   );
   gpc1_1 gpc479 (
      {stage0_19[59]},
      {stage1_19[24]}
   );
   gpc1_1 gpc480 (
      {stage0_19[60]},
      {stage1_19[25]}
   );
   gpc1_1 gpc481 (
      {stage0_19[61]},
      {stage1_19[26]}
   );
   gpc1_1 gpc482 (
      {stage0_19[62]},
      {stage1_19[27]}
   );
   gpc1_1 gpc483 (
      {stage0_19[63]},
      {stage1_19[28]}
   );
   gpc1_1 gpc484 (
      {stage0_20[49]},
      {stage1_20[26]}
   );
   gpc1_1 gpc485 (
      {stage0_20[50]},
      {stage1_20[27]}
   );
   gpc1_1 gpc486 (
      {stage0_20[51]},
      {stage1_20[28]}
   );
   gpc1_1 gpc487 (
      {stage0_20[52]},
      {stage1_20[29]}
   );
   gpc1_1 gpc488 (
      {stage0_20[53]},
      {stage1_20[30]}
   );
   gpc1_1 gpc489 (
      {stage0_20[54]},
      {stage1_20[31]}
   );
   gpc1_1 gpc490 (
      {stage0_20[55]},
      {stage1_20[32]}
   );
   gpc1_1 gpc491 (
      {stage0_20[56]},
      {stage1_20[33]}
   );
   gpc1_1 gpc492 (
      {stage0_20[57]},
      {stage1_20[34]}
   );
   gpc1_1 gpc493 (
      {stage0_20[58]},
      {stage1_20[35]}
   );
   gpc1_1 gpc494 (
      {stage0_20[59]},
      {stage1_20[36]}
   );
   gpc1_1 gpc495 (
      {stage0_20[60]},
      {stage1_20[37]}
   );
   gpc1_1 gpc496 (
      {stage0_20[61]},
      {stage1_20[38]}
   );
   gpc1_1 gpc497 (
      {stage0_20[62]},
      {stage1_20[39]}
   );
   gpc1_1 gpc498 (
      {stage0_20[63]},
      {stage1_20[40]}
   );
   gpc1_1 gpc499 (
      {stage0_21[55]},
      {stage1_21[24]}
   );
   gpc1_1 gpc500 (
      {stage0_21[56]},
      {stage1_21[25]}
   );
   gpc1_1 gpc501 (
      {stage0_21[57]},
      {stage1_21[26]}
   );
   gpc1_1 gpc502 (
      {stage0_21[58]},
      {stage1_21[27]}
   );
   gpc1_1 gpc503 (
      {stage0_21[59]},
      {stage1_21[28]}
   );
   gpc1_1 gpc504 (
      {stage0_21[60]},
      {stage1_21[29]}
   );
   gpc1_1 gpc505 (
      {stage0_21[61]},
      {stage1_21[30]}
   );
   gpc1_1 gpc506 (
      {stage0_21[62]},
      {stage1_21[31]}
   );
   gpc1_1 gpc507 (
      {stage0_21[63]},
      {stage1_21[32]}
   );
   gpc1_1 gpc508 (
      {stage0_22[52]},
      {stage1_22[19]}
   );
   gpc1_1 gpc509 (
      {stage0_22[53]},
      {stage1_22[20]}
   );
   gpc1_1 gpc510 (
      {stage0_22[54]},
      {stage1_22[21]}
   );
   gpc1_1 gpc511 (
      {stage0_22[55]},
      {stage1_22[22]}
   );
   gpc1_1 gpc512 (
      {stage0_22[56]},
      {stage1_22[23]}
   );
   gpc1_1 gpc513 (
      {stage0_22[57]},
      {stage1_22[24]}
   );
   gpc1_1 gpc514 (
      {stage0_22[58]},
      {stage1_22[25]}
   );
   gpc1_1 gpc515 (
      {stage0_22[59]},
      {stage1_22[26]}
   );
   gpc1_1 gpc516 (
      {stage0_22[60]},
      {stage1_22[27]}
   );
   gpc1_1 gpc517 (
      {stage0_22[61]},
      {stage1_22[28]}
   );
   gpc1_1 gpc518 (
      {stage0_22[62]},
      {stage1_22[29]}
   );
   gpc1_1 gpc519 (
      {stage0_22[63]},
      {stage1_22[30]}
   );
   gpc1_1 gpc520 (
      {stage0_23[48]},
      {stage1_23[19]}
   );
   gpc1_1 gpc521 (
      {stage0_23[49]},
      {stage1_23[20]}
   );
   gpc1_1 gpc522 (
      {stage0_23[50]},
      {stage1_23[21]}
   );
   gpc1_1 gpc523 (
      {stage0_23[51]},
      {stage1_23[22]}
   );
   gpc1_1 gpc524 (
      {stage0_23[52]},
      {stage1_23[23]}
   );
   gpc1_1 gpc525 (
      {stage0_23[53]},
      {stage1_23[24]}
   );
   gpc1_1 gpc526 (
      {stage0_23[54]},
      {stage1_23[25]}
   );
   gpc1_1 gpc527 (
      {stage0_23[55]},
      {stage1_23[26]}
   );
   gpc1_1 gpc528 (
      {stage0_23[56]},
      {stage1_23[27]}
   );
   gpc1_1 gpc529 (
      {stage0_23[57]},
      {stage1_23[28]}
   );
   gpc1_1 gpc530 (
      {stage0_23[58]},
      {stage1_23[29]}
   );
   gpc1_1 gpc531 (
      {stage0_23[59]},
      {stage1_23[30]}
   );
   gpc1_1 gpc532 (
      {stage0_23[60]},
      {stage1_23[31]}
   );
   gpc1_1 gpc533 (
      {stage0_23[61]},
      {stage1_23[32]}
   );
   gpc1_1 gpc534 (
      {stage0_23[62]},
      {stage1_23[33]}
   );
   gpc1_1 gpc535 (
      {stage0_23[63]},
      {stage1_23[34]}
   );
   gpc1_1 gpc536 (
      {stage0_24[62]},
      {stage1_24[25]}
   );
   gpc1_1 gpc537 (
      {stage0_24[63]},
      {stage1_24[26]}
   );
   gpc1_1 gpc538 (
      {stage0_25[42]},
      {stage1_25[23]}
   );
   gpc1_1 gpc539 (
      {stage0_25[43]},
      {stage1_25[24]}
   );
   gpc1_1 gpc540 (
      {stage0_25[44]},
      {stage1_25[25]}
   );
   gpc1_1 gpc541 (
      {stage0_25[45]},
      {stage1_25[26]}
   );
   gpc1_1 gpc542 (
      {stage0_25[46]},
      {stage1_25[27]}
   );
   gpc1_1 gpc543 (
      {stage0_25[47]},
      {stage1_25[28]}
   );
   gpc1_1 gpc544 (
      {stage0_25[48]},
      {stage1_25[29]}
   );
   gpc1_1 gpc545 (
      {stage0_25[49]},
      {stage1_25[30]}
   );
   gpc1_1 gpc546 (
      {stage0_25[50]},
      {stage1_25[31]}
   );
   gpc1_1 gpc547 (
      {stage0_25[51]},
      {stage1_25[32]}
   );
   gpc1_1 gpc548 (
      {stage0_25[52]},
      {stage1_25[33]}
   );
   gpc1_1 gpc549 (
      {stage0_25[53]},
      {stage1_25[34]}
   );
   gpc1_1 gpc550 (
      {stage0_25[54]},
      {stage1_25[35]}
   );
   gpc1_1 gpc551 (
      {stage0_25[55]},
      {stage1_25[36]}
   );
   gpc1_1 gpc552 (
      {stage0_25[56]},
      {stage1_25[37]}
   );
   gpc1_1 gpc553 (
      {stage0_25[57]},
      {stage1_25[38]}
   );
   gpc1_1 gpc554 (
      {stage0_25[58]},
      {stage1_25[39]}
   );
   gpc1_1 gpc555 (
      {stage0_25[59]},
      {stage1_25[40]}
   );
   gpc1_1 gpc556 (
      {stage0_25[60]},
      {stage1_25[41]}
   );
   gpc1_1 gpc557 (
      {stage0_25[61]},
      {stage1_25[42]}
   );
   gpc1_1 gpc558 (
      {stage0_25[62]},
      {stage1_25[43]}
   );
   gpc1_1 gpc559 (
      {stage0_25[63]},
      {stage1_25[44]}
   );
   gpc1_1 gpc560 (
      {stage0_26[53]},
      {stage1_26[18]}
   );
   gpc1_1 gpc561 (
      {stage0_26[54]},
      {stage1_26[19]}
   );
   gpc1_1 gpc562 (
      {stage0_26[55]},
      {stage1_26[20]}
   );
   gpc1_1 gpc563 (
      {stage0_26[56]},
      {stage1_26[21]}
   );
   gpc1_1 gpc564 (
      {stage0_26[57]},
      {stage1_26[22]}
   );
   gpc1_1 gpc565 (
      {stage0_26[58]},
      {stage1_26[23]}
   );
   gpc1_1 gpc566 (
      {stage0_26[59]},
      {stage1_26[24]}
   );
   gpc1_1 gpc567 (
      {stage0_26[60]},
      {stage1_26[25]}
   );
   gpc1_1 gpc568 (
      {stage0_26[61]},
      {stage1_26[26]}
   );
   gpc1_1 gpc569 (
      {stage0_26[62]},
      {stage1_26[27]}
   );
   gpc1_1 gpc570 (
      {stage0_26[63]},
      {stage1_26[28]}
   );
   gpc1_1 gpc571 (
      {stage0_27[41]},
      {stage1_27[18]}
   );
   gpc1_1 gpc572 (
      {stage0_27[42]},
      {stage1_27[19]}
   );
   gpc1_1 gpc573 (
      {stage0_27[43]},
      {stage1_27[20]}
   );
   gpc1_1 gpc574 (
      {stage0_27[44]},
      {stage1_27[21]}
   );
   gpc1_1 gpc575 (
      {stage0_27[45]},
      {stage1_27[22]}
   );
   gpc1_1 gpc576 (
      {stage0_27[46]},
      {stage1_27[23]}
   );
   gpc1_1 gpc577 (
      {stage0_27[47]},
      {stage1_27[24]}
   );
   gpc1_1 gpc578 (
      {stage0_27[48]},
      {stage1_27[25]}
   );
   gpc1_1 gpc579 (
      {stage0_27[49]},
      {stage1_27[26]}
   );
   gpc1_1 gpc580 (
      {stage0_27[50]},
      {stage1_27[27]}
   );
   gpc1_1 gpc581 (
      {stage0_27[51]},
      {stage1_27[28]}
   );
   gpc1_1 gpc582 (
      {stage0_27[52]},
      {stage1_27[29]}
   );
   gpc1_1 gpc583 (
      {stage0_27[53]},
      {stage1_27[30]}
   );
   gpc1_1 gpc584 (
      {stage0_27[54]},
      {stage1_27[31]}
   );
   gpc1_1 gpc585 (
      {stage0_27[55]},
      {stage1_27[32]}
   );
   gpc1_1 gpc586 (
      {stage0_27[56]},
      {stage1_27[33]}
   );
   gpc1_1 gpc587 (
      {stage0_27[57]},
      {stage1_27[34]}
   );
   gpc1_1 gpc588 (
      {stage0_27[58]},
      {stage1_27[35]}
   );
   gpc1_1 gpc589 (
      {stage0_27[59]},
      {stage1_27[36]}
   );
   gpc1_1 gpc590 (
      {stage0_27[60]},
      {stage1_27[37]}
   );
   gpc1_1 gpc591 (
      {stage0_27[61]},
      {stage1_27[38]}
   );
   gpc1_1 gpc592 (
      {stage0_27[62]},
      {stage1_27[39]}
   );
   gpc1_1 gpc593 (
      {stage0_27[63]},
      {stage1_27[40]}
   );
   gpc1_1 gpc594 (
      {stage0_28[62]},
      {stage1_28[25]}
   );
   gpc1_1 gpc595 (
      {stage0_28[63]},
      {stage1_28[26]}
   );
   gpc1_1 gpc596 (
      {stage0_29[60]},
      {stage1_29[25]}
   );
   gpc1_1 gpc597 (
      {stage0_29[61]},
      {stage1_29[26]}
   );
   gpc1_1 gpc598 (
      {stage0_29[62]},
      {stage1_29[27]}
   );
   gpc1_1 gpc599 (
      {stage0_29[63]},
      {stage1_29[28]}
   );
   gpc1_1 gpc600 (
      {stage0_30[59]},
      {stage1_30[21]}
   );
   gpc1_1 gpc601 (
      {stage0_30[60]},
      {stage1_30[22]}
   );
   gpc1_1 gpc602 (
      {stage0_30[61]},
      {stage1_30[23]}
   );
   gpc1_1 gpc603 (
      {stage0_30[62]},
      {stage1_30[24]}
   );
   gpc1_1 gpc604 (
      {stage0_30[63]},
      {stage1_30[25]}
   );
   gpc1_1 gpc605 (
      {stage0_32[63]},
      {stage1_32[30]}
   );
   gpc1_1 gpc606 (
      {stage0_33[53]},
      {stage1_33[27]}
   );
   gpc1_1 gpc607 (
      {stage0_33[54]},
      {stage1_33[28]}
   );
   gpc1_1 gpc608 (
      {stage0_33[55]},
      {stage1_33[29]}
   );
   gpc1_1 gpc609 (
      {stage0_33[56]},
      {stage1_33[30]}
   );
   gpc1_1 gpc610 (
      {stage0_33[57]},
      {stage1_33[31]}
   );
   gpc1_1 gpc611 (
      {stage0_33[58]},
      {stage1_33[32]}
   );
   gpc1_1 gpc612 (
      {stage0_33[59]},
      {stage1_33[33]}
   );
   gpc1_1 gpc613 (
      {stage0_33[60]},
      {stage1_33[34]}
   );
   gpc1_1 gpc614 (
      {stage0_33[61]},
      {stage1_33[35]}
   );
   gpc1_1 gpc615 (
      {stage0_33[62]},
      {stage1_33[36]}
   );
   gpc1_1 gpc616 (
      {stage0_33[63]},
      {stage1_33[37]}
   );
   gpc1_1 gpc617 (
      {stage0_34[60]},
      {stage1_34[20]}
   );
   gpc1_1 gpc618 (
      {stage0_34[61]},
      {stage1_34[21]}
   );
   gpc1_1 gpc619 (
      {stage0_34[62]},
      {stage1_34[22]}
   );
   gpc1_1 gpc620 (
      {stage0_34[63]},
      {stage1_34[23]}
   );
   gpc1_1 gpc621 (
      {stage0_35[57]},
      {stage1_35[23]}
   );
   gpc1_1 gpc622 (
      {stage0_35[58]},
      {stage1_35[24]}
   );
   gpc1_1 gpc623 (
      {stage0_35[59]},
      {stage1_35[25]}
   );
   gpc1_1 gpc624 (
      {stage0_35[60]},
      {stage1_35[26]}
   );
   gpc1_1 gpc625 (
      {stage0_35[61]},
      {stage1_35[27]}
   );
   gpc1_1 gpc626 (
      {stage0_35[62]},
      {stage1_35[28]}
   );
   gpc1_1 gpc627 (
      {stage0_35[63]},
      {stage1_35[29]}
   );
   gpc1_1 gpc628 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc629 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc630 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc631 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc632 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc633 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc634 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc635 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc636 (
      {stage0_36[54]},
      {stage1_36[34]}
   );
   gpc1_1 gpc637 (
      {stage0_36[55]},
      {stage1_36[35]}
   );
   gpc1_1 gpc638 (
      {stage0_36[56]},
      {stage1_36[36]}
   );
   gpc1_1 gpc639 (
      {stage0_36[57]},
      {stage1_36[37]}
   );
   gpc1_1 gpc640 (
      {stage0_36[58]},
      {stage1_36[38]}
   );
   gpc1_1 gpc641 (
      {stage0_36[59]},
      {stage1_36[39]}
   );
   gpc1_1 gpc642 (
      {stage0_36[60]},
      {stage1_36[40]}
   );
   gpc1_1 gpc643 (
      {stage0_36[61]},
      {stage1_36[41]}
   );
   gpc1_1 gpc644 (
      {stage0_36[62]},
      {stage1_36[42]}
   );
   gpc1_1 gpc645 (
      {stage0_36[63]},
      {stage1_36[43]}
   );
   gpc1_1 gpc646 (
      {stage0_38[41]},
      {stage1_38[19]}
   );
   gpc1_1 gpc647 (
      {stage0_38[42]},
      {stage1_38[20]}
   );
   gpc1_1 gpc648 (
      {stage0_38[43]},
      {stage1_38[21]}
   );
   gpc1_1 gpc649 (
      {stage0_38[44]},
      {stage1_38[22]}
   );
   gpc1_1 gpc650 (
      {stage0_38[45]},
      {stage1_38[23]}
   );
   gpc1_1 gpc651 (
      {stage0_38[46]},
      {stage1_38[24]}
   );
   gpc1_1 gpc652 (
      {stage0_38[47]},
      {stage1_38[25]}
   );
   gpc1_1 gpc653 (
      {stage0_38[48]},
      {stage1_38[26]}
   );
   gpc1_1 gpc654 (
      {stage0_38[49]},
      {stage1_38[27]}
   );
   gpc1_1 gpc655 (
      {stage0_38[50]},
      {stage1_38[28]}
   );
   gpc1_1 gpc656 (
      {stage0_38[51]},
      {stage1_38[29]}
   );
   gpc1_1 gpc657 (
      {stage0_38[52]},
      {stage1_38[30]}
   );
   gpc1_1 gpc658 (
      {stage0_38[53]},
      {stage1_38[31]}
   );
   gpc1_1 gpc659 (
      {stage0_38[54]},
      {stage1_38[32]}
   );
   gpc1_1 gpc660 (
      {stage0_38[55]},
      {stage1_38[33]}
   );
   gpc1_1 gpc661 (
      {stage0_38[56]},
      {stage1_38[34]}
   );
   gpc1_1 gpc662 (
      {stage0_38[57]},
      {stage1_38[35]}
   );
   gpc1_1 gpc663 (
      {stage0_38[58]},
      {stage1_38[36]}
   );
   gpc1_1 gpc664 (
      {stage0_38[59]},
      {stage1_38[37]}
   );
   gpc1_1 gpc665 (
      {stage0_38[60]},
      {stage1_38[38]}
   );
   gpc1_1 gpc666 (
      {stage0_38[61]},
      {stage1_38[39]}
   );
   gpc1_1 gpc667 (
      {stage0_38[62]},
      {stage1_38[40]}
   );
   gpc1_1 gpc668 (
      {stage0_38[63]},
      {stage1_38[41]}
   );
   gpc1_1 gpc669 (
      {stage0_39[63]},
      {stage1_39[22]}
   );
   gpc1_1 gpc670 (
      {stage0_41[54]},
      {stage1_41[26]}
   );
   gpc1_1 gpc671 (
      {stage0_41[55]},
      {stage1_41[27]}
   );
   gpc1_1 gpc672 (
      {stage0_41[56]},
      {stage1_41[28]}
   );
   gpc1_1 gpc673 (
      {stage0_41[57]},
      {stage1_41[29]}
   );
   gpc1_1 gpc674 (
      {stage0_41[58]},
      {stage1_41[30]}
   );
   gpc1_1 gpc675 (
      {stage0_41[59]},
      {stage1_41[31]}
   );
   gpc1_1 gpc676 (
      {stage0_41[60]},
      {stage1_41[32]}
   );
   gpc1_1 gpc677 (
      {stage0_41[61]},
      {stage1_41[33]}
   );
   gpc1_1 gpc678 (
      {stage0_41[62]},
      {stage1_41[34]}
   );
   gpc1_1 gpc679 (
      {stage0_41[63]},
      {stage1_41[35]}
   );
   gpc1_1 gpc680 (
      {stage0_42[54]},
      {stage1_42[19]}
   );
   gpc1_1 gpc681 (
      {stage0_42[55]},
      {stage1_42[20]}
   );
   gpc1_1 gpc682 (
      {stage0_42[56]},
      {stage1_42[21]}
   );
   gpc1_1 gpc683 (
      {stage0_42[57]},
      {stage1_42[22]}
   );
   gpc1_1 gpc684 (
      {stage0_42[58]},
      {stage1_42[23]}
   );
   gpc1_1 gpc685 (
      {stage0_42[59]},
      {stage1_42[24]}
   );
   gpc1_1 gpc686 (
      {stage0_42[60]},
      {stage1_42[25]}
   );
   gpc1_1 gpc687 (
      {stage0_42[61]},
      {stage1_42[26]}
   );
   gpc1_1 gpc688 (
      {stage0_42[62]},
      {stage1_42[27]}
   );
   gpc1_1 gpc689 (
      {stage0_42[63]},
      {stage1_42[28]}
   );
   gpc1_1 gpc690 (
      {stage0_43[50]},
      {stage1_43[22]}
   );
   gpc1_1 gpc691 (
      {stage0_43[51]},
      {stage1_43[23]}
   );
   gpc1_1 gpc692 (
      {stage0_43[52]},
      {stage1_43[24]}
   );
   gpc1_1 gpc693 (
      {stage0_43[53]},
      {stage1_43[25]}
   );
   gpc1_1 gpc694 (
      {stage0_43[54]},
      {stage1_43[26]}
   );
   gpc1_1 gpc695 (
      {stage0_43[55]},
      {stage1_43[27]}
   );
   gpc1_1 gpc696 (
      {stage0_43[56]},
      {stage1_43[28]}
   );
   gpc1_1 gpc697 (
      {stage0_43[57]},
      {stage1_43[29]}
   );
   gpc1_1 gpc698 (
      {stage0_43[58]},
      {stage1_43[30]}
   );
   gpc1_1 gpc699 (
      {stage0_43[59]},
      {stage1_43[31]}
   );
   gpc1_1 gpc700 (
      {stage0_43[60]},
      {stage1_43[32]}
   );
   gpc1_1 gpc701 (
      {stage0_43[61]},
      {stage1_43[33]}
   );
   gpc1_1 gpc702 (
      {stage0_43[62]},
      {stage1_43[34]}
   );
   gpc1_1 gpc703 (
      {stage0_43[63]},
      {stage1_43[35]}
   );
   gpc1_1 gpc704 (
      {stage0_44[58]},
      {stage1_44[27]}
   );
   gpc1_1 gpc705 (
      {stage0_44[59]},
      {stage1_44[28]}
   );
   gpc1_1 gpc706 (
      {stage0_44[60]},
      {stage1_44[29]}
   );
   gpc1_1 gpc707 (
      {stage0_44[61]},
      {stage1_44[30]}
   );
   gpc1_1 gpc708 (
      {stage0_44[62]},
      {stage1_44[31]}
   );
   gpc1_1 gpc709 (
      {stage0_44[63]},
      {stage1_44[32]}
   );
   gpc1_1 gpc710 (
      {stage0_45[36]},
      {stage1_45[20]}
   );
   gpc1_1 gpc711 (
      {stage0_45[37]},
      {stage1_45[21]}
   );
   gpc1_1 gpc712 (
      {stage0_45[38]},
      {stage1_45[22]}
   );
   gpc1_1 gpc713 (
      {stage0_45[39]},
      {stage1_45[23]}
   );
   gpc1_1 gpc714 (
      {stage0_45[40]},
      {stage1_45[24]}
   );
   gpc1_1 gpc715 (
      {stage0_45[41]},
      {stage1_45[25]}
   );
   gpc1_1 gpc716 (
      {stage0_45[42]},
      {stage1_45[26]}
   );
   gpc1_1 gpc717 (
      {stage0_45[43]},
      {stage1_45[27]}
   );
   gpc1_1 gpc718 (
      {stage0_45[44]},
      {stage1_45[28]}
   );
   gpc1_1 gpc719 (
      {stage0_45[45]},
      {stage1_45[29]}
   );
   gpc1_1 gpc720 (
      {stage0_45[46]},
      {stage1_45[30]}
   );
   gpc1_1 gpc721 (
      {stage0_45[47]},
      {stage1_45[31]}
   );
   gpc1_1 gpc722 (
      {stage0_45[48]},
      {stage1_45[32]}
   );
   gpc1_1 gpc723 (
      {stage0_45[49]},
      {stage1_45[33]}
   );
   gpc1_1 gpc724 (
      {stage0_45[50]},
      {stage1_45[34]}
   );
   gpc1_1 gpc725 (
      {stage0_45[51]},
      {stage1_45[35]}
   );
   gpc1_1 gpc726 (
      {stage0_45[52]},
      {stage1_45[36]}
   );
   gpc1_1 gpc727 (
      {stage0_45[53]},
      {stage1_45[37]}
   );
   gpc1_1 gpc728 (
      {stage0_45[54]},
      {stage1_45[38]}
   );
   gpc1_1 gpc729 (
      {stage0_45[55]},
      {stage1_45[39]}
   );
   gpc1_1 gpc730 (
      {stage0_45[56]},
      {stage1_45[40]}
   );
   gpc1_1 gpc731 (
      {stage0_45[57]},
      {stage1_45[41]}
   );
   gpc1_1 gpc732 (
      {stage0_45[58]},
      {stage1_45[42]}
   );
   gpc1_1 gpc733 (
      {stage0_45[59]},
      {stage1_45[43]}
   );
   gpc1_1 gpc734 (
      {stage0_45[60]},
      {stage1_45[44]}
   );
   gpc1_1 gpc735 (
      {stage0_45[61]},
      {stage1_45[45]}
   );
   gpc1_1 gpc736 (
      {stage0_45[62]},
      {stage1_45[46]}
   );
   gpc1_1 gpc737 (
      {stage0_45[63]},
      {stage1_45[47]}
   );
   gpc1_1 gpc738 (
      {stage0_47[46]},
      {stage1_47[23]}
   );
   gpc1_1 gpc739 (
      {stage0_47[47]},
      {stage1_47[24]}
   );
   gpc1_1 gpc740 (
      {stage0_47[48]},
      {stage1_47[25]}
   );
   gpc1_1 gpc741 (
      {stage0_47[49]},
      {stage1_47[26]}
   );
   gpc1_1 gpc742 (
      {stage0_47[50]},
      {stage1_47[27]}
   );
   gpc1_1 gpc743 (
      {stage0_47[51]},
      {stage1_47[28]}
   );
   gpc1_1 gpc744 (
      {stage0_47[52]},
      {stage1_47[29]}
   );
   gpc1_1 gpc745 (
      {stage0_47[53]},
      {stage1_47[30]}
   );
   gpc1_1 gpc746 (
      {stage0_47[54]},
      {stage1_47[31]}
   );
   gpc1_1 gpc747 (
      {stage0_47[55]},
      {stage1_47[32]}
   );
   gpc1_1 gpc748 (
      {stage0_47[56]},
      {stage1_47[33]}
   );
   gpc1_1 gpc749 (
      {stage0_47[57]},
      {stage1_47[34]}
   );
   gpc1_1 gpc750 (
      {stage0_47[58]},
      {stage1_47[35]}
   );
   gpc1_1 gpc751 (
      {stage0_47[59]},
      {stage1_47[36]}
   );
   gpc1_1 gpc752 (
      {stage0_47[60]},
      {stage1_47[37]}
   );
   gpc1_1 gpc753 (
      {stage0_47[61]},
      {stage1_47[38]}
   );
   gpc1_1 gpc754 (
      {stage0_47[62]},
      {stage1_47[39]}
   );
   gpc1_1 gpc755 (
      {stage0_47[63]},
      {stage1_47[40]}
   );
   gpc1_1 gpc756 (
      {stage0_48[58]},
      {stage1_48[26]}
   );
   gpc1_1 gpc757 (
      {stage0_48[59]},
      {stage1_48[27]}
   );
   gpc1_1 gpc758 (
      {stage0_48[60]},
      {stage1_48[28]}
   );
   gpc1_1 gpc759 (
      {stage0_48[61]},
      {stage1_48[29]}
   );
   gpc1_1 gpc760 (
      {stage0_48[62]},
      {stage1_48[30]}
   );
   gpc1_1 gpc761 (
      {stage0_48[63]},
      {stage1_48[31]}
   );
   gpc1_1 gpc762 (
      {stage0_49[60]},
      {stage1_49[21]}
   );
   gpc1_1 gpc763 (
      {stage0_49[61]},
      {stage1_49[22]}
   );
   gpc1_1 gpc764 (
      {stage0_49[62]},
      {stage1_49[23]}
   );
   gpc1_1 gpc765 (
      {stage0_49[63]},
      {stage1_49[24]}
   );
   gpc1_1 gpc766 (
      {stage0_50[62]},
      {stage1_50[23]}
   );
   gpc1_1 gpc767 (
      {stage0_50[63]},
      {stage1_50[24]}
   );
   gpc1_1 gpc768 (
      {stage0_51[59]},
      {stage1_51[27]}
   );
   gpc1_1 gpc769 (
      {stage0_51[60]},
      {stage1_51[28]}
   );
   gpc1_1 gpc770 (
      {stage0_51[61]},
      {stage1_51[29]}
   );
   gpc1_1 gpc771 (
      {stage0_51[62]},
      {stage1_51[30]}
   );
   gpc1_1 gpc772 (
      {stage0_51[63]},
      {stage1_51[31]}
   );
   gpc1_1 gpc773 (
      {stage0_52[45]},
      {stage1_52[24]}
   );
   gpc1_1 gpc774 (
      {stage0_52[46]},
      {stage1_52[25]}
   );
   gpc1_1 gpc775 (
      {stage0_52[47]},
      {stage1_52[26]}
   );
   gpc1_1 gpc776 (
      {stage0_52[48]},
      {stage1_52[27]}
   );
   gpc1_1 gpc777 (
      {stage0_52[49]},
      {stage1_52[28]}
   );
   gpc1_1 gpc778 (
      {stage0_52[50]},
      {stage1_52[29]}
   );
   gpc1_1 gpc779 (
      {stage0_52[51]},
      {stage1_52[30]}
   );
   gpc1_1 gpc780 (
      {stage0_52[52]},
      {stage1_52[31]}
   );
   gpc1_1 gpc781 (
      {stage0_52[53]},
      {stage1_52[32]}
   );
   gpc1_1 gpc782 (
      {stage0_52[54]},
      {stage1_52[33]}
   );
   gpc1_1 gpc783 (
      {stage0_52[55]},
      {stage1_52[34]}
   );
   gpc1_1 gpc784 (
      {stage0_52[56]},
      {stage1_52[35]}
   );
   gpc1_1 gpc785 (
      {stage0_52[57]},
      {stage1_52[36]}
   );
   gpc1_1 gpc786 (
      {stage0_52[58]},
      {stage1_52[37]}
   );
   gpc1_1 gpc787 (
      {stage0_52[59]},
      {stage1_52[38]}
   );
   gpc1_1 gpc788 (
      {stage0_52[60]},
      {stage1_52[39]}
   );
   gpc1_1 gpc789 (
      {stage0_52[61]},
      {stage1_52[40]}
   );
   gpc1_1 gpc790 (
      {stage0_52[62]},
      {stage1_52[41]}
   );
   gpc1_1 gpc791 (
      {stage0_52[63]},
      {stage1_52[42]}
   );
   gpc1_1 gpc792 (
      {stage0_53[58]},
      {stage1_53[21]}
   );
   gpc1_1 gpc793 (
      {stage0_53[59]},
      {stage1_53[22]}
   );
   gpc1_1 gpc794 (
      {stage0_53[60]},
      {stage1_53[23]}
   );
   gpc1_1 gpc795 (
      {stage0_53[61]},
      {stage1_53[24]}
   );
   gpc1_1 gpc796 (
      {stage0_53[62]},
      {stage1_53[25]}
   );
   gpc1_1 gpc797 (
      {stage0_53[63]},
      {stage1_53[26]}
   );
   gpc1_1 gpc798 (
      {stage0_54[54]},
      {stage1_54[23]}
   );
   gpc1_1 gpc799 (
      {stage0_54[55]},
      {stage1_54[24]}
   );
   gpc1_1 gpc800 (
      {stage0_54[56]},
      {stage1_54[25]}
   );
   gpc1_1 gpc801 (
      {stage0_54[57]},
      {stage1_54[26]}
   );
   gpc1_1 gpc802 (
      {stage0_54[58]},
      {stage1_54[27]}
   );
   gpc1_1 gpc803 (
      {stage0_54[59]},
      {stage1_54[28]}
   );
   gpc1_1 gpc804 (
      {stage0_54[60]},
      {stage1_54[29]}
   );
   gpc1_1 gpc805 (
      {stage0_54[61]},
      {stage1_54[30]}
   );
   gpc1_1 gpc806 (
      {stage0_54[62]},
      {stage1_54[31]}
   );
   gpc1_1 gpc807 (
      {stage0_54[63]},
      {stage1_54[32]}
   );
   gpc1_1 gpc808 (
      {stage0_56[62]},
      {stage1_56[24]}
   );
   gpc1_1 gpc809 (
      {stage0_56[63]},
      {stage1_56[25]}
   );
   gpc1_1 gpc810 (
      {stage0_58[47]},
      {stage1_58[24]}
   );
   gpc1_1 gpc811 (
      {stage0_58[48]},
      {stage1_58[25]}
   );
   gpc1_1 gpc812 (
      {stage0_58[49]},
      {stage1_58[26]}
   );
   gpc1_1 gpc813 (
      {stage0_58[50]},
      {stage1_58[27]}
   );
   gpc1_1 gpc814 (
      {stage0_58[51]},
      {stage1_58[28]}
   );
   gpc1_1 gpc815 (
      {stage0_58[52]},
      {stage1_58[29]}
   );
   gpc1_1 gpc816 (
      {stage0_58[53]},
      {stage1_58[30]}
   );
   gpc1_1 gpc817 (
      {stage0_58[54]},
      {stage1_58[31]}
   );
   gpc1_1 gpc818 (
      {stage0_58[55]},
      {stage1_58[32]}
   );
   gpc1_1 gpc819 (
      {stage0_58[56]},
      {stage1_58[33]}
   );
   gpc1_1 gpc820 (
      {stage0_58[57]},
      {stage1_58[34]}
   );
   gpc1_1 gpc821 (
      {stage0_58[58]},
      {stage1_58[35]}
   );
   gpc1_1 gpc822 (
      {stage0_58[59]},
      {stage1_58[36]}
   );
   gpc1_1 gpc823 (
      {stage0_58[60]},
      {stage1_58[37]}
   );
   gpc1_1 gpc824 (
      {stage0_58[61]},
      {stage1_58[38]}
   );
   gpc1_1 gpc825 (
      {stage0_58[62]},
      {stage1_58[39]}
   );
   gpc1_1 gpc826 (
      {stage0_58[63]},
      {stage1_58[40]}
   );
   gpc1_1 gpc827 (
      {stage0_59[42]},
      {stage1_59[20]}
   );
   gpc1_1 gpc828 (
      {stage0_59[43]},
      {stage1_59[21]}
   );
   gpc1_1 gpc829 (
      {stage0_59[44]},
      {stage1_59[22]}
   );
   gpc1_1 gpc830 (
      {stage0_59[45]},
      {stage1_59[23]}
   );
   gpc1_1 gpc831 (
      {stage0_59[46]},
      {stage1_59[24]}
   );
   gpc1_1 gpc832 (
      {stage0_59[47]},
      {stage1_59[25]}
   );
   gpc1_1 gpc833 (
      {stage0_59[48]},
      {stage1_59[26]}
   );
   gpc1_1 gpc834 (
      {stage0_59[49]},
      {stage1_59[27]}
   );
   gpc1_1 gpc835 (
      {stage0_59[50]},
      {stage1_59[28]}
   );
   gpc1_1 gpc836 (
      {stage0_59[51]},
      {stage1_59[29]}
   );
   gpc1_1 gpc837 (
      {stage0_59[52]},
      {stage1_59[30]}
   );
   gpc1_1 gpc838 (
      {stage0_59[53]},
      {stage1_59[31]}
   );
   gpc1_1 gpc839 (
      {stage0_59[54]},
      {stage1_59[32]}
   );
   gpc1_1 gpc840 (
      {stage0_59[55]},
      {stage1_59[33]}
   );
   gpc1_1 gpc841 (
      {stage0_59[56]},
      {stage1_59[34]}
   );
   gpc1_1 gpc842 (
      {stage0_59[57]},
      {stage1_59[35]}
   );
   gpc1_1 gpc843 (
      {stage0_59[58]},
      {stage1_59[36]}
   );
   gpc1_1 gpc844 (
      {stage0_59[59]},
      {stage1_59[37]}
   );
   gpc1_1 gpc845 (
      {stage0_59[60]},
      {stage1_59[38]}
   );
   gpc1_1 gpc846 (
      {stage0_59[61]},
      {stage1_59[39]}
   );
   gpc1_1 gpc847 (
      {stage0_59[62]},
      {stage1_59[40]}
   );
   gpc1_1 gpc848 (
      {stage0_59[63]},
      {stage1_59[41]}
   );
   gpc1_1 gpc849 (
      {stage0_60[52]},
      {stage1_60[21]}
   );
   gpc1_1 gpc850 (
      {stage0_60[53]},
      {stage1_60[22]}
   );
   gpc1_1 gpc851 (
      {stage0_60[54]},
      {stage1_60[23]}
   );
   gpc1_1 gpc852 (
      {stage0_60[55]},
      {stage1_60[24]}
   );
   gpc1_1 gpc853 (
      {stage0_60[56]},
      {stage1_60[25]}
   );
   gpc1_1 gpc854 (
      {stage0_60[57]},
      {stage1_60[26]}
   );
   gpc1_1 gpc855 (
      {stage0_60[58]},
      {stage1_60[27]}
   );
   gpc1_1 gpc856 (
      {stage0_60[59]},
      {stage1_60[28]}
   );
   gpc1_1 gpc857 (
      {stage0_60[60]},
      {stage1_60[29]}
   );
   gpc1_1 gpc858 (
      {stage0_60[61]},
      {stage1_60[30]}
   );
   gpc1_1 gpc859 (
      {stage0_60[62]},
      {stage1_60[31]}
   );
   gpc1_1 gpc860 (
      {stage0_60[63]},
      {stage1_60[32]}
   );
   gpc1_1 gpc861 (
      {stage0_61[58]},
      {stage1_61[25]}
   );
   gpc1_1 gpc862 (
      {stage0_61[59]},
      {stage1_61[26]}
   );
   gpc1_1 gpc863 (
      {stage0_61[60]},
      {stage1_61[27]}
   );
   gpc1_1 gpc864 (
      {stage0_61[61]},
      {stage1_61[28]}
   );
   gpc1_1 gpc865 (
      {stage0_61[62]},
      {stage1_61[29]}
   );
   gpc1_1 gpc866 (
      {stage0_61[63]},
      {stage1_61[30]}
   );
   gpc1_1 gpc867 (
      {stage0_62[51]},
      {stage1_62[20]}
   );
   gpc1_1 gpc868 (
      {stage0_62[52]},
      {stage1_62[21]}
   );
   gpc1_1 gpc869 (
      {stage0_62[53]},
      {stage1_62[22]}
   );
   gpc1_1 gpc870 (
      {stage0_62[54]},
      {stage1_62[23]}
   );
   gpc1_1 gpc871 (
      {stage0_62[55]},
      {stage1_62[24]}
   );
   gpc1_1 gpc872 (
      {stage0_62[56]},
      {stage1_62[25]}
   );
   gpc1_1 gpc873 (
      {stage0_62[57]},
      {stage1_62[26]}
   );
   gpc1_1 gpc874 (
      {stage0_62[58]},
      {stage1_62[27]}
   );
   gpc1_1 gpc875 (
      {stage0_62[59]},
      {stage1_62[28]}
   );
   gpc1_1 gpc876 (
      {stage0_62[60]},
      {stage1_62[29]}
   );
   gpc1_1 gpc877 (
      {stage0_62[61]},
      {stage1_62[30]}
   );
   gpc1_1 gpc878 (
      {stage0_62[62]},
      {stage1_62[31]}
   );
   gpc1_1 gpc879 (
      {stage0_62[63]},
      {stage1_62[32]}
   );
   gpc1_1 gpc880 (
      {stage0_63[54]},
      {stage1_63[18]}
   );
   gpc1_1 gpc881 (
      {stage0_63[55]},
      {stage1_63[19]}
   );
   gpc1_1 gpc882 (
      {stage0_63[56]},
      {stage1_63[20]}
   );
   gpc1_1 gpc883 (
      {stage0_63[57]},
      {stage1_63[21]}
   );
   gpc1_1 gpc884 (
      {stage0_63[58]},
      {stage1_63[22]}
   );
   gpc1_1 gpc885 (
      {stage0_63[59]},
      {stage1_63[23]}
   );
   gpc1_1 gpc886 (
      {stage0_63[60]},
      {stage1_63[24]}
   );
   gpc1_1 gpc887 (
      {stage0_63[61]},
      {stage1_63[25]}
   );
   gpc1_1 gpc888 (
      {stage0_63[62]},
      {stage1_63[26]}
   );
   gpc1_1 gpc889 (
      {stage0_63[63]},
      {stage1_63[27]}
   );
   gpc1163_5 gpc890 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc891 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc892 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc893 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc894 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc895 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], 1'b0, 1'b0},
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc896 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc897 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc898 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc899 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc900 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc901 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[12]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[11],stage2_3[11]}
   );
   gpc1163_5 gpc902 (
      {stage1_4[13], stage1_4[14], stage1_4[15]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[12]}
   );
   gpc606_5 gpc903 (
      {stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[13]}
   );
   gpc1325_5 gpc904 (
      {stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_5[12], stage1_5[13]},
      {stage1_6[7], stage1_6[8], stage1_6[9]},
      {stage1_7[1]},
      {stage2_8[2],stage2_7[3],stage2_6[5],stage2_5[8],stage2_4[14]}
   );
   gpc615_5 gpc905 (
      {stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13], stage1_6[14]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[3],stage2_7[4],stage2_6[6]}
   );
   gpc117_4 gpc906 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage1_8[6]},
      {stage1_9[0]},
      {stage2_10[1],stage2_9[1],stage2_8[4],stage2_7[5]}
   );
   gpc615_5 gpc907 (
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14]},
      {stage1_8[7]},
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[5],stage2_7[6]}
   );
   gpc615_5 gpc908 (
      {stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage1_8[8]},
      {stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11], stage1_9[12]},
      {stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[6],stage2_7[7]}
   );
   gpc615_5 gpc909 (
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage1_8[9]},
      {stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18]},
      {stage2_11[2],stage2_10[4],stage2_9[4],stage2_8[7],stage2_7[8]}
   );
   gpc606_5 gpc910 (
      {stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[3],stage2_10[5],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc911 (
      {stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc912 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[5],stage2_10[7]}
   );
   gpc615_5 gpc913 (
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[6]}
   );
   gpc615_5 gpc914 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4],stage2_11[7]}
   );
   gpc615_5 gpc915 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[4],stage2_12[5],stage2_11[8]}
   );
   gpc615_5 gpc916 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[5],stage2_12[6],stage2_11[9]}
   );
   gpc606_5 gpc917 (
      {stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[4],stage2_14[5],stage2_13[6],stage2_12[7]}
   );
   gpc615_5 gpc918 (
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28]},
      {stage1_14[6]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[5],stage2_14[6],stage2_13[7]}
   );
   gpc615_5 gpc919 (
      {stage1_13[29], stage1_13[30], 1'b0, 1'b0, 1'b0},
      {stage1_14[7]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[2],stage2_15[6],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc920 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[3],stage2_15[7],stage2_14[8]}
   );
   gpc615_5 gpc921 (
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[12]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[4],stage2_15[8],stage2_14[9]}
   );
   gpc615_5 gpc922 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[12]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[5],stage2_15[9]}
   );
   gpc615_5 gpc923 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22]},
      {stage1_16[13]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[6],stage2_15[10]}
   );
   gpc615_5 gpc924 (
      {stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage1_16[14]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[7],stage2_15[11]}
   );
   gpc615_5 gpc925 (
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32]},
      {stage1_16[15]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[8],stage2_15[12]}
   );
   gpc615_5 gpc926 (
      {stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[16]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[9],stage2_15[13]}
   );
   gpc615_5 gpc927 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21]},
      {stage1_17[30]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[10]}
   );
   gpc615_5 gpc928 (
      {stage1_16[22], stage1_16[23], stage1_16[24], stage1_16[25], stage1_16[26]},
      {stage1_17[31]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[11]}
   );
   gpc623_5 gpc929 (
      {stage1_17[32], stage1_17[33], stage1_17[34]},
      {stage1_18[12], stage1_18[13]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[7],stage2_18[9],stage2_17[11]}
   );
   gpc615_5 gpc930 (
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[8]}
   );
   gpc615_5 gpc931 (
      {stage1_19[11], stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[2],stage2_20[4],stage2_19[9]}
   );
   gpc615_5 gpc932 (
      {stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19], stage1_19[20]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[3],stage2_20[5],stage2_19[10]}
   );
   gpc615_5 gpc933 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[4],stage2_20[6],stage2_19[11]}
   );
   gpc606_5 gpc934 (
      {stage1_20[4], stage1_20[5], stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[4],stage2_22[4],stage2_21[5],stage2_20[7]}
   );
   gpc606_5 gpc935 (
      {stage1_20[10], stage1_20[11], stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[5],stage2_22[5],stage2_21[6],stage2_20[8]}
   );
   gpc606_5 gpc936 (
      {stage1_20[16], stage1_20[17], stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[6],stage2_22[6],stage2_21[7],stage2_20[9]}
   );
   gpc606_5 gpc937 (
      {stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[7],stage2_22[7],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc938 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[4],stage2_23[8],stage2_22[8],stage2_21[9]}
   );
   gpc1415_5 gpc939 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[6]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[1],stage2_24[5],stage2_23[9],stage2_22[9]}
   );
   gpc623_5 gpc940 (
      {stage1_22[29], stage1_22[30], 1'b0},
      {stage1_23[7], stage1_23[8]},
      {stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9]},
      {stage2_26[1],stage2_25[2],stage2_24[6],stage2_23[10],stage2_22[10]}
   );
   gpc615_5 gpc941 (
      {stage1_23[9], stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13]},
      {stage1_24[10]},
      {stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[7],stage2_23[11]}
   );
   gpc615_5 gpc942 (
      {stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17], stage1_23[18]},
      {stage1_24[11]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[8],stage2_23[12]}
   );
   gpc615_5 gpc943 (
      {stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage1_24[12]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[9],stage2_23[13]}
   );
   gpc615_5 gpc944 (
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28]},
      {stage1_24[13]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[3],stage2_26[5],stage2_25[6],stage2_24[10],stage2_23[14]}
   );
   gpc615_5 gpc945 (
      {stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33]},
      {stage1_24[14]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[4],stage2_26[6],stage2_25[7],stage2_24[11],stage2_23[15]}
   );
   gpc606_5 gpc946 (
      {stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19], stage1_24[20]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[7],stage2_25[8],stage2_24[12]}
   );
   gpc606_5 gpc947 (
      {stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25], stage1_24[26]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[8],stage2_25[9],stage2_24[13]}
   );
   gpc606_5 gpc948 (
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[9],stage2_25[10]}
   );
   gpc606_5 gpc949 (
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[10],stage2_25[11]}
   );
   gpc615_5 gpc950 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16]},
      {stage1_27[12]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[11]}
   );
   gpc615_5 gpc951 (
      {stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21]},
      {stage1_27[13]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[12]}
   );
   gpc615_5 gpc952 (
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18]},
      {stage1_28[12]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[2],stage2_29[4],stage2_28[6],stage2_27[11]}
   );
   gpc615_5 gpc953 (
      {stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage1_28[13]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[3],stage2_29[5],stage2_28[7],stage2_27[12]}
   );
   gpc615_5 gpc954 (
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28]},
      {stage1_28[14]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[4],stage2_29[6],stage2_28[8],stage2_27[13]}
   );
   gpc606_5 gpc955 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[3],stage2_30[5],stage2_29[7],stage2_28[9]}
   );
   gpc606_5 gpc956 (
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[4],stage2_30[6],stage2_29[8]}
   );
   gpc606_5 gpc957 (
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], 1'b0},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[5],stage2_30[7],stage2_29[9]}
   );
   gpc615_5 gpc958 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10]},
      {stage1_31[12]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[2],stage2_32[3],stage2_31[6],stage2_30[8]}
   );
   gpc615_5 gpc959 (
      {stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15]},
      {stage1_31[13]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[3],stage2_32[4],stage2_31[7],stage2_30[9]}
   );
   gpc615_5 gpc960 (
      {stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17], stage1_31[18]},
      {stage1_32[12]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[4],stage2_32[5],stage2_31[8]}
   );
   gpc606_5 gpc961 (
      {stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17], stage1_32[18]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[1],stage2_34[3],stage2_33[5],stage2_32[6]}
   );
   gpc606_5 gpc962 (
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[1],stage2_35[2],stage2_34[4],stage2_33[6]}
   );
   gpc606_5 gpc963 (
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[2],stage2_35[3],stage2_34[5],stage2_33[7]}
   );
   gpc606_5 gpc964 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[3],stage2_35[4],stage2_34[6],stage2_33[8]}
   );
   gpc615_5 gpc965 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[18]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[3],stage2_36[4],stage2_35[5],stage2_34[7]}
   );
   gpc615_5 gpc966 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[19]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[4],stage2_36[5],stage2_35[6],stage2_34[8]}
   );
   gpc615_5 gpc967 (
      {stage1_34[16], stage1_34[17], stage1_34[18], stage1_34[19], stage1_34[20]},
      {stage1_35[20]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[5],stage2_36[6],stage2_35[7],stage2_34[9]}
   );
   gpc615_5 gpc968 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[6],stage2_36[7],stage2_35[8]}
   );
   gpc606_5 gpc969 (
      {stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[1],stage2_38[4],stage2_37[7],stage2_36[8]}
   );
   gpc606_5 gpc970 (
      {stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30]},
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11]},
      {stage2_40[1],stage2_39[2],stage2_38[5],stage2_37[8],stage2_36[9]}
   );
   gpc606_5 gpc971 (
      {stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36]},
      {stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17]},
      {stage2_40[2],stage2_39[3],stage2_38[6],stage2_37[9],stage2_36[10]}
   );
   gpc606_5 gpc972 (
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[3],stage2_39[4],stage2_38[7],stage2_37[10]}
   );
   gpc606_5 gpc973 (
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[4],stage2_39[5],stage2_38[8],stage2_37[11]}
   );
   gpc1406_5 gpc974 (
      {stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3]},
      {stage1_41[0]},
      {stage2_42[0],stage2_41[2],stage2_40[5],stage2_39[6],stage2_38[9]}
   );
   gpc1325_5 gpc975 (
      {stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28]},
      {stage1_39[12], stage1_39[13]},
      {stage1_40[4], stage1_40[5], stage1_40[6]},
      {stage1_41[1]},
      {stage2_42[1],stage2_41[3],stage2_40[6],stage2_39[7],stage2_38[10]}
   );
   gpc615_5 gpc976 (
      {stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage1_40[7]},
      {stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5], stage1_41[6], stage1_41[7]},
      {stage2_43[0],stage2_42[2],stage2_41[4],stage2_40[7],stage2_39[8]}
   );
   gpc606_5 gpc977 (
      {stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11], stage1_40[12], stage1_40[13]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[1],stage2_42[3],stage2_41[5],stage2_40[8]}
   );
   gpc606_5 gpc978 (
      {stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17], stage1_40[18], stage1_40[19]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[2],stage2_42[4],stage2_41[6],stage2_40[9]}
   );
   gpc606_5 gpc979 (
      {stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23], stage1_40[24], stage1_40[25]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[3],stage2_42[5],stage2_41[7],stage2_40[10]}
   );
   gpc7_3 gpc980 (
      {stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11], stage1_41[12], stage1_41[13], stage1_41[14]},
      {stage2_43[4],stage2_42[6],stage2_41[8]}
   );
   gpc606_5 gpc981 (
      {stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19], stage1_41[20]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[3],stage2_43[5],stage2_42[7],stage2_41[9]}
   );
   gpc606_5 gpc982 (
      {stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24], stage1_41[25], stage1_41[26]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[4],stage2_43[6],stage2_42[8],stage2_41[10]}
   );
   gpc606_5 gpc983 (
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[2],stage2_44[5],stage2_43[7],stage2_42[9]}
   );
   gpc615_5 gpc984 (
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[3],stage2_44[6],stage2_43[8]}
   );
   gpc615_5 gpc985 (
      {stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[4],stage2_44[7],stage2_43[9]}
   );
   gpc615_5 gpc986 (
      {stage1_43[22], stage1_43[23], stage1_43[24], stage1_43[25], stage1_43[26]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[5],stage2_44[8],stage2_43[10]}
   );
   gpc615_5 gpc987 (
      {stage1_43[27], stage1_43[28], stage1_43[29], stage1_43[30], stage1_43[31]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[6],stage2_44[9],stage2_43[11]}
   );
   gpc615_5 gpc988 (
      {stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35], 1'b0},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[7],stage2_44[10],stage2_43[12]}
   );
   gpc606_5 gpc989 (
      {stage1_44[11], stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[5],stage2_46[6],stage2_45[8],stage2_44[11]}
   );
   gpc606_5 gpc990 (
      {stage1_44[17], stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[6],stage2_46[7],stage2_45[9],stage2_44[12]}
   );
   gpc606_5 gpc991 (
      {stage1_44[23], stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], 1'b0},
      {stage2_48[2],stage2_47[7],stage2_46[8],stage2_45[10],stage2_44[13]}
   );
   gpc606_5 gpc992 (
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[8],stage2_46[9],stage2_45[11]}
   );
   gpc606_5 gpc993 (
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[9],stage2_46[10],stage2_45[12]}
   );
   gpc606_5 gpc994 (
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[5],stage2_47[10],stage2_46[11],stage2_45[13]}
   );
   gpc606_5 gpc995 (
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[3],stage2_48[6],stage2_47[11]}
   );
   gpc606_5 gpc996 (
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[4],stage2_48[7],stage2_47[12]}
   );
   gpc606_5 gpc997 (
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[2],stage2_49[5],stage2_48[8],stage2_47[13]}
   );
   gpc117_4 gpc998 (
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6]},
      {stage1_49[18]},
      {stage1_50[0]},
      {stage2_51[3],stage2_50[3],stage2_49[6],stage2_48[9]}
   );
   gpc117_4 gpc999 (
      {stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_49[19]},
      {stage1_50[1]},
      {stage2_51[4],stage2_50[4],stage2_49[7],stage2_48[10]}
   );
   gpc117_4 gpc1000 (
      {stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17], stage1_48[18], stage1_48[19], stage1_48[20]},
      {stage1_49[20]},
      {stage1_50[2]},
      {stage2_51[5],stage2_50[5],stage2_49[8],stage2_48[11]}
   );
   gpc207_4 gpc1001 (
      {stage1_48[21], stage1_48[22], stage1_48[23], stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27]},
      {stage1_50[3], stage1_50[4]},
      {stage2_51[6],stage2_50[6],stage2_49[9],stage2_48[12]}
   );
   gpc606_5 gpc1002 (
      {stage1_49[21], stage1_49[22], stage1_49[23], stage1_49[24], 1'b0, 1'b0},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[0],stage2_51[7],stage2_50[7],stage2_49[10]}
   );
   gpc615_5 gpc1003 (
      {stage1_50[5], stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9]},
      {stage1_51[6]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[1],stage2_52[1],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc1004 (
      {stage1_50[10], stage1_50[11], stage1_50[12], stage1_50[13], stage1_50[14]},
      {stage1_51[7]},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage2_54[1],stage2_53[2],stage2_52[2],stage2_51[9],stage2_50[9]}
   );
   gpc615_5 gpc1005 (
      {stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18], stage1_50[19]},
      {stage1_51[8]},
      {stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17]},
      {stage2_54[2],stage2_53[3],stage2_52[3],stage2_51[10],stage2_50[10]}
   );
   gpc615_5 gpc1006 (
      {stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_51[9]},
      {stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23]},
      {stage2_54[3],stage2_53[4],stage2_52[4],stage2_51[11],stage2_50[11]}
   );
   gpc2116_5 gpc1007 (
      {stage1_51[10], stage1_51[11], stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15]},
      {stage1_52[24]},
      {stage1_53[0]},
      {stage1_54[0], stage1_54[1]},
      {stage2_55[0],stage2_54[4],stage2_53[5],stage2_52[5],stage2_51[12]}
   );
   gpc2116_5 gpc1008 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_52[25]},
      {stage1_53[1]},
      {stage1_54[2], stage1_54[3]},
      {stage2_55[1],stage2_54[5],stage2_53[6],stage2_52[6],stage2_51[13]}
   );
   gpc615_5 gpc1009 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26]},
      {stage1_52[26]},
      {stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5], stage1_53[6], stage1_53[7]},
      {stage2_55[2],stage2_54[6],stage2_53[7],stage2_52[7],stage2_51[14]}
   );
   gpc615_5 gpc1010 (
      {stage1_51[27], stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31]},
      {stage1_52[27]},
      {stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13]},
      {stage2_55[3],stage2_54[7],stage2_53[8],stage2_52[8],stage2_51[15]}
   );
   gpc615_5 gpc1011 (
      {stage1_52[28], stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32]},
      {stage1_53[14]},
      {stage1_54[4], stage1_54[5], stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9]},
      {stage2_56[0],stage2_55[4],stage2_54[8],stage2_53[9],stage2_52[9]}
   );
   gpc615_5 gpc1012 (
      {stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36], stage1_52[37]},
      {stage1_53[15]},
      {stage1_54[10], stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage2_56[1],stage2_55[5],stage2_54[9],stage2_53[10],stage2_52[10]}
   );
   gpc615_5 gpc1013 (
      {stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_53[16]},
      {stage1_54[16], stage1_54[17], stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21]},
      {stage2_56[2],stage2_55[6],stage2_54[10],stage2_53[11],stage2_52[11]}
   );
   gpc615_5 gpc1014 (
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage1_54[22]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[3],stage2_55[7],stage2_54[11],stage2_53[12]}
   );
   gpc1163_5 gpc1015 (
      {stage1_54[23], stage1_54[24], stage1_54[25]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage1_56[0]},
      {stage1_57[0]},
      {stage2_58[0],stage2_57[1],stage2_56[4],stage2_55[8],stage2_54[12]}
   );
   gpc1163_5 gpc1016 (
      {stage1_54[26], stage1_54[27], stage1_54[28]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[1]},
      {stage1_57[1]},
      {stage2_58[1],stage2_57[2],stage2_56[5],stage2_55[9],stage2_54[13]}
   );
   gpc615_5 gpc1017 (
      {stage1_54[29], stage1_54[30], stage1_54[31], stage1_54[32], 1'b0},
      {stage1_55[18]},
      {stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5], stage1_56[6], stage1_56[7]},
      {stage2_58[2],stage2_57[3],stage2_56[6],stage2_55[10],stage2_54[14]}
   );
   gpc606_5 gpc1018 (
      {stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11], stage1_56[12], stage1_56[13]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[0],stage2_58[3],stage2_57[4],stage2_56[7]}
   );
   gpc606_5 gpc1019 (
      {stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17], stage1_56[18], stage1_56[19]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[1],stage2_58[4],stage2_57[5],stage2_56[8]}
   );
   gpc606_5 gpc1020 (
      {stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[2],stage2_58[5],stage2_57[6],stage2_56[9]}
   );
   gpc606_5 gpc1021 (
      {stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5], stage1_57[6], stage1_57[7]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[3],stage2_59[3],stage2_58[6],stage2_57[7]}
   );
   gpc615_5 gpc1022 (
      {stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11], stage1_57[12]},
      {stage1_58[18]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[4],stage2_59[4],stage2_58[7],stage2_57[8]}
   );
   gpc615_5 gpc1023 (
      {stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage1_58[19]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[5],stage2_59[5],stage2_58[8],stage2_57[9]}
   );
   gpc615_5 gpc1024 (
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22]},
      {stage1_58[20]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[6],stage2_59[6],stage2_58[9],stage2_57[10]}
   );
   gpc615_5 gpc1025 (
      {stage1_58[21], stage1_58[22], stage1_58[23], stage1_58[24], stage1_58[25]},
      {stage1_59[24]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[4],stage2_60[7],stage2_59[7],stage2_58[10]}
   );
   gpc615_5 gpc1026 (
      {stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29], stage1_58[30]},
      {stage1_59[25]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[5],stage2_60[8],stage2_59[8],stage2_58[11]}
   );
   gpc615_5 gpc1027 (
      {stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage1_59[26]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[6],stage2_60[9],stage2_59[9],stage2_58[12]}
   );
   gpc606_5 gpc1028 (
      {stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30], stage1_59[31], stage1_59[32]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[3],stage2_61[7],stage2_60[10],stage2_59[10]}
   );
   gpc615_5 gpc1029 (
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22]},
      {stage1_61[6]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[1],stage2_62[4],stage2_61[8],stage2_60[11]}
   );
   gpc615_5 gpc1030 (
      {stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage1_61[7]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[2],stage2_62[5],stage2_61[9],stage2_60[12]}
   );
   gpc615_5 gpc1031 (
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32]},
      {stage1_61[8]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[3],stage2_62[6],stage2_61[10],stage2_60[13]}
   );
   gpc2135_5 gpc1032 (
      {stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12], stage1_61[13]},
      {stage1_62[18], stage1_62[19], stage1_62[20]},
      {stage1_63[0]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[0],stage2_64[3],stage2_63[4],stage2_62[7],stage2_61[11]}
   );
   gpc2135_5 gpc1033 (
      {stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage1_63[1]},
      {stage1_64[2], stage1_64[3]},
      {stage2_65[1],stage2_64[4],stage2_63[5],stage2_62[8],stage2_61[12]}
   );
   gpc606_5 gpc1034 (
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6], stage1_63[7]},
      {stage2_65[2],stage2_64[5],stage2_63[6],stage2_62[9],stage2_61[13]}
   );
   gpc606_5 gpc1035 (
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12], stage1_63[13]},
      {stage2_65[3],stage2_64[6],stage2_63[7],stage2_62[10],stage2_61[14]}
   );
   gpc606_5 gpc1036 (
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9]},
      {stage2_66[0],stage2_65[4],stage2_64[7],stage2_63[8],stage2_62[11]}
   );
   gpc615_5 gpc1037 (
      {stage1_62[30], stage1_62[31], stage1_62[32], 1'b0, 1'b0},
      {stage1_63[14]},
      {stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15]},
      {stage2_66[1],stage2_65[5],stage2_64[8],stage2_63[9],stage2_62[12]}
   );
   gpc606_5 gpc1038 (
      {stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_65[0], stage1_65[1], stage1_65[2], stage1_65[3], stage1_65[4], stage1_65[5]},
      {stage2_67[0],stage2_66[2],stage2_65[6],stage2_64[9],stage2_63[10]}
   );
   gpc606_5 gpc1039 (
      {stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_65[6], stage1_65[7], stage1_65[8], 1'b0, 1'b0, 1'b0},
      {stage2_67[1],stage2_66[3],stage2_65[7],stage2_64[10],stage2_63[11]}
   );
   gpc1_1 gpc1040 (
      {stage1_2[23]},
      {stage2_2[11]}
   );
   gpc1_1 gpc1041 (
      {stage1_4[27]},
      {stage2_4[15]}
   );
   gpc1_1 gpc1042 (
      {stage1_4[28]},
      {stage2_4[16]}
   );
   gpc1_1 gpc1043 (
      {stage1_4[29]},
      {stage2_4[17]}
   );
   gpc1_1 gpc1044 (
      {stage1_4[30]},
      {stage2_4[18]}
   );
   gpc1_1 gpc1045 (
      {stage1_4[31]},
      {stage2_4[19]}
   );
   gpc1_1 gpc1046 (
      {stage1_4[32]},
      {stage2_4[20]}
   );
   gpc1_1 gpc1047 (
      {stage1_4[33]},
      {stage2_4[21]}
   );
   gpc1_1 gpc1048 (
      {stage1_4[34]},
      {stage2_4[22]}
   );
   gpc1_1 gpc1049 (
      {stage1_4[35]},
      {stage2_4[23]}
   );
   gpc1_1 gpc1050 (
      {stage1_4[36]},
      {stage2_4[24]}
   );
   gpc1_1 gpc1051 (
      {stage1_4[37]},
      {stage2_4[25]}
   );
   gpc1_1 gpc1052 (
      {stage1_5[14]},
      {stage2_5[9]}
   );
   gpc1_1 gpc1053 (
      {stage1_5[15]},
      {stage2_5[10]}
   );
   gpc1_1 gpc1054 (
      {stage1_5[16]},
      {stage2_5[11]}
   );
   gpc1_1 gpc1055 (
      {stage1_5[17]},
      {stage2_5[12]}
   );
   gpc1_1 gpc1056 (
      {stage1_5[18]},
      {stage2_5[13]}
   );
   gpc1_1 gpc1057 (
      {stage1_5[19]},
      {stage2_5[14]}
   );
   gpc1_1 gpc1058 (
      {stage1_5[20]},
      {stage2_5[15]}
   );
   gpc1_1 gpc1059 (
      {stage1_5[21]},
      {stage2_5[16]}
   );
   gpc1_1 gpc1060 (
      {stage1_5[22]},
      {stage2_5[17]}
   );
   gpc1_1 gpc1061 (
      {stage1_5[23]},
      {stage2_5[18]}
   );
   gpc1_1 gpc1062 (
      {stage1_5[24]},
      {stage2_5[19]}
   );
   gpc1_1 gpc1063 (
      {stage1_5[25]},
      {stage2_5[20]}
   );
   gpc1_1 gpc1064 (
      {stage1_5[26]},
      {stage2_5[21]}
   );
   gpc1_1 gpc1065 (
      {stage1_6[15]},
      {stage2_6[7]}
   );
   gpc1_1 gpc1066 (
      {stage1_6[16]},
      {stage2_6[8]}
   );
   gpc1_1 gpc1067 (
      {stage1_6[17]},
      {stage2_6[9]}
   );
   gpc1_1 gpc1068 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc1069 (
      {stage1_6[19]},
      {stage2_6[11]}
   );
   gpc1_1 gpc1070 (
      {stage1_6[20]},
      {stage2_6[12]}
   );
   gpc1_1 gpc1071 (
      {stage1_6[21]},
      {stage2_6[13]}
   );
   gpc1_1 gpc1072 (
      {stage1_7[25]},
      {stage2_7[9]}
   );
   gpc1_1 gpc1073 (
      {stage1_7[26]},
      {stage2_7[10]}
   );
   gpc1_1 gpc1074 (
      {stage1_7[27]},
      {stage2_7[11]}
   );
   gpc1_1 gpc1075 (
      {stage1_7[28]},
      {stage2_7[12]}
   );
   gpc1_1 gpc1076 (
      {stage1_7[29]},
      {stage2_7[13]}
   );
   gpc1_1 gpc1077 (
      {stage1_7[30]},
      {stage2_7[14]}
   );
   gpc1_1 gpc1078 (
      {stage1_7[31]},
      {stage2_7[15]}
   );
   gpc1_1 gpc1079 (
      {stage1_7[32]},
      {stage2_7[16]}
   );
   gpc1_1 gpc1080 (
      {stage1_7[33]},
      {stage2_7[17]}
   );
   gpc1_1 gpc1081 (
      {stage1_7[34]},
      {stage2_7[18]}
   );
   gpc1_1 gpc1082 (
      {stage1_7[35]},
      {stage2_7[19]}
   );
   gpc1_1 gpc1083 (
      {stage1_8[16]},
      {stage2_8[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_8[17]},
      {stage2_8[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_8[18]},
      {stage2_8[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_8[19]},
      {stage2_8[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_8[20]},
      {stage2_8[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_8[21]},
      {stage2_8[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_8[22]},
      {stage2_8[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_8[23]},
      {stage2_8[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_8[24]},
      {stage2_8[17]}
   );
   gpc1_1 gpc1092 (
      {stage1_8[25]},
      {stage2_8[18]}
   );
   gpc1_1 gpc1093 (
      {stage1_8[26]},
      {stage2_8[19]}
   );
   gpc1_1 gpc1094 (
      {stage1_9[25]},
      {stage2_9[7]}
   );
   gpc1_1 gpc1095 (
      {stage1_9[26]},
      {stage2_9[8]}
   );
   gpc1_1 gpc1096 (
      {stage1_9[27]},
      {stage2_9[9]}
   );
   gpc1_1 gpc1097 (
      {stage1_9[28]},
      {stage2_9[10]}
   );
   gpc1_1 gpc1098 (
      {stage1_10[11]},
      {stage2_10[8]}
   );
   gpc1_1 gpc1099 (
      {stage1_10[12]},
      {stage2_10[9]}
   );
   gpc1_1 gpc1100 (
      {stage1_10[13]},
      {stage2_10[10]}
   );
   gpc1_1 gpc1101 (
      {stage1_10[14]},
      {stage2_10[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_10[15]},
      {stage2_10[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_10[16]},
      {stage2_10[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_10[17]},
      {stage2_10[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_10[18]},
      {stage2_10[15]}
   );
   gpc1_1 gpc1106 (
      {stage1_10[19]},
      {stage2_10[16]}
   );
   gpc1_1 gpc1107 (
      {stage1_10[20]},
      {stage2_10[17]}
   );
   gpc1_1 gpc1108 (
      {stage1_10[21]},
      {stage2_10[18]}
   );
   gpc1_1 gpc1109 (
      {stage1_10[22]},
      {stage2_10[19]}
   );
   gpc1_1 gpc1110 (
      {stage1_10[23]},
      {stage2_10[20]}
   );
   gpc1_1 gpc1111 (
      {stage1_10[24]},
      {stage2_10[21]}
   );
   gpc1_1 gpc1112 (
      {stage1_10[25]},
      {stage2_10[22]}
   );
   gpc1_1 gpc1113 (
      {stage1_10[26]},
      {stage2_10[23]}
   );
   gpc1_1 gpc1114 (
      {stage1_10[27]},
      {stage2_10[24]}
   );
   gpc1_1 gpc1115 (
      {stage1_10[28]},
      {stage2_10[25]}
   );
   gpc1_1 gpc1116 (
      {stage1_10[29]},
      {stage2_10[26]}
   );
   gpc1_1 gpc1117 (
      {stage1_10[30]},
      {stage2_10[27]}
   );
   gpc1_1 gpc1118 (
      {stage1_10[31]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1119 (
      {stage1_10[32]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1120 (
      {stage1_10[33]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1121 (
      {stage1_11[27]},
      {stage2_11[10]}
   );
   gpc1_1 gpc1122 (
      {stage1_11[28]},
      {stage2_11[11]}
   );
   gpc1_1 gpc1123 (
      {stage1_11[29]},
      {stage2_11[12]}
   );
   gpc1_1 gpc1124 (
      {stage1_11[30]},
      {stage2_11[13]}
   );
   gpc1_1 gpc1125 (
      {stage1_11[31]},
      {stage2_11[14]}
   );
   gpc1_1 gpc1126 (
      {stage1_11[32]},
      {stage2_11[15]}
   );
   gpc1_1 gpc1127 (
      {stage1_12[16]},
      {stage2_12[8]}
   );
   gpc1_1 gpc1128 (
      {stage1_12[17]},
      {stage2_12[9]}
   );
   gpc1_1 gpc1129 (
      {stage1_12[18]},
      {stage2_12[10]}
   );
   gpc1_1 gpc1130 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc1131 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc1132 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc1133 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc1134 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc1135 (
      {stage1_12[24]},
      {stage2_12[16]}
   );
   gpc1_1 gpc1136 (
      {stage1_12[25]},
      {stage2_12[17]}
   );
   gpc1_1 gpc1137 (
      {stage1_12[26]},
      {stage2_12[18]}
   );
   gpc1_1 gpc1138 (
      {stage1_14[19]},
      {stage2_14[10]}
   );
   gpc1_1 gpc1139 (
      {stage1_14[20]},
      {stage2_14[11]}
   );
   gpc1_1 gpc1140 (
      {stage1_14[21]},
      {stage2_14[12]}
   );
   gpc1_1 gpc1141 (
      {stage1_14[22]},
      {stage2_14[13]}
   );
   gpc1_1 gpc1142 (
      {stage1_14[23]},
      {stage2_14[14]}
   );
   gpc1_1 gpc1143 (
      {stage1_14[24]},
      {stage2_14[15]}
   );
   gpc1_1 gpc1144 (
      {stage1_15[38]},
      {stage2_15[14]}
   );
   gpc1_1 gpc1145 (
      {stage1_15[39]},
      {stage2_15[15]}
   );
   gpc1_1 gpc1146 (
      {stage1_15[40]},
      {stage2_15[16]}
   );
   gpc1_1 gpc1147 (
      {stage1_15[41]},
      {stage2_15[17]}
   );
   gpc1_1 gpc1148 (
      {stage1_15[42]},
      {stage2_15[18]}
   );
   gpc1_1 gpc1149 (
      {stage1_15[43]},
      {stage2_15[19]}
   );
   gpc1_1 gpc1150 (
      {stage1_15[44]},
      {stage2_15[20]}
   );
   gpc1_1 gpc1151 (
      {stage1_16[27]},
      {stage2_16[12]}
   );
   gpc1_1 gpc1152 (
      {stage1_16[28]},
      {stage2_16[13]}
   );
   gpc1_1 gpc1153 (
      {stage1_16[29]},
      {stage2_16[14]}
   );
   gpc1_1 gpc1154 (
      {stage1_16[30]},
      {stage2_16[15]}
   );
   gpc1_1 gpc1155 (
      {stage1_17[35]},
      {stage2_17[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_17[36]},
      {stage2_17[13]}
   );
   gpc1_1 gpc1157 (
      {stage1_17[37]},
      {stage2_17[14]}
   );
   gpc1_1 gpc1158 (
      {stage1_17[38]},
      {stage2_17[15]}
   );
   gpc1_1 gpc1159 (
      {stage1_17[39]},
      {stage2_17[16]}
   );
   gpc1_1 gpc1160 (
      {stage1_17[40]},
      {stage2_17[17]}
   );
   gpc1_1 gpc1161 (
      {stage1_17[41]},
      {stage2_17[18]}
   );
   gpc1_1 gpc1162 (
      {stage1_17[42]},
      {stage2_17[19]}
   );
   gpc1_1 gpc1163 (
      {stage1_17[43]},
      {stage2_17[20]}
   );
   gpc1_1 gpc1164 (
      {stage1_17[44]},
      {stage2_17[21]}
   );
   gpc1_1 gpc1165 (
      {stage1_18[14]},
      {stage2_18[10]}
   );
   gpc1_1 gpc1166 (
      {stage1_18[15]},
      {stage2_18[11]}
   );
   gpc1_1 gpc1167 (
      {stage1_18[16]},
      {stage2_18[12]}
   );
   gpc1_1 gpc1168 (
      {stage1_18[17]},
      {stage2_18[13]}
   );
   gpc1_1 gpc1169 (
      {stage1_18[18]},
      {stage2_18[14]}
   );
   gpc1_1 gpc1170 (
      {stage1_18[19]},
      {stage2_18[15]}
   );
   gpc1_1 gpc1171 (
      {stage1_18[20]},
      {stage2_18[16]}
   );
   gpc1_1 gpc1172 (
      {stage1_18[21]},
      {stage2_18[17]}
   );
   gpc1_1 gpc1173 (
      {stage1_18[22]},
      {stage2_18[18]}
   );
   gpc1_1 gpc1174 (
      {stage1_19[26]},
      {stage2_19[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_19[27]},
      {stage2_19[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_19[28]},
      {stage2_19[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_20[28]},
      {stage2_20[11]}
   );
   gpc1_1 gpc1178 (
      {stage1_20[29]},
      {stage2_20[12]}
   );
   gpc1_1 gpc1179 (
      {stage1_20[30]},
      {stage2_20[13]}
   );
   gpc1_1 gpc1180 (
      {stage1_20[31]},
      {stage2_20[14]}
   );
   gpc1_1 gpc1181 (
      {stage1_20[32]},
      {stage2_20[15]}
   );
   gpc1_1 gpc1182 (
      {stage1_20[33]},
      {stage2_20[16]}
   );
   gpc1_1 gpc1183 (
      {stage1_20[34]},
      {stage2_20[17]}
   );
   gpc1_1 gpc1184 (
      {stage1_20[35]},
      {stage2_20[18]}
   );
   gpc1_1 gpc1185 (
      {stage1_20[36]},
      {stage2_20[19]}
   );
   gpc1_1 gpc1186 (
      {stage1_20[37]},
      {stage2_20[20]}
   );
   gpc1_1 gpc1187 (
      {stage1_20[38]},
      {stage2_20[21]}
   );
   gpc1_1 gpc1188 (
      {stage1_20[39]},
      {stage2_20[22]}
   );
   gpc1_1 gpc1189 (
      {stage1_20[40]},
      {stage2_20[23]}
   );
   gpc1_1 gpc1190 (
      {stage1_21[30]},
      {stage2_21[10]}
   );
   gpc1_1 gpc1191 (
      {stage1_21[31]},
      {stage2_21[11]}
   );
   gpc1_1 gpc1192 (
      {stage1_21[32]},
      {stage2_21[12]}
   );
   gpc1_1 gpc1193 (
      {stage1_23[34]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1194 (
      {stage1_25[43]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1195 (
      {stage1_25[44]},
      {stage2_25[13]}
   );
   gpc1_1 gpc1196 (
      {stage1_26[22]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1197 (
      {stage1_26[23]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1198 (
      {stage1_26[24]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1199 (
      {stage1_26[25]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1200 (
      {stage1_26[26]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1201 (
      {stage1_26[27]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1202 (
      {stage1_26[28]},
      {stage2_26[19]}
   );
   gpc1_1 gpc1203 (
      {stage1_27[29]},
      {stage2_27[14]}
   );
   gpc1_1 gpc1204 (
      {stage1_27[30]},
      {stage2_27[15]}
   );
   gpc1_1 gpc1205 (
      {stage1_27[31]},
      {stage2_27[16]}
   );
   gpc1_1 gpc1206 (
      {stage1_27[32]},
      {stage2_27[17]}
   );
   gpc1_1 gpc1207 (
      {stage1_27[33]},
      {stage2_27[18]}
   );
   gpc1_1 gpc1208 (
      {stage1_27[34]},
      {stage2_27[19]}
   );
   gpc1_1 gpc1209 (
      {stage1_27[35]},
      {stage2_27[20]}
   );
   gpc1_1 gpc1210 (
      {stage1_27[36]},
      {stage2_27[21]}
   );
   gpc1_1 gpc1211 (
      {stage1_27[37]},
      {stage2_27[22]}
   );
   gpc1_1 gpc1212 (
      {stage1_27[38]},
      {stage2_27[23]}
   );
   gpc1_1 gpc1213 (
      {stage1_27[39]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1214 (
      {stage1_27[40]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1215 (
      {stage1_28[21]},
      {stage2_28[10]}
   );
   gpc1_1 gpc1216 (
      {stage1_28[22]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1217 (
      {stage1_28[23]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1218 (
      {stage1_28[24]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1219 (
      {stage1_28[25]},
      {stage2_28[14]}
   );
   gpc1_1 gpc1220 (
      {stage1_28[26]},
      {stage2_28[15]}
   );
   gpc1_1 gpc1221 (
      {stage1_30[16]},
      {stage2_30[10]}
   );
   gpc1_1 gpc1222 (
      {stage1_30[17]},
      {stage2_30[11]}
   );
   gpc1_1 gpc1223 (
      {stage1_30[18]},
      {stage2_30[12]}
   );
   gpc1_1 gpc1224 (
      {stage1_30[19]},
      {stage2_30[13]}
   );
   gpc1_1 gpc1225 (
      {stage1_30[20]},
      {stage2_30[14]}
   );
   gpc1_1 gpc1226 (
      {stage1_30[21]},
      {stage2_30[15]}
   );
   gpc1_1 gpc1227 (
      {stage1_30[22]},
      {stage2_30[16]}
   );
   gpc1_1 gpc1228 (
      {stage1_30[23]},
      {stage2_30[17]}
   );
   gpc1_1 gpc1229 (
      {stage1_30[24]},
      {stage2_30[18]}
   );
   gpc1_1 gpc1230 (
      {stage1_30[25]},
      {stage2_30[19]}
   );
   gpc1_1 gpc1231 (
      {stage1_31[19]},
      {stage2_31[9]}
   );
   gpc1_1 gpc1232 (
      {stage1_31[20]},
      {stage2_31[10]}
   );
   gpc1_1 gpc1233 (
      {stage1_31[21]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1234 (
      {stage1_31[22]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1235 (
      {stage1_32[19]},
      {stage2_32[7]}
   );
   gpc1_1 gpc1236 (
      {stage1_32[20]},
      {stage2_32[8]}
   );
   gpc1_1 gpc1237 (
      {stage1_32[21]},
      {stage2_32[9]}
   );
   gpc1_1 gpc1238 (
      {stage1_32[22]},
      {stage2_32[10]}
   );
   gpc1_1 gpc1239 (
      {stage1_32[23]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1240 (
      {stage1_32[24]},
      {stage2_32[12]}
   );
   gpc1_1 gpc1241 (
      {stage1_32[25]},
      {stage2_32[13]}
   );
   gpc1_1 gpc1242 (
      {stage1_32[26]},
      {stage2_32[14]}
   );
   gpc1_1 gpc1243 (
      {stage1_32[27]},
      {stage2_32[15]}
   );
   gpc1_1 gpc1244 (
      {stage1_32[28]},
      {stage2_32[16]}
   );
   gpc1_1 gpc1245 (
      {stage1_32[29]},
      {stage2_32[17]}
   );
   gpc1_1 gpc1246 (
      {stage1_32[30]},
      {stage2_32[18]}
   );
   gpc1_1 gpc1247 (
      {stage1_33[24]},
      {stage2_33[9]}
   );
   gpc1_1 gpc1248 (
      {stage1_33[25]},
      {stage2_33[10]}
   );
   gpc1_1 gpc1249 (
      {stage1_33[26]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1250 (
      {stage1_33[27]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1251 (
      {stage1_33[28]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1252 (
      {stage1_33[29]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1253 (
      {stage1_33[30]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1254 (
      {stage1_33[31]},
      {stage2_33[16]}
   );
   gpc1_1 gpc1255 (
      {stage1_33[32]},
      {stage2_33[17]}
   );
   gpc1_1 gpc1256 (
      {stage1_33[33]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1257 (
      {stage1_33[34]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1258 (
      {stage1_33[35]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1259 (
      {stage1_33[36]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1260 (
      {stage1_33[37]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1261 (
      {stage1_34[21]},
      {stage2_34[10]}
   );
   gpc1_1 gpc1262 (
      {stage1_34[22]},
      {stage2_34[11]}
   );
   gpc1_1 gpc1263 (
      {stage1_34[23]},
      {stage2_34[12]}
   );
   gpc1_1 gpc1264 (
      {stage1_35[26]},
      {stage2_35[9]}
   );
   gpc1_1 gpc1265 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1266 (
      {stage1_35[28]},
      {stage2_35[11]}
   );
   gpc1_1 gpc1267 (
      {stage1_35[29]},
      {stage2_35[12]}
   );
   gpc1_1 gpc1268 (
      {stage1_36[37]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1269 (
      {stage1_36[38]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1270 (
      {stage1_36[39]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1271 (
      {stage1_36[40]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1272 (
      {stage1_36[41]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1273 (
      {stage1_36[42]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1274 (
      {stage1_36[43]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1275 (
      {stage1_37[18]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1276 (
      {stage1_37[19]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1277 (
      {stage1_37[20]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1278 (
      {stage1_37[21]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1279 (
      {stage1_37[22]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1280 (
      {stage1_37[23]},
      {stage2_37[17]}
   );
   gpc1_1 gpc1281 (
      {stage1_38[29]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1282 (
      {stage1_38[30]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1283 (
      {stage1_38[31]},
      {stage2_38[13]}
   );
   gpc1_1 gpc1284 (
      {stage1_38[32]},
      {stage2_38[14]}
   );
   gpc1_1 gpc1285 (
      {stage1_38[33]},
      {stage2_38[15]}
   );
   gpc1_1 gpc1286 (
      {stage1_38[34]},
      {stage2_38[16]}
   );
   gpc1_1 gpc1287 (
      {stage1_38[35]},
      {stage2_38[17]}
   );
   gpc1_1 gpc1288 (
      {stage1_38[36]},
      {stage2_38[18]}
   );
   gpc1_1 gpc1289 (
      {stage1_38[37]},
      {stage2_38[19]}
   );
   gpc1_1 gpc1290 (
      {stage1_38[38]},
      {stage2_38[20]}
   );
   gpc1_1 gpc1291 (
      {stage1_38[39]},
      {stage2_38[21]}
   );
   gpc1_1 gpc1292 (
      {stage1_38[40]},
      {stage2_38[22]}
   );
   gpc1_1 gpc1293 (
      {stage1_38[41]},
      {stage2_38[23]}
   );
   gpc1_1 gpc1294 (
      {stage1_39[19]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1295 (
      {stage1_39[20]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1296 (
      {stage1_39[21]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1297 (
      {stage1_39[22]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1298 (
      {stage1_40[26]},
      {stage2_40[11]}
   );
   gpc1_1 gpc1299 (
      {stage1_41[27]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1300 (
      {stage1_41[28]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1301 (
      {stage1_41[29]},
      {stage2_41[13]}
   );
   gpc1_1 gpc1302 (
      {stage1_41[30]},
      {stage2_41[14]}
   );
   gpc1_1 gpc1303 (
      {stage1_41[31]},
      {stage2_41[15]}
   );
   gpc1_1 gpc1304 (
      {stage1_41[32]},
      {stage2_41[16]}
   );
   gpc1_1 gpc1305 (
      {stage1_41[33]},
      {stage2_41[17]}
   );
   gpc1_1 gpc1306 (
      {stage1_41[34]},
      {stage2_41[18]}
   );
   gpc1_1 gpc1307 (
      {stage1_41[35]},
      {stage2_41[19]}
   );
   gpc1_1 gpc1308 (
      {stage1_42[24]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1309 (
      {stage1_42[25]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1310 (
      {stage1_42[26]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1311 (
      {stage1_42[27]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1312 (
      {stage1_42[28]},
      {stage2_42[14]}
   );
   gpc1_1 gpc1313 (
      {stage1_44[29]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1314 (
      {stage1_44[30]},
      {stage2_44[15]}
   );
   gpc1_1 gpc1315 (
      {stage1_44[31]},
      {stage2_44[16]}
   );
   gpc1_1 gpc1316 (
      {stage1_44[32]},
      {stage2_44[17]}
   );
   gpc1_1 gpc1317 (
      {stage1_47[36]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1318 (
      {stage1_47[37]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1319 (
      {stage1_47[38]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1320 (
      {stage1_47[39]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1321 (
      {stage1_47[40]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1322 (
      {stage1_48[28]},
      {stage2_48[13]}
   );
   gpc1_1 gpc1323 (
      {stage1_48[29]},
      {stage2_48[14]}
   );
   gpc1_1 gpc1324 (
      {stage1_48[30]},
      {stage2_48[15]}
   );
   gpc1_1 gpc1325 (
      {stage1_48[31]},
      {stage2_48[16]}
   );
   gpc1_1 gpc1326 (
      {stage1_53[22]},
      {stage2_53[13]}
   );
   gpc1_1 gpc1327 (
      {stage1_53[23]},
      {stage2_53[14]}
   );
   gpc1_1 gpc1328 (
      {stage1_53[24]},
      {stage2_53[15]}
   );
   gpc1_1 gpc1329 (
      {stage1_53[25]},
      {stage2_53[16]}
   );
   gpc1_1 gpc1330 (
      {stage1_53[26]},
      {stage2_53[17]}
   );
   gpc1_1 gpc1331 (
      {stage1_55[19]},
      {stage2_55[11]}
   );
   gpc1_1 gpc1332 (
      {stage1_55[20]},
      {stage2_55[12]}
   );
   gpc1_1 gpc1333 (
      {stage1_55[21]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1334 (
      {stage1_55[22]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1335 (
      {stage1_55[23]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1336 (
      {stage1_55[24]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1337 (
      {stage1_57[23]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1338 (
      {stage1_57[24]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1339 (
      {stage1_57[25]},
      {stage2_57[13]}
   );
   gpc1_1 gpc1340 (
      {stage1_58[36]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1341 (
      {stage1_58[37]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1342 (
      {stage1_58[38]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1343 (
      {stage1_58[39]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1344 (
      {stage1_58[40]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1345 (
      {stage1_59[33]},
      {stage2_59[11]}
   );
   gpc1_1 gpc1346 (
      {stage1_59[34]},
      {stage2_59[12]}
   );
   gpc1_1 gpc1347 (
      {stage1_59[35]},
      {stage2_59[13]}
   );
   gpc1_1 gpc1348 (
      {stage1_59[36]},
      {stage2_59[14]}
   );
   gpc1_1 gpc1349 (
      {stage1_59[37]},
      {stage2_59[15]}
   );
   gpc1_1 gpc1350 (
      {stage1_59[38]},
      {stage2_59[16]}
   );
   gpc1_1 gpc1351 (
      {stage1_59[39]},
      {stage2_59[17]}
   );
   gpc1_1 gpc1352 (
      {stage1_59[40]},
      {stage2_59[18]}
   );
   gpc1_1 gpc1353 (
      {stage1_59[41]},
      {stage2_59[19]}
   );
   gpc1_1 gpc1354 (
      {stage1_63[27]},
      {stage2_63[12]}
   );
   gpc606_5 gpc1355 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc1356 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc1357 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1358 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc606_5 gpc1359 (
      {stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4]}
   );
   gpc606_5 gpc1360 (
      {stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5]}
   );
   gpc606_5 gpc1361 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc606_5 gpc1362 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc1325_5 gpc1363 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], 1'b0},
      {stage2_6[12], stage2_6[13]},
      {stage2_7[12], stage2_7[13], stage2_7[14]},
      {stage2_8[0]},
      {stage3_9[2],stage3_8[4],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc606_5 gpc1364 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc1365 (
      {stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc1366 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[7]}
   );
   gpc606_5 gpc1367 (
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[3],stage3_10[3],stage3_9[6]}
   );
   gpc1163_5 gpc1368 (
      {stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[1],stage3_12[4],stage3_11[4],stage3_10[4]}
   );
   gpc615_5 gpc1369 (
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25]},
      {stage2_11[12]},
      {stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6]},
      {stage3_14[1],stage3_13[2],stage3_12[5],stage3_11[5],stage3_10[5]}
   );
   gpc615_5 gpc1370 (
      {stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_11[13]},
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage3_14[2],stage3_13[3],stage3_12[6],stage3_11[6],stage3_10[6]}
   );
   gpc606_5 gpc1371 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[7]}
   );
   gpc615_5 gpc1372 (
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_14[6]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[1],stage3_14[4],stage3_13[5]}
   );
   gpc615_5 gpc1373 (
      {stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[2],stage3_15[2],stage3_14[5]}
   );
   gpc615_5 gpc1374 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], 1'b0},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[3],stage3_15[3],stage3_14[6]}
   );
   gpc615_5 gpc1375 (
      {stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12]},
      {stage2_16[12]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[3],stage3_16[4],stage3_15[4]}
   );
   gpc615_5 gpc1376 (
      {stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage2_16[13]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[3],stage3_17[4],stage3_16[5],stage3_15[5]}
   );
   gpc606_5 gpc1377 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[2],stage3_18[4],stage3_17[5]}
   );
   gpc606_5 gpc1378 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], 1'b0, 1'b0},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[3],stage3_18[5],stage3_17[6]}
   );
   gpc615_5 gpc1379 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[2],stage3_20[2],stage3_19[4],stage3_18[6]}
   );
   gpc615_5 gpc1380 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[13]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[3],stage3_20[3],stage3_19[5],stage3_18[7]}
   );
   gpc615_5 gpc1381 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[14]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[4],stage3_20[4],stage3_19[6],stage3_18[8]}
   );
   gpc606_5 gpc1382 (
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[3],stage3_21[5],stage3_20[5]}
   );
   gpc606_5 gpc1383 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[1],stage3_22[4],stage3_21[6]}
   );
   gpc606_5 gpc1384 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[2],stage3_22[5],stage3_21[7]}
   );
   gpc615_5 gpc1385 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[3],stage3_23[3],stage3_22[6]}
   );
   gpc606_5 gpc1386 (
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[3],stage3_24[4]}
   );
   gpc606_5 gpc1387 (
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[4]}
   );
   gpc606_5 gpc1388 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[5]}
   );
   gpc135_4 gpc1389 (
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10]},
      {stage2_27[12], stage2_27[13], stage2_27[14]},
      {stage2_28[0]},
      {stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc135_4 gpc1390 (
      {stage2_26[11], stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15]},
      {stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage2_28[1]},
      {stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc135_4 gpc1391 (
      {stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20]},
      {stage2_28[2]},
      {stage3_29[4],stage3_28[5],stage3_27[5],stage3_26[6]}
   );
   gpc615_5 gpc1392 (
      {stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25]},
      {stage2_28[3]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[5],stage3_28[6],stage3_27[6]}
   );
   gpc606_5 gpc1393 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[1],stage3_29[6],stage3_28[7]}
   );
   gpc606_5 gpc1394 (
      {stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[2],stage3_29[7],stage3_28[8]}
   );
   gpc606_5 gpc1395 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], 1'b0, 1'b0},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[2],stage3_31[3],stage3_30[3],stage3_29[8]}
   );
   gpc615_5 gpc1396 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[3],stage3_31[4],stage3_30[4]}
   );
   gpc615_5 gpc1397 (
      {stage2_30[17], stage2_30[18], stage2_30[19], 1'b0, 1'b0},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[4],stage3_31[5],stage3_30[5]}
   );
   gpc615_5 gpc1398 (
      {stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12]},
      {stage2_32[12]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[2],stage3_33[3],stage3_32[5],stage3_31[6]}
   );
   gpc606_5 gpc1399 (
      {stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[1],stage3_34[3],stage3_33[4],stage3_32[6]}
   );
   gpc606_5 gpc1400 (
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[2],stage3_34[4],stage3_33[5]}
   );
   gpc615_5 gpc1401 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10]},
      {stage2_35[6]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[2],stage3_35[3],stage3_34[5]}
   );
   gpc615_5 gpc1402 (
      {stage2_34[11], stage2_34[12], 1'b0, 1'b0, 1'b0},
      {stage2_35[7]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[3],stage3_35[4],stage3_34[6]}
   );
   gpc615_5 gpc1403 (
      {stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[4],stage3_35[5]}
   );
   gpc606_5 gpc1404 (
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4]}
   );
   gpc606_5 gpc1405 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc207_4 gpc1406 (
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6]},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[2],stage3_39[3],stage3_38[5]}
   );
   gpc207_4 gpc1407 (
      {stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage2_40[2], stage2_40[3]},
      {stage3_41[3],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc207_4 gpc1408 (
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_40[4], stage2_40[5]},
      {stage3_41[4],stage3_40[4],stage3_39[5],stage3_38[7]}
   );
   gpc606_5 gpc1409 (
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[0],stage3_42[0],stage3_41[5],stage3_40[5]}
   );
   gpc135_4 gpc1410 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4]},
      {stage2_42[6], stage2_42[7], stage2_42[8]},
      {stage2_43[0]},
      {stage3_44[1],stage3_43[1],stage3_42[1],stage3_41[6]}
   );
   gpc135_4 gpc1411 (
      {stage2_41[5], stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9]},
      {stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage2_43[1]},
      {stage3_44[2],stage3_43[2],stage3_42[2],stage3_41[7]}
   );
   gpc135_4 gpc1412 (
      {stage2_41[10], stage2_41[11], stage2_41[12], stage2_41[13], stage2_41[14]},
      {stage2_42[12], stage2_42[13], stage2_42[14]},
      {stage2_43[2]},
      {stage3_44[3],stage3_43[3],stage3_42[3],stage3_41[8]}
   );
   gpc615_5 gpc1413 (
      {stage2_43[3], stage2_43[4], stage2_43[5], stage2_43[6], stage2_43[7]},
      {stage2_44[0]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[4]}
   );
   gpc615_5 gpc1414 (
      {stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11], stage2_43[12]},
      {stage2_44[1]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[5]}
   );
   gpc606_5 gpc1415 (
      {stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5], stage2_44[6], stage2_44[7]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[2],stage3_46[2],stage3_45[2],stage3_44[6]}
   );
   gpc1163_5 gpc1416 (
      {stage2_46[6], stage2_46[7], stage2_46[8]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[0],stage3_48[1],stage3_47[3],stage3_46[3]}
   );
   gpc1325_5 gpc1417 (
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10]},
      {stage2_48[1], stage2_48[2]},
      {stage2_49[1], stage2_49[2], stage2_49[3]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[1],stage3_49[1],stage3_48[2],stage3_47[4]}
   );
   gpc1325_5 gpc1418 (
      {stage2_47[11], stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15]},
      {stage2_48[3], stage2_48[4]},
      {stage2_49[4], stage2_49[5], stage2_49[6]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[2],stage3_49[2],stage3_48[3],stage3_47[5]}
   );
   gpc1406_5 gpc1419 (
      {stage2_48[5], stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[2],stage3_50[3],stage3_49[3],stage3_48[4]}
   );
   gpc1406_5 gpc1420 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9]},
      {stage2_51[1]},
      {stage3_52[1],stage3_51[3],stage3_50[4],stage3_49[4],stage3_48[5]}
   );
   gpc615_5 gpc1421 (
      {stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], 1'b0},
      {stage2_50[10]},
      {stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7]},
      {stage3_53[0],stage3_52[2],stage3_51[4],stage3_50[5],stage3_49[5]}
   );
   gpc615_5 gpc1422 (
      {stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[1],stage3_52[3],stage3_51[5]}
   );
   gpc615_5 gpc1423 (
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage2_53[6]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[1],stage3_54[1],stage3_53[2],stage3_52[4]}
   );
   gpc615_5 gpc1424 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10]},
      {stage2_53[7]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[2],stage3_54[2],stage3_53[3],stage3_52[5]}
   );
   gpc615_5 gpc1425 (
      {stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11], stage2_53[12]},
      {stage2_54[12]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[2],stage3_55[3],stage3_54[3],stage3_53[4]}
   );
   gpc615_5 gpc1426 (
      {stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage2_54[13]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[3],stage3_55[4],stage3_54[4],stage3_53[5]}
   );
   gpc615_5 gpc1427 (
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[2],stage3_56[4]}
   );
   gpc615_5 gpc1428 (
      {stage2_56[5], stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[3],stage3_56[5]}
   );
   gpc615_5 gpc1429 (
      {stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6]},
      {stage2_58[12]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[4]}
   );
   gpc615_5 gpc1430 (
      {stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage2_58[13]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[5]}
   );
   gpc615_5 gpc1431 (
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16]},
      {stage2_60[0]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[0],stage3_61[2],stage3_60[4],stage3_59[4]}
   );
   gpc615_5 gpc1432 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_61[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[1],stage3_62[1],stage3_61[3],stage3_60[5]}
   );
   gpc606_5 gpc1433 (
      {stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[1],stage3_63[2],stage3_62[2],stage3_61[4]}
   );
   gpc606_5 gpc1434 (
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[2],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1435 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[3],stage3_63[4]}
   );
   gpc1406_5 gpc1436 (
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], 1'b0},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3]},
      {stage2_67[0]},
      {stage3_68[0],stage3_67[1],stage3_66[2],stage3_65[3],stage3_64[4]}
   );
   gpc1_1 gpc1437 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc1438 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1439 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1440 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1441 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1442 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1443 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc1444 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1445 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1446 (
      {stage2_3[11]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1447 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1448 (
      {stage2_7[15]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1449 (
      {stage2_7[16]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1450 (
      {stage2_7[17]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1451 (
      {stage2_7[18]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1452 (
      {stage2_7[19]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1453 (
      {stage2_8[19]},
      {stage3_8[8]}
   );
   gpc1_1 gpc1454 (
      {stage2_9[6]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1455 (
      {stage2_9[7]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1456 (
      {stage2_9[8]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1457 (
      {stage2_9[9]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1458 (
      {stage2_9[10]},
      {stage3_9[11]}
   );
   gpc1_1 gpc1459 (
      {stage2_11[14]},
      {stage3_11[7]}
   );
   gpc1_1 gpc1460 (
      {stage2_11[15]},
      {stage3_11[8]}
   );
   gpc1_1 gpc1461 (
      {stage2_13[6]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1462 (
      {stage2_13[7]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1463 (
      {stage2_13[8]},
      {stage3_13[8]}
   );
   gpc1_1 gpc1464 (
      {stage2_15[18]},
      {stage3_15[6]}
   );
   gpc1_1 gpc1465 (
      {stage2_15[19]},
      {stage3_15[7]}
   );
   gpc1_1 gpc1466 (
      {stage2_15[20]},
      {stage3_15[8]}
   );
   gpc1_1 gpc1467 (
      {stage2_16[14]},
      {stage3_16[6]}
   );
   gpc1_1 gpc1468 (
      {stage2_16[15]},
      {stage3_16[7]}
   );
   gpc1_1 gpc1469 (
      {stage2_18[15]},
      {stage3_18[9]}
   );
   gpc1_1 gpc1470 (
      {stage2_18[16]},
      {stage3_18[10]}
   );
   gpc1_1 gpc1471 (
      {stage2_18[17]},
      {stage3_18[11]}
   );
   gpc1_1 gpc1472 (
      {stage2_18[18]},
      {stage3_18[12]}
   );
   gpc1_1 gpc1473 (
      {stage2_21[12]},
      {stage3_21[8]}
   );
   gpc1_1 gpc1474 (
      {stage2_23[13]},
      {stage3_23[4]}
   );
   gpc1_1 gpc1475 (
      {stage2_23[14]},
      {stage3_23[5]}
   );
   gpc1_1 gpc1476 (
      {stage2_23[15]},
      {stage3_23[6]}
   );
   gpc1_1 gpc1477 (
      {stage2_23[16]},
      {stage3_23[7]}
   );
   gpc1_1 gpc1478 (
      {stage2_24[12]},
      {stage3_24[5]}
   );
   gpc1_1 gpc1479 (
      {stage2_24[13]},
      {stage3_24[6]}
   );
   gpc1_1 gpc1480 (
      {stage2_25[12]},
      {stage3_25[6]}
   );
   gpc1_1 gpc1481 (
      {stage2_25[13]},
      {stage3_25[7]}
   );
   gpc1_1 gpc1482 (
      {stage2_33[12]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1483 (
      {stage2_33[13]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1484 (
      {stage2_33[14]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1485 (
      {stage2_33[15]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1486 (
      {stage2_33[16]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1487 (
      {stage2_33[17]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1488 (
      {stage2_33[18]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1489 (
      {stage2_33[19]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1490 (
      {stage2_33[20]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1491 (
      {stage2_33[21]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1492 (
      {stage2_33[22]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1493 (
      {stage2_36[13]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1494 (
      {stage2_36[14]},
      {stage3_36[6]}
   );
   gpc1_1 gpc1495 (
      {stage2_36[15]},
      {stage3_36[7]}
   );
   gpc1_1 gpc1496 (
      {stage2_36[16]},
      {stage3_36[8]}
   );
   gpc1_1 gpc1497 (
      {stage2_36[17]},
      {stage3_36[9]}
   );
   gpc1_1 gpc1498 (
      {stage2_38[21]},
      {stage3_38[8]}
   );
   gpc1_1 gpc1499 (
      {stage2_38[22]},
      {stage3_38[9]}
   );
   gpc1_1 gpc1500 (
      {stage2_38[23]},
      {stage3_38[10]}
   );
   gpc1_1 gpc1501 (
      {stage2_39[12]},
      {stage3_39[6]}
   );
   gpc1_1 gpc1502 (
      {stage2_41[15]},
      {stage3_41[9]}
   );
   gpc1_1 gpc1503 (
      {stage2_41[16]},
      {stage3_41[10]}
   );
   gpc1_1 gpc1504 (
      {stage2_41[17]},
      {stage3_41[11]}
   );
   gpc1_1 gpc1505 (
      {stage2_41[18]},
      {stage3_41[12]}
   );
   gpc1_1 gpc1506 (
      {stage2_41[19]},
      {stage3_41[13]}
   );
   gpc1_1 gpc1507 (
      {stage2_44[8]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1508 (
      {stage2_44[9]},
      {stage3_44[8]}
   );
   gpc1_1 gpc1509 (
      {stage2_44[10]},
      {stage3_44[9]}
   );
   gpc1_1 gpc1510 (
      {stage2_44[11]},
      {stage3_44[10]}
   );
   gpc1_1 gpc1511 (
      {stage2_44[12]},
      {stage3_44[11]}
   );
   gpc1_1 gpc1512 (
      {stage2_44[13]},
      {stage3_44[12]}
   );
   gpc1_1 gpc1513 (
      {stage2_44[14]},
      {stage3_44[13]}
   );
   gpc1_1 gpc1514 (
      {stage2_44[15]},
      {stage3_44[14]}
   );
   gpc1_1 gpc1515 (
      {stage2_44[16]},
      {stage3_44[15]}
   );
   gpc1_1 gpc1516 (
      {stage2_44[17]},
      {stage3_44[16]}
   );
   gpc1_1 gpc1517 (
      {stage2_45[12]},
      {stage3_45[3]}
   );
   gpc1_1 gpc1518 (
      {stage2_45[13]},
      {stage3_45[4]}
   );
   gpc1_1 gpc1519 (
      {stage2_46[9]},
      {stage3_46[4]}
   );
   gpc1_1 gpc1520 (
      {stage2_46[10]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1521 (
      {stage2_46[11]},
      {stage3_46[6]}
   );
   gpc1_1 gpc1522 (
      {stage2_47[16]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1523 (
      {stage2_47[17]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1524 (
      {stage2_47[18]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1525 (
      {stage2_50[11]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1526 (
      {stage2_51[13]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1527 (
      {stage2_51[14]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1528 (
      {stage2_51[15]},
      {stage3_51[8]}
   );
   gpc1_1 gpc1529 (
      {stage2_52[11]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1530 (
      {stage2_54[14]},
      {stage3_54[5]}
   );
   gpc1_1 gpc1531 (
      {stage2_55[12]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1532 (
      {stage2_55[13]},
      {stage3_55[6]}
   );
   gpc1_1 gpc1533 (
      {stage2_55[14]},
      {stage3_55[7]}
   );
   gpc1_1 gpc1534 (
      {stage2_55[15]},
      {stage3_55[8]}
   );
   gpc1_1 gpc1535 (
      {stage2_55[16]},
      {stage3_55[9]}
   );
   gpc1_1 gpc1536 (
      {stage2_57[12]},
      {stage3_57[6]}
   );
   gpc1_1 gpc1537 (
      {stage2_57[13]},
      {stage3_57[7]}
   );
   gpc1_1 gpc1538 (
      {stage2_58[14]},
      {stage3_58[4]}
   );
   gpc1_1 gpc1539 (
      {stage2_58[15]},
      {stage3_58[5]}
   );
   gpc1_1 gpc1540 (
      {stage2_58[16]},
      {stage3_58[6]}
   );
   gpc1_1 gpc1541 (
      {stage2_58[17]},
      {stage3_58[7]}
   );
   gpc1_1 gpc1542 (
      {stage2_59[17]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1543 (
      {stage2_59[18]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1544 (
      {stage2_59[19]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1545 (
      {stage2_60[6]},
      {stage3_60[6]}
   );
   gpc1_1 gpc1546 (
      {stage2_60[7]},
      {stage3_60[7]}
   );
   gpc1_1 gpc1547 (
      {stage2_60[8]},
      {stage3_60[8]}
   );
   gpc1_1 gpc1548 (
      {stage2_60[9]},
      {stage3_60[9]}
   );
   gpc1_1 gpc1549 (
      {stage2_60[10]},
      {stage3_60[10]}
   );
   gpc1_1 gpc1550 (
      {stage2_60[11]},
      {stage3_60[11]}
   );
   gpc1_1 gpc1551 (
      {stage2_60[12]},
      {stage3_60[12]}
   );
   gpc1_1 gpc1552 (
      {stage2_60[13]},
      {stage3_60[13]}
   );
   gpc1_1 gpc1553 (
      {stage2_61[13]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1554 (
      {stage2_61[14]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1555 (
      {stage2_62[12]},
      {stage3_62[4]}
   );
   gpc1_1 gpc1556 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1557 (
      {stage2_65[6]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1558 (
      {stage2_65[7]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1559 (
      {stage2_67[1]},
      {stage3_67[2]}
   );
   gpc135_4 gpc1560 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[0]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1325_5 gpc1561 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[1]}
   );
   gpc1163_5 gpc1562 (
      {stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[1]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc1563 (
      {stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc1564 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1565 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc207_4 gpc1566 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1567 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4]},
      {stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3]}
   );
   gpc135_4 gpc1568 (
      {stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], 1'b0},
      {stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[1]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4]}
   );
   gpc117_4 gpc1569 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc7_3 gpc1570 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], 1'b0},
      {stage4_16[1],stage4_15[1],stage4_14[3]}
   );
   gpc117_4 gpc1571 (
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7]},
      {stage3_16[0]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[2],stage4_15[2]}
   );
   gpc606_5 gpc1572 (
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1],stage4_16[3]}
   );
   gpc606_5 gpc1573 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[2]}
   );
   gpc117_4 gpc1574 (
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage3_19[6]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[2],stage4_19[2],stage4_18[3]}
   );
   gpc606_5 gpc1575 (
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5], 1'b0},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[3]}
   );
   gpc215_4 gpc1576 (
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4]},
      {stage3_22[6]},
      {stage3_23[0], stage3_23[1]},
      {stage4_24[1],stage4_23[1],stage4_22[1],stage4_21[3]}
   );
   gpc615_5 gpc1577 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[2]}
   );
   gpc606_5 gpc1578 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[1],stage4_26[1],stage4_25[1],stage4_24[3]}
   );
   gpc606_5 gpc1579 (
      {stage3_25[6], stage3_25[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[1],stage4_27[2],stage4_26[2],stage4_25[2]}
   );
   gpc2135_5 gpc1580 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[2]}
   );
   gpc2135_5 gpc1581 (
      {stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8], 1'b0},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[2],stage4_28[3]}
   );
   gpc1343_5 gpc1582 (
      {stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc7_3 gpc1583 (
      {stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5], stage3_32[6], 1'b0},
      {stage4_34[0],stage4_33[1],stage4_32[3]}
   );
   gpc2135_5 gpc1584 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[2]}
   );
   gpc2135_5 gpc1585 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[3]}
   );
   gpc606_5 gpc1586 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15]},
      {stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5], 1'b0, 1'b0},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1587 (
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3],stage4_36[3]}
   );
   gpc606_5 gpc1588 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[1],stage4_39[1],stage4_38[1],stage4_37[4]}
   );
   gpc615_5 gpc1589 (
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10]},
      {stage3_39[6]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[1],stage4_40[2],stage4_39[2],stage4_38[2]}
   );
   gpc207_4 gpc1590 (
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[1],stage4_41[2]}
   );
   gpc207_4 gpc1591 (
      {stage3_41[7], stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[2],stage4_41[3]}
   );
   gpc615_5 gpc1592 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], 1'b0},
      {stage3_43[4]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[3]}
   );
   gpc2135_5 gpc1593 (
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10]},
      {stage3_45[0], stage3_45[1], stage3_45[2]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc2135_5 gpc1594 (
      {stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage3_45[3], stage3_45[4], 1'b0},
      {stage3_46[1]},
      {stage3_47[2], stage3_47[3]},
      {stage4_48[1],stage4_47[1],stage4_46[2],stage4_45[2],stage4_44[4]}
   );
   gpc615_5 gpc1595 (
      {stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_47[4]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[2],stage4_47[2],stage4_46[3]}
   );
   gpc1406_5 gpc1596 (
      {stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8], 1'b0, 1'b0},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3]},
      {stage3_50[0]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[3],stage4_47[3]}
   );
   gpc615_5 gpc1597 (
      {stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[0],stage4_51[1],stage4_50[2]}
   );
   gpc615_5 gpc1598 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage3_52[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[1],stage4_51[2]}
   );
   gpc606_5 gpc1599 (
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[0],stage4_55[1],stage4_54[2]}
   );
   gpc606_5 gpc1600 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[1],stage4_55[2]}
   );
   gpc615_5 gpc1601 (
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4]},
      {stage3_59[0]},
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage4_62[0],stage4_61[0],stage4_60[0],stage4_59[1],stage4_58[2]}
   );
   gpc7_3 gpc1602 (
      {stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7]},
      {stage4_61[1],stage4_60[1],stage4_59[2]}
   );
   gpc615_5 gpc1603 (
      {stage3_60[6], stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10]},
      {stage3_61[0]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], 1'b0},
      {stage4_64[0],stage4_63[0],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc615_5 gpc1604 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {1'b0},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[1],stage4_63[1],stage4_62[2],stage4_61[3]}
   );
   gpc1325_5 gpc1605 (
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4]},
      {stage3_66[0], stage3_66[1]},
      {stage3_67[0], stage3_67[1], stage3_67[2]},
      {stage3_68[0]},
      {stage4_69[0],stage4_68[0],stage4_67[0],stage4_66[0],stage4_65[1]}
   );
   gpc1_1 gpc1606 (
      {stage3_0[5]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1607 (
      {stage3_1[3]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1608 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc1609 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1610 (
      {stage3_4[5]},
      {stage4_4[2]}
   );
   gpc1_1 gpc1611 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1612 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc1613 (
      {stage3_15[8]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1614 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc1615 (
      {stage3_21[5]},
      {stage4_21[4]}
   );
   gpc1_1 gpc1616 (
      {stage3_21[6]},
      {stage4_21[5]}
   );
   gpc1_1 gpc1617 (
      {stage3_21[7]},
      {stage4_21[6]}
   );
   gpc1_1 gpc1618 (
      {stage3_21[8]},
      {stage4_21[7]}
   );
   gpc1_1 gpc1619 (
      {stage3_23[7]},
      {stage4_23[3]}
   );
   gpc1_1 gpc1620 (
      {stage3_26[6]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1621 (
      {stage3_27[6]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1622 (
      {stage3_33[16]},
      {stage4_33[5]}
   );
   gpc1_1 gpc1623 (
      {stage3_34[6]},
      {stage4_34[4]}
   );
   gpc1_1 gpc1624 (
      {stage3_43[5]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1625 (
      {stage3_44[16]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1626 (
      {stage3_49[4]},
      {stage4_49[2]}
   );
   gpc1_1 gpc1627 (
      {stage3_49[5]},
      {stage4_49[3]}
   );
   gpc1_1 gpc1628 (
      {stage3_50[6]},
      {stage4_50[3]}
   );
   gpc1_1 gpc1629 (
      {stage3_51[6]},
      {stage4_51[3]}
   );
   gpc1_1 gpc1630 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1631 (
      {stage3_51[8]},
      {stage4_51[5]}
   );
   gpc1_1 gpc1632 (
      {stage3_55[6]},
      {stage4_55[3]}
   );
   gpc1_1 gpc1633 (
      {stage3_55[7]},
      {stage4_55[4]}
   );
   gpc1_1 gpc1634 (
      {stage3_55[8]},
      {stage4_55[5]}
   );
   gpc1_1 gpc1635 (
      {stage3_55[9]},
      {stage4_55[6]}
   );
   gpc1_1 gpc1636 (
      {stage3_57[6]},
      {stage4_57[2]}
   );
   gpc1_1 gpc1637 (
      {stage3_57[7]},
      {stage4_57[3]}
   );
   gpc1_1 gpc1638 (
      {stage3_58[5]},
      {stage4_58[3]}
   );
   gpc1_1 gpc1639 (
      {stage3_58[6]},
      {stage4_58[4]}
   );
   gpc1_1 gpc1640 (
      {stage3_58[7]},
      {stage4_58[5]}
   );
   gpc1_1 gpc1641 (
      {stage3_60[11]},
      {stage4_60[3]}
   );
   gpc1_1 gpc1642 (
      {stage3_60[12]},
      {stage4_60[4]}
   );
   gpc1_1 gpc1643 (
      {stage3_60[13]},
      {stage4_60[5]}
   );
   gpc1_1 gpc1644 (
      {stage3_61[6]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1645 (
      {stage3_64[0]},
      {stage4_64[2]}
   );
   gpc1_1 gpc1646 (
      {stage3_64[1]},
      {stage4_64[3]}
   );
   gpc1_1 gpc1647 (
      {stage3_64[2]},
      {stage4_64[4]}
   );
   gpc1_1 gpc1648 (
      {stage3_64[3]},
      {stage4_64[5]}
   );
   gpc1_1 gpc1649 (
      {stage3_64[4]},
      {stage4_64[6]}
   );
   gpc1_1 gpc1650 (
      {stage3_65[5]},
      {stage4_65[2]}
   );
   gpc1_1 gpc1651 (
      {stage3_66[2]},
      {stage4_66[1]}
   );
   gpc1343_5 gpc1652 (
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0], stage4_3[1], 1'b0, 1'b0},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc623_5 gpc1653 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], 1'b0},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1]}
   );
   gpc3_2 gpc1654 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage5_8[1],stage5_7[1]}
   );
   gpc1343_5 gpc1655 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1423_5 gpc1656 (
      {stage4_11[3], stage4_11[4], 1'b0},
      {stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1343_5 gpc1657 (
      {stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc1658 (
      {stage4_16[3], stage4_16[4], 1'b0},
      {stage4_17[1], stage4_17[2]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc1659 (
      {stage4_19[1], stage4_19[2], 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc615_5 gpc1660 (
      {stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6], stage4_21[7]},
      {stage4_22[1]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], 1'b0, 1'b0},
      {stage5_25[0],stage5_24[0],stage5_23[1],stage5_22[1],stage5_21[1]}
   );
   gpc135_4 gpc1661 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc1343_5 gpc1662 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1], stage4_28[2]},
      {stage4_29[0]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[1],stage5_26[1]}
   );
   gpc135_4 gpc1663 (
      {stage4_29[1], stage4_29[2], stage4_29[3], 1'b0, 1'b0},
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[1]}
   );
   gpc1343_5 gpc1664 (
      {stage4_31[1], stage4_31[2], 1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0], stage4_33[1], stage4_33[2]},
      {stage4_34[0]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[1],stage5_31[1]}
   );
   gpc1343_5 gpc1665 (
      {stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[1],stage5_33[1]}
   );
   gpc1163_5 gpc1666 (
      {stage4_36[1], stage4_36[2], stage4_36[3]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], 1'b0},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc1423_5 gpc1667 (
      {stage4_38[1], stage4_38[2], 1'b0},
      {stage4_39[1], stage4_39[2]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1668 (
      {stage4_41[1], stage4_41[2], stage4_41[3]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3]},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1669 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1670 (
      {stage4_46[1], stage4_46[2], stage4_46[3]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1163_5 gpc1671 (
      {stage4_49[1], stage4_49[2], stage4_49[3]},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], 1'b0, 1'b0},
      {stage4_51[0]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc215_4 gpc1672 (
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5]},
      {stage4_52[1]},
      {stage4_53[0], stage4_53[1]},
      {stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc3_2 gpc1673 (
      {stage4_54[0], stage4_54[1], stage4_54[2]},
      {stage5_55[0],stage5_54[1]}
   );
   gpc7_3 gpc1674 (
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5], stage4_55[6]},
      {stage5_57[0],stage5_56[0],stage5_55[1]}
   );
   gpc1343_5 gpc1675 (
      {stage4_56[0], stage4_56[1], 1'b0},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3]},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[0],stage5_57[1],stage5_56[1]}
   );
   gpc623_5 gpc1676 (
      {stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage4_59[1], stage4_59[2]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[1]}
   );
   gpc2135_5 gpc1677 (
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc2135_5 gpc1678 (
      {stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2]},
      {stage4_66[0]},
      {stage4_67[0], 1'b0},
      {stage5_68[0],stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1]}
   );
   gpc1_1 gpc1679 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1680 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1681 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1682 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1683 (
      {stage4_4[3]},
      {stage5_4[1]}
   );
   gpc1_1 gpc1684 (
      {stage4_5[1]},
      {stage5_5[1]}
   );
   gpc1_1 gpc1685 (
      {stage4_28[3]},
      {stage5_28[1]}
   );
   gpc1_1 gpc1686 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1687 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
   gpc1_1 gpc1688 (
      {stage4_63[1]},
      {stage5_63[1]}
   );
   gpc1_1 gpc1689 (
      {stage4_66[1]},
      {stage5_66[1]}
   );
   gpc1_1 gpc1690 (
      {stage4_68[0]},
      {stage5_68[1]}
   );
   gpc1_1 gpc1691 (
      {stage4_69[0]},
      {stage5_69[0]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor_CLA64_64 compressor_CLA64_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h670398822a5899e84c65922986b2a185f5980f7702bb1d5764e304318a62de5bafb4817b6d67b4cbe6598cbc969bd923a088d93bc9cb8f9eb7e37850fd107a1aff592da8af21dd1c3a21fd8ca34b0af453ceec5424315beb02cf3703e54aa8e719c4d5766ec87f5b5b9a617ee299fca40bf3cb11cc9b63b2fb3c294c126c2f661f6b7ef93346b037e12398aa57ff13b85338718c09e90614c491c77eac2926b674f469dd3f5106d1a342451efce31939d4eca2e8dcc21f373c91ef72ecbce25876a8133824b68976b96b2ce576600ec7be24553fd2f00cdbd756e3098f61eaf61198c56ee2201a9cda15b06f6df7f04abf427cbf85628a6ea432a6280c72fa5efe5465536b6e4cfc576e7373136a2d95106f3b872b0608c156c2fd108d4d0ca8e959a5f021a5da1adca8632e00ac3cea306a22a69b8193b4548839b2858590e954438b73277afac7c0ec77e382bb4bfbc5e429df018f161978d533747c8efa639dcc6608c828b657aa03eac8c9470483d097b2fb6c8be7912ba0232ad5caaf652b1f5b16af9ec53123d82438bc74e5e3e9e523df713039bf7ce8e6a53c40a592587741558c03a4b74eb08297791195ca06e7a6ff016e25fb9b005a0ac21d805c936010364dcf8d0c5891d7b45f33ae86d105868496544c2db3d089b66ab0fa899a32218b6759f19c52371bacaa89cda7893efabb50673a1e43748453269f2f8b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3fbd74838079c745e9ff6a5acae7576f7d84b97c2ea444ba57cd4ec7e2b961aa01f28c9822689e0ccab1d62d157ee6d75caab222a509ac6c51ffe93741f10fb1d8e55bba2b2f014f1898284516470c4b78206f6c2d609cbdce094699fa5b489aee24bea2dd00eeda9ad7b0f50f33957cd46d436733d65da5c300dc0419aa5c1a60a122573f02b2924e12b47985729a6d90b43775b251cf1947a911a99459b27811999c2c3a37c8d0bc1b0da3f18e78a0d3aaaa7045c799a2343311bbb601b65a8f5a056664bf5aa3e6b046b39ee31870334dfebbf392b3f7b23552e4caefbdb19c21556415b0b2abb98d78cfa95e13e502afbc6f81bc6616c6398d4ec1eaa0afd42c498a63fdc36d76e9a3b1b71bf5b757de837c41bf5cb9f302180e0e3a51810772ad83f3ec4cc7d9ed1aff0418d50f97fa0db71d92de2f5d1570043ff05586d67dfbb4d613da79db4aee918f081fdef0bc023c1a2ff05c8f38d54d2327e1f69f8c645b9b5c047a66996032377567e275b954fe9f65d7288ec7b91b18253ed5cec5fd58369d8e8bba46a6e8efe29e87fbd102586d893d5bad9cfcf23f4c6326c4a432175e6d9773886d4f37f458d29beff467340114f57da87f5e3c135f8b8326d5ab7987c8765a9c1a3c98d1021c1b12ef343c47741b58949a6391a6b2fde86bf5c087421f70c4ecbbf31490c6f3eb376f54761b236848eb3e838336da70c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha2d826e387aeaccf3f5454c6ff5c6b1720dc35b76954c0242b9cc02875a3ec358c68bebb92327b0204ae5fede3963526fe7bf6eb0e2cfa7093b324f7ded2524a820637a952a2e6f8366ef399cc882c1cdd18ef606bc03eeab1798e929a7a925f03876dd0ea4f4f099fe8ac294811f482bf0d41b094e69736bb2abe553f807607a7f8fcf1510bb1f867f7336c72cccbe58f409749174105ca3d4c974279fbf942d915b7a78d3bc4cb14af44d6b0d25d4211e44e6ee71053b44a715b943337cd2b2e266a589d97df36a50c89e8ad5246851b875d64a5baac0d45908e22d5cce575e061f71fb10225e90dc28ac7af3f78d1f8eda9735856fa4021647d1c56b3446baf13746250afa7bbfe4fa10d8c902932b85a342a2e9c28da04dad7489c33ffedda7453ffdc2955ed0e5a165f05ba173b505d0327a13d0cc3ccdcdd52de56f8f3b4efdc27571c404dcc06eebe60518b5432b22ab6dbfd6328a3cf0cb0b41910ea271413e245ee479eabc5e5942ce8044352cbd82d825a940ea697e85fa507b93b5d4b4bcef5f9f32fab7c9ee38e64e9b220b6c827256c9f1970be37438a7a6c6e47301b3ef93a1cf11ba07aa3cda424135259d1a62a63c47d513967ce5a77de8581303ef6ab10675907b908068ba3b206b0f3ab63411157b8d5e8bda8f190eb5f38eb64b453f9d7d1cd48bbc07ca1aab90acece3aafeb9b719d3c8eac72bf08f6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hadcb1842e1c235742f7d680e0a4ebe9d50764008b394b0b4a9dcae56b385a8bb118e69d37b19b67beba831bac5100bc76eda5494d89e2fe3b2cda5fae01176fe54468a35f4e1a074b8298a55830b3bd949ae936f4b9c15a5b67350e1db6c4b195ca75588fdf4f7378fe054017ef49e4ec15999bdd4a394db1b5f470331b96cf0aee6549dcf63790ffea979ee1331b25b24197dd361470c38e5a33e342b4c73b01f2c77b4dee44c5b2b9f66963e55011be8fbc8c159907930352f97a98cc03c557afee28619f4ca6e5c347b4457f864398b4b41aa9ead6116687d0e210777b38cfcc34414dc78585c684fa13921ab03d683f5f75a30f0dbdd81b950655ad9c09e53af294350c80c028dc79fea27656de964284fc2da1217f8f0eae45e337498b00224bd4343fb6bae95d3607fcfd35aaaaf08c6c69ce4e934ac364add56b77e5f79e7b135a3ca2d49bc9ead947fc28e40d7bc5eecd57f227ac9770912d946a5562c9b28030fe15a37fe8ff27110d50096cab12857092faa80f962d9396067a7e8c8f5e3a6d7fc346c6f68e0e1487914470b813734d17cd39c4cf8d1432b75104846f9faf1794ec5ddb7ba00725a9fef3caaf175b164a86e108d2b74b94bff2ebc0f7f8f9f646489307fa34c601083134b67db7cbd3aea83978c69e1c25c7385adbbecd52ba9c9ca6867a4748f518cb2e9b781b7f26b06f0016310c4a1fe6d9b73;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf232b028eb90749dcf0836ca78e702cd3bff77baa206edcb1ebb207619572803f3070848f4856a7ef46b1162fcc0b05bf9ff53e3c4bab94029a18499e4ee960a174fb520c5665821fed971145aa7d71912c736de1645117f0c0b3abfa8a9ba3d9e98a7cd5eacd60bde9fc025af430eec9b51add0abb9f41a6cf40d6869935df1cc180be3cf56317fe59481063a781a2abe1c060d033fe7724dfeb030fad72e55949b46b532b5d44e722e6b40eb12e5cbabc978454bba5eabe84fe9c6de707516060f2e363ee3f093966c7f4addde1e6837797729f4ed784b1bcaa2359245ca32a277d46db2a487fac91118ec6a16f429ff7e947ebd6bbfddedab459cef142aad3fa2bc1e10c195922c46e40bef224556d58502cf75f91df54601b99e1afc4abd6a5a30966ba284d26d5d40a2c62aca3d9de35a357ec1e66b3beea5f28cf57a5a11c1ea6770272f33231349774e9a206b68ad2c67ad9059b01d9779522415efefe5bf4770366863a3a369bd4ed30d77862c9a48b7d3240d1f1720ae842e3179f9ca1cc27315572ed9ca18fc51285c4150c03864a4127e0585dfadab036027b47ca6d41d09631d6976f1fef534909095ea8d8cc8a4d2a28987be6743b8c3d450871f930ab0c121e28ba6a8e773d1ac8f80c9115a6ae1c34c61d0d3a057d3cd721477e527507cdf97fca1295c088a2af8b1f4693c109dfc1877fe92536f3e1f5652;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h28e99499ddb17e0ce92993ca8552786f52841aeb6c9a21aebf4b886d8fbbb7b9769c82f77141a643eb6efdd4b9f0a68cb548ce07bdd3f0b530e91c05c4c705020f4586c4351cd3b69bb7f8c2580a409dd8fc8259b8379b877e6279e84e26b6ef427063d4c2d445e7454e50825f6acec2265553b227d4477182b434a43137a29ae62fe174a3753622d9f16e65738ef0cad28ce217f9d7235d20ba586c09f0ec2e9f734d4011fe47eb3e6e4d7d8a72df371c1a4a3f2ca1a4fcfe4c667f41f9a588209e33b65c6d0b2251835d49ff2291b303521fa0df1f226e0feac954a99b3032240214c1fc423d7431a8afa02235fede7120a92972f7812f98fb8cb62bfb70b06e8654fc7b96eb722769959e67e8abdacca337653cf2cb29084688fed603bce992cb4e7071128c3c5c59a5a1b07f7fc9d437019484d5fd05bbaef743111e02e88b53800724b927168b50d76eed413025e9debe91716e8678952ee1217be8c9de16b82aec8e75f60331ba3de089e11db62a6c1f8f6d9779efba81162fd59374a3911e4c2d2e2d4176b4deae76d38f1387160cc27ed7681e9f55b0970fda75ef0745e3f389490031190d839c071f5e66e9398d142d066d3e6bb74d2a0a9c386630ca1595f9476d3535c9de21b286c1ee93729a776868399686c5abe09c06a57cbcd996e69db32d2f0858730aae669273340da7c6203e77adbe5cc0c7e4f5ca722;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h74991c2d68595038622bf4276db87a7a9b1b79ab063662a136eb05823f2c045a8fb9e9e861d28d3e6bafbb4e08e99ba9c90e5fa60777d41092767dd84ef846c27f296904c62d654b198178e06d5be6ae5dae45f29b66c28d131905758a02a1060a7caadd96726e6c226785d326f79e0b8f720543083922545e4e6060bb7676ef7bd4d7338099b24819d0727f8afa8bc8b32bc26b3ffd50a996d9a2f112260fc09e250de7ca99f99fef47942ecf2fe7d27e589fb4059ae4400044ff333ebb2ff000b6bacfd915d598d1da1ce1061c2af4d37fda9d5297c845b0b4870171c0189eb2465328cdfb53a2d0d5df57f63d83136fc51f5fc2c1ebb70309cf33da423cb03f9f123f37a1b036519bcf9f6a177a7db3c31c30e7dcea1a297a23ecc19fe9da415dfd155276779634b4d286edf9ab65922a3c06dd3e8c68af0c13727b3ec2325ecbaabdb8752ff901b86ab51946817c27c5bcfd8b164782dfb760928437b5aef09363a4eab1bed3091b11b8e278b8595bee168b802fac0e3e7d7c99d5892d0b06e80e1a66bc2eacdccea01874ca6f59d36402c7128af744c8622d7065ec55d91cea7eb088b7d127fca0a1b38e7427d0d7997618408ccfa61169f5805af2de7172cb73b1d971871be5d8af8b92f5bf97cb028ebab148e7125fa3b9cd1b3c2930202221690c987286115b0f9ca8ed0a5cad2f661c3ce626f7c2235fd69369641f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h99484d576ac899b396ce24fa39acb6949243c208ff35758c762a9da1296a5f3519a3488f8a304e1febfce749741530715b6988faa82277d1c36e8b7d59bd0d89f023eb28611e962178fefdc1b46415b5508496e70983b27d30d42585c9f2045e0d46387ab42152e8049143392d1a58e007f504f3c4c7a759b1fa43b94ff9fd07e929ecbed22c646fec839f2b5f3953db808e0d56ccb85c370fbd6d6ca6a16df1d0b434b6c227a9887edfa9b198c52757df9c0b822338684f6abe2d8151a92f6a1329207be33016dd1e3b6b8b935c8d6d5d715c199453dfbe3939463b38ba334e25a2bf83d7cc2ca597cd74ca69f53cea23e332048e66c684788c0c7600a3c08a3fff03e736242e40b81793c2b7dc2edac472ac4a3d38c137c4acef9f5743aa8ef7ef80b15ab29577f162aaf5d274f28b806763574fac8b6acf76a9f1eaba25dee3cae4cf350dafd448712fee82ea9f222f24cf828af78fb0e13b25e51a9b5616fd36f920bb49ebfafc892bcfd13a1a0532ed040b455d488c565cb195a9d73cc94a96d8f18b6c02c2b4351a3d37d39dc20e137d50c5c58c40c7e61c2570e5071b9aba7e54e788fbfebeefc77521a86d9754b8431f2ee6327ad6f0ae4f244e0204a0af0c9c928a1c8822c3a090ae9c34d9807b760af69296ec6592f45104ce04a6d3cc0f8ddb9c6f393fd82743ed1dfe5e39ee0d8a0e7c25852a4f40f8b720ea89;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7a36253d6a894c0f28628fbaa5cf0275326606c5adfaa0a7ecefdc2fb5fb58fc27add7dc202b95a9016bba0fe53e37c33ce6262b72c1d8e0908b7f8b2ea1eba753dd3bc30f6e3f8f895ac1d3f865ee9739a6712fbd6e9ed4bd467b7df65a7f347f5475e4e5469a7b3a0d15d9e3872cde6a3962406d4c5eb99ad0cb478c01292d00eac02858a610b8167f620c0b32d55f7177710084b5c784cfd029954894b09ff143f382ddefcf4fd5530c304a55cc87c34ae1c8fac05f77365bf5560be8a9adba353445cd3a471951d06d0e817da0bcf001e63ec16dd762c5b262912b278b5ee4ca1633fb6e94cbc283d353e478a11f583716302a9dcd241dcfaa485443fd2e5d7eee145eba6de275fcc5dbcd75ca9e8ad0140128818ca2d51131de97214dba5b99e4f706e00a4181ec54d911a5afbab4215ec4173c057c0391378bbb9ab56de7af6762ef524d15512122ab7794ef6da1ad76702b3ef1576253ed48da7ee977b42e7edaafabda475a198f04e8ce6b515539ca8f0c25ea79b0ed331b76379681fd38722a65ce27d838fa74693cfd97d27f062ca139dc27ff388fd01cd7820dbf670b96d0e250af999dae3d56be50ee3b09322bb085d9077bd62673bbb16e5f410fdcadd9a9a04518ebb7d8487e28c3ed1e3ab326643d1f431eab033a2d14754abc750c800de991aefb9369bfdc82a614b0eb564bced9abca48de3d009e52dcac;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd8b15f4fc7ecd2598c69543099d2f0e3740be22327f6dfd19508f557538a2a732efdd19a661f93b370ed641dd94139d4a8bc29046ea3776292e350cf3b7e2dad7a8fda56f956d3f1d809dc5608c696fa057c73b0527e0f29bda46c2fdb80e3658ad0f8516b2d52d6015ebcf34957ee65b3a382ce8fec619940c8308775526a386b067aa389a722bfa6cae91b26aa31858b2f2e3fe1fd239921dab8747088b87f58c02d2f63b3c629946ebe653815cbcb2f47db65d75dfd3edc04a879bf670e787072ae0a1b9c8ea377a9c9ef74b006ad1c2e2180dd850010f2c7d3844969e4faa96663a13fc67bc921a8c0d210f1acdd46163a75d3141cb4232c71a0b3454a34ce19e03e33020829dc4ba1ac31e98a201314f09eae84e70954d18915ae0dfc863e04ed48f5e6021ebbec799f585c6c04c32e7219c02f15c9f53a92511fd480fab10ea14dcbaae310139c66cbc3922b53b97410632926cf3522d53045c754fe93948b4e2bff41ea7f030c6fc4ba03d495f855afb9c36725e38f41581009d76e4338b9a114031f60b6dd7fec1b176b41df5aefce4fca267d3bf7846355fcd6650f84f87d6ff43d08cd55db1eb8df42a3ae9c728a96cbfa7fc862f63d16fe37ae7da546b290c1fa5105cb2b9f1b803703f8f805e5ec73ba6f89e4a9eeb48dffadc33912b8709bbe1cafab61a2cbd4540ae590f2441638b8a00b1d24771e6b88e832;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4f9934fc674d3428431a7a7470e97c11ff70c92c26530d39dfa9d54a4a77df4db5ac7156f1500f37e06507b5ae8415966b3f21a3f4b7ad1a2daf6cc0bb604587c7c799bae7534e10c34e3a00579dc992c136d64f6a1e13a524223eb718e21db89a96de52a35a83d0425fa7f19b281d8f9d56ea9e90fc8598dc923f4af92f3224db3e829c20733b10f1af925ea5d8e8bd5ac397597447e9fe03b0af3d683de8183664cb0dd8fe0ca27b3612699282b99227e803032aecada8933238b9f50af43151d0ff4786f5de40afe59674a616cfe0a6800f361998d0f64740b7b622c47228658b67095d299b736d78670ffc9101f175ffceb84b8de7d2c0383b6d651c1f450a2de7682f97b47aa593a5a3cef13df123b47f71440a57927a9ed1e3b3d2dca669381e088d42c780b3b8c2c01e281750971361a462dd7d64c2801b4cf4d6eee491bb8db788d53681654124c1d0e4d4635aa5075e24358fb3e6da8abbadc8d01f5cfc3c578df4e13a259c0258fd65b2e7ee46f0a83e0f7b27d56bef7af056a978f61c8e67b1642945616c69ed849fbc737ce55b9141abe900079061fce68e5531821176cd2f21efaff06c2ac70734ce64ce640533784a6400662f3a0ccc2c86b481aa97468058ebaabaad57c5b7752edfb71a85008a0bea8855ec3f517d83796e08cf8065ae6e9bddedab3bc7d0616b675b3ad12682300551c79eff69b038f02e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf7a5762e4df7fa53975041ed92add03256ce6688572d5be70559edfd1f4ccb02e99759187368a2c569b6e3bafb434d9885a7abe5b48dba1e48d597872f10184de61213d1afbd4989ba6dc7a49e01846b5d6a443fa7a7200a06285587a84045903296b3e618709f948b77bb115abde626c618b338c07bab3417ef38279f66b265faff5eb5de7c9a947e9e0d1afe139b2be123af9d261bd28ac96a6d020fbe3442ec123aa850afa5efc25308358251980cf8f7ddfeeb937a49431b4d525229f81f9524d98504c262d37859db8657e2aeba4d7424bcbee5d845175f858b26df1c4306b2dc5c734f22cf736b5c32b617042258b1f2c8172fd004229675df8741bca2bcf532be4dfe74681d6c2861d30744a72b0bdc777626899089f03c523dad21695290d6e3df7c560f4db8a24276b67bbae28ab7ce8459596deae3699f95d3e1f0c20cf8fae8a61dd712c6c0e88273b55484f99e18730fd95ce48421c17b5cc2c61ffd609859fb44e724cf9a4de730ad99305589cf2d95639284e686df794422a8b4948d79cfcba8bccfbfa988ae4d731887c23c3a1776076cf5609460d7b8245a615eca0f2df77f031bb0f9ad28af69912c07699b6960b3beebd4d47e92daead69ae437dedb7cffe4db16c63353f0fb4499d55755fb2e85ab7475c393ae0eff0a19903807984c6557b4c546958d859fb5cf13dfad179ff27a041bc81da3c0110b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h16c18ca7639a609c1e046a9367280714f70db552b9106f0e267a6bc437333436a0e29780729038f5d84e0c1c6e6c359d42be49600fe98452d2ec245e725c572a9956c222ac608d588b22d5e9a66455b3d2a49e52ba7dfe300a4025d20d79f58f4d69daeb11e4d4110b8d6d0c47bea3a92d3c8e1cd5abccd35c2faef478d56affe7b05532b2625c8f977d50c9ff7cd9d90e41b6ecbe7a8ef27efb0ec2e280c2309561c6b101225d4e7989c48ca3c50c252f38de184a2d5e83ae0620f88f66538db4e6cc5bfcd98aeeebd5bd566806bae991ea0df6d92969ddd1bc0f76f726c747dd514bbd322fb949b6d6985a732d6849b9966a2b116c43df9b8f4111503d343fbec9a756ea97eff253419e7713305f90c182408d2a150cf5e37ea36cc085e766bb2887f4af1ab81a461f8b7ec2ebdbd0c4f2fef5613d76e09a447e46b0403008790bd674c86d24ecc99c05dc4b9bcd0914134c5eda4546e0679d91ac641c4521a072e8ac6c39002691a683ace823c242c40783ce4e9d2b1dc418b6d48619b80a855698df6c86861c5fb16f32369b02744022161d27757f8b17de51afb3dc3f3c3a264023a99c141a9e0f14758177c55706ba4436ff22f3019235cf75d80e97a6bdf82b137f76f8185da810be3b2a9ee0c8781a441d7ec00bf384ace8913ad765552b2aa785ea1bca0a89d5e8ac47313ad92f767786319e72c67d9b964b72b5c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha40e8292d4ed61d1acaedb804be770260e1344251cc6438ba13896ef2021f8f1557888462bf2384f7d65358c9012abb8e3ef068a8199cbf7a0bf24f4373d89393e76b59cca53aa6e25f93de77400763f47465097a88724f020bd28b343c8994641b613da3ff523286af180d164cfde5af736862d19daee32b6006e8958e69cc20b3bc7de99da352b7d702b183932683ea8ede484517c53f5af6e9a3d65f1d0ea7c5e2fc9e7018b23bc05d3bcca0ddddf62edff04d71fac43030a169ffe3f007ae6ada93e90074752d89afe3b5410ad64259773faee753486a4c260ca9377930a5205182e1def32884fe9cc625c5e333941923e91ae617e3a9224cd6bc7116dc9e6620dddbcaa2c14ee6a5307ece1a5bc306622faef15843a537be891455ee6ca9dca4196ae309df71426b6d9cdf0b2a3bedd57ac5af013f82baff4d7fc9a7fcd58517db8f597a60451709b65bff8d757445fbb43ec8fbde74750758775c8b17ed7ab8184a5929b589816c06ffe0596ba294be575345c8833fbb696f0176d8765529b6970c3cdaeb2fbfcbef5c1ccc93a834dfbc66c22c42145eeaa0b76591096961c84ed087d5e0e1d30434c272f70693f4d77d12879b6b58be9b2fb2b17c23fa850faed0e8ad6edd668dab9c570d11119e9f72f78409f7376d5dd6d6fde97db9dc4f5c7fcc0149b3b7fbc24b84353b098f782681b24dccf1e16c2d741f84566;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he898fa7f52999e8cf55e27228d1f36f4d3d3cecbfdcdd0c4954aa2e10ae75d10b2f8bcc71febb8eacd88ee503c31dc7798e98fd4273743bd35297423a65181bf1450e6b55e9ff7020241ec0501b90e0e67eee316146b96e2997fde161c561f8252cf38ede3aa6ba047da44fa2fc3659e455be6380a9130644025ebe0734d0bc01178ee446326ec168ca877f6f23c54fd971b43a7cbfe6a2be744c17f96628aa32b8f4634e0428fa2af540cbfb4e1462a9bcce9459d88c41a859c4c8cf313c3c38430d2cac7b37540101caca7250863749f8b771551cd8009eb28b68f2ec9bf76d55d33aa79db1cf54d18febf030f9c1af94926b01afbada10b1dbc8bfcfe0ba1d03ce86d62e462ca5ea45ec75f620f6617fa88efe2dee28f549baa4a595baa14fccca7b439272611a7aece65fb7cd7751a4cead13ed2892cc334e361d47f0653e67176bb784fd3d323e56fc67a9ca17e7c768c2462679caacff7a62aabd13989729bc755adc152b4f0f9c2e37f6692a822217cc0ae895d86ee8b85b8a3b298ecd2fec4f34f3c4db4fa0b1609ec5d213b62ec37e7d9844a906deaac74dc2807d1e810fdc5d298eb3bbe535f9ab2cb21ff370cb78f913238d31e80fb895cb42c299a6dea85773839a7726d1a78ec2210e3825f7d35017d0cbc1dc22bb02c807648b2d0f77d821cc519875f5190c5cb08e0f6ec72a2e8c13459ae2b528b9a64511c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1081f8ca4bc0956fda9cf255a0e798a6f66841d8e5a4c38593110023474859cc7f7176150ff3a1951b27fbec0c8d93d51a8c831d00ebaf865901eef20c085b3211297ef9626f660c87ef6891dc07087f4bd28d3f15e08a464acb06524bf7f06c9df2174e8ea2d47bbdac9811d149689e329b4d6c14bdab44fd80ffc0063a1d89fd8b684ec593bff183dc0d4a7ecf48ff4899d2a883584cdea346e1da2d59bc33b50e415b4b57cc632f31ff34b4ed11d0acf442d28dc1500317f7be7a65ab7a8079e0c8f97f938cee2a67aea885d522b1df2e2fc7a1123078bb94d60829c834554e728645bb59347167869ab835dfccdcdf499e03e33a8c6d5ba6ca48200a3a748d1c13bea11e72a59e01fd9678bfd51025d7c1e00139926ebfdd89efb5f79b2645c6cea30fd0c661028620bf14991d9e99582f22f11dfb650af07417bce86945d765136ba0b91ecc00a77c8b9ec36118feafdb6f3181b536c9916263f84345786800c93a6a71bd23f85631cdd6e7cc8f7d6a55c692e43848e2b17d4b3ce73f85c66fa7d6de8f2998631f9c2c9c2ac7829e608568eedea16fa4c862353cbefeba85479aa170770afa26ad98be4b6e25cd423777a7fee1a5591bda0a42a0953d917ad0f7acc824da94998717a5d54814295cedffdc2c18bfadef4a282126327cdab92ea904d71a7eda6662c7fc9efde8e341e611487f1101f3a3d94b396bb20b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h15a66c0e649093f8078608cb99a2956831c1f671c2d1f5a670867a9704faf17e2655691ae916aa0b893de9e46b7741e7c52b9cb5abcea988b9a8581c755f91abf4451532f792374c754dd876008cdfed19e12ad307e96b5fd3790ee75952d7c3cb656ff3cbb18acea0082032a37712a792deb187f4b2b5731670e4dbb2f528c61a32ae331d87029e1e7cb544b4152fd0ac54b770a3bdac08c5300de37fb68e6a4e125a7bbd711655fedf7b87159d7c521b635fb5bf93bb8230b27174021a5d011349ad1429923dbf2011d406db88ae65e4ad7be91271b77a44d4be4e6be288e0ccfbf1bebb906bdea7b910c9aff42d334c674b6fd1c7e6f5fad2875c6e458920c276067483cba5795b54491cb7f629f03bcb872460421f9e99af5668531a8904d2bdcf0db4018a70e1b08389c753565c7d8c9d9f978c199567c6b922b888179afd3edd0e4f4bc02cdedd10583c38c38f737b1128489a8b6a6c729ef8792b1e4b3b043271eec9abdccb3c46875685335518806508344fe8628d4c803fee4a7a1776c3b6bcdf3ae5f8ca39908e7834c08b45e9eac76049531cb852147951320f3c7d013260d9cd24ffd1f32729769145a91eceb70902703a701e769e228ea4eaa54bcf67c8eddd2ac1f6ef63a1a913d226018abd9e46724c7e554164f56c3742684ce4c056bc430d0e3f02d1f8e651909a18e85042861fcee6d4da5d6b4f9c6c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he254cc3c9ef49513a746c2cb3309e8c1d7cc9b97c1fe3030a280f454c678f2d7d7061bc4ec9de27a596e10a6b9ba42c854914b3da87b92375993a4d27bc0b362f7abdbaea949d414312378ed0ce49c1704e5ff2beb6c85fd98df215179eeed75ba0292d4477c0675fae1f2f7702d06ac70bca6a6ae9308955796cc404b73aef89b5c777172689843701bce6f80973527e65f3af60c48987793abede6f49a44fb74accabf803a89cc887b58bb76cf6ecedc5584a6bdc81e2922cdf495b0f26b84f64412765fcad6fae7bc10f608b1f433dc3a012f0724d708846782f1f74bab7b20d38c806434e938e7545e8cc94e84a1bf9078657b022b2a00b71e48f6c7516eaf20c47b0cb777543d5581522e3e1ea8626c1c18f661e945d64c6e506f985073fc9d6f44d22072dfad6a3c07f97084705a8b3724178c5adeb1efe4257f2e17be5d26f619c5bfc33b3f5a7653fa9620d7dc2ed1723bd4810d6054f8b4ba405bdec9c4606446cca61ec78521ae80341dd25b0facccce54470c10e7312534246c558b0723795c8b851d47316f172e1758746d3b8278e517df8bbcd56bf6765d4bda82f275c3d0c6a297fce6969625695507fa72d15c88d1bfc5fd9e6b08d3c681cdeee0b2630732d282ecf6af23f38370095cd561023b785966e7e2a5fcbed5d3ac0384ab16a4fd7bd9a35a6420e159db4faa08e70e892c0794485dee5b9de81097;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2dda0ceae16d2926b15a5aadd690117bc97d87dc5df60bc0f7fe8116a0caf7d5b6d6f2cd5d5764b68629d29d65e6a048b1a948f6cb93d4280d5497396437d5a99a2a572b8bb8f8a917fa6a71e9fb0d3ea71175625d1b970e7b73cb4c4a20b95bb2707cc477d4a92849bf34484c7dbdde2d84658a87d05219fa9ae9dc85c7a004ed23c8d51fa6618fa804be96e6710acb1736cbaf654da32c094e5703cecb0169db9375d67d319be3f7ec11531bb625679ddedfdde17164b9c7df2434d17b79697cfa23d540144d367a06f9d5b8a8c3e6106a36acb3906017716aefd7bacc931e7d4c147747de8abc59b48a84902676f5ca99e5cfbae16f1aaf2efd99f74da6dfabdf76c0a0fe93fee9e9b2a872ef1b7ab0849d38ab6b58a7a538adde93b2c42962c82d3c7376f586356a6d6983d584cf6ad0a91b807409c4c8ee4bf78a80db10627fa4109c513941866894df61c339300b547ced04b26bd0bdd4c9e44bed2f9361fe6a76c2aeabba2d8e83cdf8d59e1515a15ac66f9db59c89d999a73b69ef2725988f0277c4c1a2e7fab5b0891916bf686ab6dc1049474e4cecf9225cb3275c758f5a96df17847a02329717b359b5051588c99902ea5f2ee7e20f80af26e2cbbe497a67d6f91da5fa84ad0531c7eba506676622066461db030bba98b4254341687bf4e1992c01254fe6b3aba6d9a3626dbccd287cf810813964b5485280a607;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2bcffcf8fdf55306735a0ff4945250efe15c7757435fbc231becae7d7fd681f33c2dbde7e52a2eaebd2edc76b4a7d7c9d5fcbcfdeeb78b1bb44c18ccae0fdad1f40fa489c483b437214f88bdcafb7686f0f96753338b0c591986fc129b6f03e3909c1252e2b069c0fef95f0255014512aa86d9234cd25cb91e9ac4a70a83e4bec87722f43bf5861fd5e38241384ce84b865dc210c90f7b0d5f9d028893879205388b1f6861b729cda14667cc94dbf136715db0c3c51dcc2e928ab06f4a105d2ddf6d6454108d4af6d8965a456a82084da8bafb25322756faa1191a1056449b6f6f863fea2f16a4b48be38c130af544b824099b8ab66cd92495d0278ee2e9e5a6b7308b4ba1fe1de10e554b8989812b21bbf0836066d5374097467d44655d6bd20e96b2a30abfd38a4fb58c388415def9dabd13b82d87ab3bccbea80c0e70959ee26001abcd77aa769830b6c31af45c9f2331be7007cd7b62ca06671ba6ebb7fb57be9613cb0cc3437460c3a36f97c8b04309a3a957a17254b71e3d96edb798e8150c56dd0740c977a5f7ae22bd63b062f7c98480fe2d6f5f3c7dd08120cf12e26962caf54e8e40bd5d1eb59b9d8b3507f34d55ec898713ad0db548b19d6a94d608b1b6db4a006c7b4d4337897c06ee9b2f32d8e21788ab7f7f671de9cc623209f7c2a6b841788f4db4a94d5efebd085981b9bb0f37b57927dafdf2ab5566b3a9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h43d3d98ccb4f7f401ca72ce3a0b4be4791ac3922b9f124809502cdca128fcd7b10f2cd9df8a4ba97dbd51816a9d554bbe16e7c8252787a60c5ae156fbadd9efe14c3b4258f09d59e1fc193f1729d5d1cec25aec65406bcc3f8138676dff419dd21922324f48fa421d473ed2595016ef9412917e17906ba3702214f76e6f9064596220dd3a1c08967de1e3522aba336926eb84a82302c5c3b1fd3595f194c50c3f496405e4c3138d18a481cf9814924f1336c6c0b8da6cff27fd97cfd469d454f95e1f0ae2849946403a51983616634c94d8f8f5c085b94641e828f661815de040f496dd066f7c5827fad9a67d52aaadc6ed29e7665693136d3bf7943b3cdd26864be18e74d5f85e36e96d01745fe55352b91de075a7d00040db0e3cec15066db9dc112fb5e54382ea9efd15cd33b5e4abcd8314f9a90f521d6284a5469bbb39977686a23f672b92a4c0f88de86fbec92947f7cc1608404c36e9775cf7dd8c55132173e8af8758a2dc01ddf798ecbaa2bbd07d0f1ff58dc749bd38833a11f7bbe2ac3cec42233343d0cd0e364a7801fb4e0e6a94e63e4ae093326acae5ce2c008b3f38a85ca1cb2f94993d5a08ffd89ca812c71914e344724da77858cec6b25d9a651ee44415bc68e60ec0f6c6f112215619c88c7c79821f4b0620aabbdba7ed5035589d51fb686f04047689fabe21d6ce6876ec9496617122e143ed9ec43b95b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5983f24fa4f3b1657dd3adef4e0b33169e88966c2274958e34b8ff834883af8bf1d7ace91c4e31038cadd5a8547cf4240569d52135ca4ee7d83b216f199b3dd898f41e748f292419a043e2f6e8751ec34c1afc6b1e5534f72db1f33cd92d3133d7b26e7a063ff230beaf8a64f83d70d859253ad6088fe0ebcac4c0e161bc82a14eeebb7c6615c0342dd572a95b38efe4016cd26e0cd43af08d57356bd5d799c80e04834054977e37913513ff19e7b7a709814f79daf118fb67b4362c396b2146adfa84992b838769554b4f52f2ba7b7abe535a745a197cba1e996b4c64b096419582b8f330cdef0895702e66231ca6a5960eb3bf6949b22e8e63ec14ba06b75aecaf8e516eb6165d4887a3c99614eb2fde24c695a8e631dd528bc2fd2f518a18481a0bf0f0d10fe4770f4b73aad0455cfa6287f8a5a4ebe053d5f46f4aea72fc0b18e4c9b422347f546b6e7f850d7a026cb85dc822ba29412bd276a3b4b92f87a8f93e9df813199cca5c1b4868e05ad2381f4a1c368ce0e992356834cdde6a5bb14b35c6c5ca5576fed03faca257f5b6a125fb39493a8b4263f04a9a356200c6a5788561187ed6f465f758b4d68652a2fd9433cd62333182295fea948079997ed6550f6eb5f4fdad2a39107744a89d9014bca7f95d55ec3f30a76723c7154a5dc1ac654b60dd2d5ccf139449d769b9483973622c82d2bf33ba581ea19d2e22e7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6ca0cc3d37a01d943699581814330ef1100cb4625174bbc9ffb22b99c420641ac804a01e759a5d9b71db2a0dfcfd7e3c1ffdc8699862a204dddb601f5f8b9d525d37053f93e2815c1c673da3e136c28e0cef6e5d1d1720694d4b85d763419bf5ec84f4caf9cb2e1326581931491e53473cbe508868eae8ea18a519d82f770bef2a21555f2f7b3a95ffe7f3cace5e196edd55675980bb69a8d7549f6ffd3d51d3ce44d45de19c17861ac78336d6bac41d9109ee85173d929f15cb2c64533cedf21d182065be42cc75c235eb93550bdaf3f6d14d8db3d019eab6f080ac01f9299335e1954c16f1c94be0f886b970789fa97a73b7e8832543c32f009227fe631995f15165126e1b1ae42ea1ebeb89c424d37fff7700fd9281580f3cce335169b37a8b3ba2fced69a01db912327a3e9f5157e16fd0c4cff864b214cf3ef244eb8e7ca018f57c0f5848045bea882ac6ab8a78249dcd8c2a0b7e0f95970e1fe7cdc566763233f1efbabdb11ba80b2da656294c95549dc99670267336e4004eae5f818f41e446114c37b9b238232b71b7c1e10fde2aadef7d763b9fd54b4854dcad3dd4a47b508ab906796b93da5630016ce8287378a6da649e768f6c4ffb90392257ada0d608966de517ba2b841787a8a0f0c87683949b8db12bcee337e8b3778e863a81a253ac3c62a9ea0d7b3dde1c6a8574535ca928edbca636f07a2855e3341455;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5037b77c5a31f427b96fb470409e010de655c02334e1867aa7850c1d8eab30f527d811ed20f051ed78a8011b7f885006a6eb10f5eaec01ce62e8da6c77ed83befff1151af58f4dbb542992328cc01e49a786470022d50ca81b4f0ee0b48f60d6dfc1c43c11e18cca9e5015f9d6a5a396294845575096a51f6078e513245bccbd3390841e59fff15fb358597299f44bcc1366e0cbcd3509815d0d5df3d026c601805faee836c7c85c76c420de5a68d05bdddae51328e9e3cc1b0a61369483cf65e9f82f9684ff5d18594c7311eb5422e1036e60098592c71b56b984a10f06618507a4d264f4a3acf753f9a3bc62629e4b28d9a555b7303f7540523bb1312c832660f1e8c78bace36d070c476946b7abc7b64a52cd69db0667947d66cedd6c2adb3eb539500c09304fb6bfda43532ca06a6ee6731f74e7ea57eba5e5a5736a00b52cb17dff092f51ceec550c81b9f5086dd8115c98589ab15505a31f79cbcc924ac0786556e61ce04971f8ba1ce63750cc032e7c81c29abf042bda4cad34cf2ef11646a7a94922609aa6f589e6d693e22aae6bbf6d65be1d8d971219fb0271339cae66677cb749cc64530eae4e4be8db7e69106f055dbc03ea4dcf930d2c1448f10d28ecc891cb3c19937b3db7ae72ecf8a6d0893d08ff7b8931940bda1a76154cb8d21221ae2859f7416043f356da81a6c446d09e1790c36e655f415c25f28371;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he23c51fad6ebd1b8a003911ee8dbb0fbc2ca1105f081f78958a12a8ad1e4042ff6013262870b66b638e9857a28c09fae16764ee534be4197ea97ee20976de97bebfccef81f41cc39a5633aabe77129baa4be452150ec9a43f1650ed29e7878c60cda585953fde0ec04cc1c92c84b0b98f01a141bc7e6f8a839a20e40c3942db1fca6d4d432cb4551dbe3ebf8c4cb3090a966a374cf80d7ca21dfa448f3fc79c984ef687c479c80736a5355611b08dd2c2113b1395b419e05d1bdf694b2f58ad0fe7c191cd29169fc285cb61230bf756403d69fb8e0ced25182f5e63b870f9bf9a09924e00b29f3318c8d26799cf73538021ba180fbc9fa1df57d6d4d002b7b9d260a1ad993c945ae3898e613dfe1145e39d4d51a736e64ef0e0b632dd19880670aab804bb1a02a4c7d3b2c0d5c8db0b358130fa14da8048a92a402d42f1ab1b884b48bd529464bb71ea18e07545aac113efd692e28aa6a5e1342ab00ba04cc4d38bdb765ecb0ca7e6757a7ecbc2427c64b1a7a6a55b13d6da3917f92ad0d9fed6eaf48d8f3744623c5573347693513b60e34697c120f3d95711b3ce8baf5dff45e409d6cc396f13bfa35afc701d3a1dc654990bc5fbba53b6860d286193af9b10b19083b70fa9a1b74f7f56bf2360b4a98b02df4d0e37ad46640d98664d1d102fd41684a14fe5be08df8961f2ffd6bac154ee3463035b7fc1c0b038c6d9ce8f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6dfc1ae597534d55d3d973cede62f86a8b2aa54b1d1be54f3f0975c325977dfe79e8ed2be1aabb6486f73466ec237c7958680bfdedc946f873f8d8b904662cfde1db3951672efaf4db25fa25d68eb467e283272a053a116ff85c1f48c3b1b0b93f4e1b00cc8d255b6d1d9f3842f1fbf6936fed3cd4b7e4b0339ea5a1ebb7a158afbc345d28161441477c771ae504f34e339f2ad22fa822f0c859bf904abef4b36bd072f50f1c7794f9fc252c7f94d04ee5ad096525e0eb01f02fbbad6613d511304d507a748e27c1d06b9934ec5a19a05f082e0d2537e594f76d3e22f6bc68de1ecf3d593cbfd350f4bdf4c5402a2f5cac7e35ace6fd7d8247712ce35973764bb420b350016ad09dbfc20f08a20cbfc07c8365471da98dea20e598d44a2ed168a26ae15459d8900c96248f3c21093cf55e5406ea6f8de2f2a83732da2aa9c8f7815f92817b9d4fbc9b507e40837345557c5157f04f8c872148bdb341fbc004a67c81f4c43211d67451b144095b337d25f00a2ef477ac0823d46df646bc6b16fd5b2a2ff4cc351c80a004688582dfd56caa0bed6cedc2ac3e9d0b84c151d10a02cc75f647461f857618ccc6a196224cf73b40d94fd30c1ba5715a9f973203b8c39bff6efe5bb47fa6ad7d430ec0694d1245655a8d12f411a495cea1efab6be1574c722ddc9aa1c539a8415cec37a4dadc56f28ecea6ab3c4d932fead5af325b40;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h184bdb26a6408049b5eeb541baa29c2e56b616d530c5df9f32e55f42010916c9019e95858d9de2452aea71f47c62c5c1cf8c7cc7eae41351811207bcae2c28c94436f4a24c886d15d88d471b3319233afb62880855facd2d2e2a6f01be910aa6015d742cf459a96312b7e0fda4241dbee2efd9f3b1be27cef54814733f4fa4d42a75531edfb81da542bb39d69cc2f8d60fe620fd70d07130a30dba8098c55ea97d8d364aa0cc39a8a5d1ea666b43adc2b9b7498e4eac2d6da4a56ff9b9d3538730201857c42c1f90aff83c23ece1cdf176a669798ecd676d3475a1b1180811fef42a74a1287c3c824c6849d8654b2c6be35149f5cd60f5e06376aae820924b16bbd40a51294fabde9888e0bb9c82c33ccacfa3bbf23cc070dd861ffdf63e23112791ea1cf7bc17f1b836e42df8dd63bc43061bd7d40e809ffa39f93c779c33f0e528d6bbec3bd7c159efed9744c3b4f10d17dcf78a74f28b6779026bc6db2f724b9d187498d5909e37529ed8821f1c896c89b3a6669929408fa7a180cd01c482892eca57d6c9223352e026856a0af06d423c74fc345a1808960a2d80a370f7910d94f2db5d95b88471e3119d84e15fa75961f191f359a246b9c0f9bfca880ef8a6ed87bd1b5d804d7e40cd65ba2fc0bb0a63ac679b4792bbc2784ca7e802ac56b5af4db67239feb18896c2effd263bb3668e447e94e7601974b66e11cfbcd58f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hea1f294e59ce3e362f1552abe6260b15b2260feb03b9860b840efb12fd1b2dc87e74e9c5428807d62384a3acdbfd694a9925865c51f7f91b7ae145472336f683d3140aed30ce3a37ad2c531693c1dea2c3e0b923a30522016a55cc234d523cc92f5354947b53836545840d99ceea13ddda56f1900a1d7a3de5891f2f3329d2d53991b8b6be36ae36a0c4e54a7e0fc76ef4966e5ff7ffc54dbe1f24a3ce086e9596172166581b5cf70dbfbf35d8aac28bacf065673347c56ca6585977c2a1eaf3e7f1809aad10156994339ed38427992f9dea820bfbf0f2db53e625efae58cffa07d6869ce0c9d22c501c649e770397579c8e262413f6a8197778794bd55724f4df365d25059c719357df3abb4a20d8b118ee01f14d1c4a352ad9854ca8184149b4d57ed92f5c17aced8b4b66e0905b39a07029e24e001b954505b9c29501a8fe9c21f9d3876402cc6f1cba9302099d00d43008cd5973de68d22ca04cf1275704bc269dbd5a156fda78ccd7eec0d0578d25075d1bfc687793a079df4ce6012b0162821ae2b46f3514073d0b862c8f655c0a8c1860b5e7263248d4956decb094fb6464071239869a578f9897883e1fe2e7b680c265f4bf60f1eaff3f3df5219cc3e4dce83102dcb4bb247599633836b9ec83c32644fc6ddc2053e70d0e34a3e6e6fbfaa0cbab1afbbdfcee7e25776234efa728b177de4a6025d0874e4e1485252b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h64e35dbe35d1e63447917e1365844cd578d3f471ab38de8a7249778c23d0f5950b36ee55f16f40bbe0e3a6cdd52e4295a85828d7602e097c5d18b6d434d1732c952106ba1f189fef95d6e46dce78e15c2d7c5d74074960ace8a7e8b308d59d7210c98d20d5e60e1dc9f2d976a3650f42a710e34fdfd6049faf43dcc05ed20d149a36feac28a4ef89559d41ec85fedf713b9d8e9336692a21a73372988d96cd82777bff1ac89d1619ce4f1274cad73752c036554420bf48105eb070c5ce08e86cd9dacd00289d7ea29a0a75972bb12a0a0deef7105e20f66c5cd40216d494d5994278281e527e264d7ce7afa9824fda7afe9eaa459508b2c72719c09451fb18f561048812b65dff14289926a2f395dc95f50b423c82a6d3af17c0cf1cea32a41076af3edcf56a90f1767656549b468044b4078bae4706b2fb7f9839492b4985d5b44fb9fc75fbdcbab7d01e5f8ce88e86cfc8c7bc23f18b8fd901a2e29d893c651af0c010be1213da80ecf2e42cd4501e5a9b1f4005d3d39c09a4a74bc06208b15b1f1608d1250368ab6f84da73843a23b99930139f388f5de0570c63de86c3738615297818bff787b7cfd07ffc447eb9ce4dfb2fc054fd3be249514e43c1c6bfa8fd5a1ee4c42d973b45ec72d46048aa2aa1b55b8c7345ab1bf11fb0a834f430ab8251d9efb478f426e9d0dacad60541c07f3a549a8d0e86a7cd1b9f27f32a19;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h11069465dca243f24434be610d04ac44e01c6d1c099eb28829624fd4af4cd5b59d4adb2671491f38bc5d11cd1a07a21a6be1901d43f9d6458352d87b666b7ab616600ebb79b1652b53d674fa91838bfc1b92843adebb3501b62d68f7c0abc0681c020e2c4b222d518ee81841a8ac8602d0390726709c26704843d287ceaf7814537d67b62bb978cc5d2979452fe20082848c4f2a793a2d3d8d5fed5553c59b3a18ee5d639cd85234514f6d8ca71958d9991c629d88efcab7358084226c28db7759805241ac65da341db2f4cc2ab01b01e7324dc0ae6474b13417999291e023d6292663a0cf80680d43aaf5e8fe67edeaf8e54e6e2cd64bee44d056038d5a7db57fde87a8a10071e5d5b23472568cc4692d87b36a69d23dfcdb8d88193e1452029df75e60b8677db76e898f10ea5f5886a49f1aef30a996743c4c8a8d76c4306e039135cc9f35f025c98dad185ec2536809697979269a48d3b1b30a493a21a3aff53957d50ada031b75213739b4792f4384eb44ff47fe5d772048be09bd68ab690f7c28f6c94919e44465d8d9e3d6ab7f8f3396d9a3f35001d75cac08a621f7d9e7a86ffe92c3672cdb83a2bc17eca39d82c0a3fbe4f8c4c6482a41e36409e84a57fe4f44f704bfdf2028314b260774f1e9762b7dc006bcb2d30ea0185d653ae49b0bbc33c38a3d4727b7c325f2a08c730024f65aae7348a22a38b8a8ec3326eb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h154fb76aa31248a51a8368da357c97e3908c2df98fa101f38470f947a00b6b68f210ab6816b00d90d6922bb223ec243876b8ca20f2d47aeec100abcf5731279418d19367db0bdfe54839b07cfd8e3727950c211dffcf6a6e4e01b284a24bb2e64fee12cf49ac351525d5bda9850c06cd80a9561457b536aabd9f2b18a2e3173c7e5648d93433eb26b30db6c9ca80517a2d4004428d16c862a72caabc31e6b1c5e1a3feecb10ec5f6b860844085d3b17c1367a039dd6ec6e5f1a602e558bd6d9936957db0429517c3ef2b7e587008d5bbc0282c6b93f72c2846b9471a8afc537bc3d9f9f10658762af9859cb466ed727d2c561770c19d556b4969c8e22f993d5e0fca4f329f9575e715bc64225b8bc4d1cc7b6410b85796f69b7ed7cf45af53997c0cfd69ac178b69a38609fea79c9b30b99bd6a24fd33fe2e33c24ee85a6d70530a758b2be3d389e61d823662fe69dd966844782e6266a95a6d627283561271214d1e1fa894da2213b1b2f14ac4bbb13d9e9c353a1e238d50c26c01e90d77afcdb7447b174ecea077257be4e423ddf576c4c9306e1511a1d6a248975c5043f11cf31a7d7a340f68ee1f76f8f8bb32d705bd03b0794e42b98ae966aeebab2d86821419e9095ffc154d6d789cff6e09312193e97c1367e687a4b3583b031848236d9e2da4c1725850b369ec9b24e51080b79c1135b55ab81fb7b3498c33b468aa0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb53c749705196fbc7a5fe58d4568949f91ced9c88aa46bb0cc3fdf0a9bbe124e87e844fb8c716ba4ddbb3340932d34ce7f0e0fe0e7aff7e2889397d65b2371f23fb47ef20fe0ef521ab37c818078d137d5189f7d78080ebed045018197ce551aa6d8cddd5f60e540431254decc7e7dbcef9df4a1eea5c256cb2c2682d84ff08dac5b7b2a99f56b8b343c82096a14e0ad4e915374919dda05355b316da2331bb3f0d8363274c3ca4391b190dae6590613a59e29070f54a9f4de58ab1a8c4faaa88445682ae47270e0d9019b1e93f236ff55f960fe39d681c6f6a0f74a73d519c448b1e281c0eb2bbe283bd31a0d9735dd718f3fef9808adde5a44c79f0e511c8c941748c37fe403e64d4bde8c2cb0ccbb42b9d6a470610bf715560fad46757c931c912f40a528504fdf5068339d10f904e24e585d1d0a307fd57bced7a19b9cc8ca5fffb64b63f4bab9b18bcb12cdca84f37281b7058b802cb9d124ae145abcccd7e4a8b2f69491fb9ce8862c18a2d30fed7315b3e69f3af72f1985d3cbb14d078f5cc370a468a983afc987470d989a27ed8d1d23e1522df102cd73d0a5582481eacc6cb75edf2d4489f2db84cd91e9b680fee1c275545c2d89ddaebb1bdcfab01e4ce1d5ee460e3f5495ef50656f467c6a4d2186549bba0303a0bc6e04421305c65e855ef0a19ca697caef47d95d73be672797a49bc8478ba29f5618d45a59a4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he7cbdd938726a49faedc22e05ac617b3e84c9397fe2ea20c99d753a222b21e87e6334764151089e6e4ad930442af8c758ee8ed28749bb0bd25057f821608849c5643891f241d368c6b109c83afe3d1a24867b3640f72442bec9c1c9916de59123fcf79d481cbbf9f04de044e00d1cf6e28d47f131944d1b60ed64081013263b6baca7469e3f6fbc2f52c24de3ff934b40a5a35314da90e157d73d2e591614b965b77c77811d050822267782f65365736358b1c2e854f87f7f7b51afd637597d98edc48502f093a402ccf0aba1ff397a5e6912b858a6ac8234592031273e0f6ef04cbb8c41bc0613deeb2ddc19193d6922d1abba3638ce8d1d7432e18c6c7120e168250aa5a5c6df3411fb749fc0f574e032ee0a265a44335166ac75f0faf654f7fe537f3b6dd024572515b90dc8c0318bb010c5bd1b701c7e7a449a10df63649857ba72af825378acee10e8e8bb8511bc9dd7ece7a2fc927075420e7e39536a189c950a0760260e376ec5e602c6a3065b9f250f6e7a4f12b77d6d9e7ec57ad8a8a14a69793b248d5e59989ddec7700bd67244b3365b3e3e8db06cd18f29b03bf360ca545968987a247e95a1eebfba80d621bb6c6812d480228f8568790a5ffe2759531d6090f445e598e7e66ac33ce4f4f4ea7eac5c517e7ffd56f192ad36e24a67dd6676185c3420ae73e533ba010c8e81ac52571aeb017b8978e206c4d6f6d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8fe1aef1eff73e85f7f6e91b3b05ad04107d2a85d428ec5760bff7f73af19fae270e2efa5df890d53e96ebc6cb4c820b973f58758610a442dc3db37ad1bad52cebea5019bb374f0f1b9fe27a29bb22536cf2727528e294f144bed8b9984991b59ad109bc1f8a6d419275851d4ffb6c00f95f0b66990d9faa8d5877fe7459ee00807ef5180c5d80f9ce94679beb147e55e0c6fffba57f483a139b746fcc8dd265f22ff618629ae95d30ad2d609ca89aca3118427e13e662ab39bb05c4f3095655d525a5c4895d183683b9e0747eac78176fd7e6dcc0b0679cb572fc30732ee4c6f6a3a9d757fc6bd355e5912e95846938246c47eee765146a6f79063472604c8b06a420b9ce256f68fcb088d53099b160fd2156079bf4fa37b68e64f514b266624b215c07e356d6d00e6e1dbe2afb4d1955fb98b55676bb4c99dc43d079ea910b743da14c52bf4460008bdc5e6355912eca2ce3173e18592a81c5c8aa2d4cfacfce569da7592395411c29fd5626d5191829374c3f26d747f9ec269d1ff50ea5f9c5a810108493000aefd2eed04b7ce18b0f980dfa3d4b7e60b10033cbf74949a36765885d9e8acc8b7510c64e17e8a104d24c2206942cc01cb1af8b5ef6c881f65c5a6e5c6b6f07a0a8a8c7fcc67c0f1313d69990e3652b6c8b6c5a41674056c141bd35a7314a9e70d3a39b6416c4a636ce5269637e57ffde1a134ed3e4ba2a3a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h287cdfcb074ce0ee580c9c7bf9096d6c289f7dc0ab72117d0df0c1ffe8c6c45ae97eb67de8fbe89cbfdb8fa8f7e749983a623fe52e6fe16a1cf2fb2755717b9b0ae53d368d9b0abb5631169e480025be07800b8c67341721340d7027b5a834b5817a36dfa4ee4c57bb6b4630cc0b9385a2afb7be72c51db59719eee2739dbe3cee4c212aec8c45405ec21ef6693e29d04e5722433b65d6482821f1c3e98a7bcc1cc9b2dda040869aaf2e256b3af972ba4f5685c0e04aa7439677c8d03380aae7ee6b4a14e0a542efdf9308c78db9011d490e4de332c6053b72c8e0ff7cd5ada5696d54fcd5945f9e7efc0a9caa30682ebe2d8b96f7d2b5cef7d7d1eaf0645092d101c908fa323d3eff3cb4af045b411fe844d81681a60647b053838b443b00dca68b6725750509f8a288b467edbd625365b2daffc8ebc5239caac4763c5e482a2f498f020e174a5e4a97bebc33024b1b6767ff7fee466d4c1aa3067de12ecfe70b1418a7e998c4733826289af6df0aaf37fc35db28bae77f95bd88871739721cb5a94aca6ea9492d48ff2470d91b49c6f8f2c636e4b5af64da7e2d7510c8aaa5208fa2103ca065c7347f88fb23adf0e3343524ee7ca7d4f495af045ff296a9c0509e0015e4ebf29260c36542d68c44e9ce7ef41292525059ef879e16fb738d5b4bc8e2a9275c3b04c18d706235838874768b7d5164ef652834b0673ae852f359;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1ff07223781b714deba09802a19de2535554adb4addbb84c41a33dda703c54d688336d6de068db778420acf57fd97e16bb02f3b884d275e3dcb582001b37ba79228c490ee29cd925d8228059696b6504a86f8860bd1fa762d17d842b3ea3414f972946b49d5b61b73b523dca8a0b511ac79bdf929d8d08695dbe71f9aa04e1091d581aa3628ab0a81bcaff8f15cdf1c90e7fae437aebe9c51528143c1b61edcb62127d51b41d42520a45af722395e2de5fc0ba958b2761536ea690a2a3c35de6178adb3bb1c9994fe639f3fca2c920fd7e53e8a326e7bce492da0640deb21c33c5be9dd5bc077c26595793d7cc8b67f31d05844d4fafad257afa1d9ba0d4cdabe1ddbbfc05f6fc18bf7cf646a15fc2ed888eb0a2ac7556095ca8f393cf25571b79ef49439727058a54bb6954ee420f01d342e8d4538310d4f47b471e4950ae9d1be7f1b33159c035469e5cdab2823d50c1c6878520badb7270b532328050f30d2034c03dd76ee8129ef795f9bdbf5b1dc04770a98ce15624ec3399b66c6ad61d4f8b72e820f12cb8c4d20905fc6cd391b325163e9e635ba74a7761dc869886dd6a1c1863bd6ccc9fe42d54d7d32668a9d62845d211366d2ac9cf12adcdb5b1627b4b266ec6fd84e83d4784722928e14cbeb3b7ad5778ad6bc4ea3e8ba75211b8cc27839ca4b5d2bce6b75409d3914cb93e9eab0e8d03e6a21604f8bfb05f4f0f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h484c8a33317f4335107d5d88db7c7c7625b58b7d375a04ad10f06e968899940f45e88e7474f829f8c20291e04dda836349a46efb9bd223c18f4242c0b70f88b68ee4c26ed148de9da462ffe12324ca81d527b05736c0223baa7ce65ac4513ce4cb6ec4c8d3a9341b2c31b94eae0dd5b4a0341cb4152528a5e175bac2ed3a0370a27f27a4c1add8047ec099254924bef7267a590df8e3a70503371640ad758fca53a3d2d9a6a123913b5f4a0a5f1ab20864a740e0447f3662e5560a5da2c9ffe46b640ef71afbd0c6c509292297cf9d9689b9057bfbbf6d8df7d727b795ec55e2c446a6fb763cdc7c2a85057f0ad1bad9df8b0708c89e497695ae51e49c92bbaa613b4a2a68cf62e21c8029d7ecf408fd6cc2f999f4c5367e3f21ae98a3937628e1a5d5721a12e1c034ba974272b363e06b0a6c9ca92e4e96df84cdef36fd414c44673c777fdc5e1eac008c52587244f81beb60e2bae24d476ec62ac5009dbc1355359cfdee7e85102509122b12224e852a80e064572725ef7a8bb9a664a1912eecd35cd646fffd8e56845c56533c8e52375db93e17c325775419763d841d88fb14a2a668857c65217c6e9e7f1f037670437e5941cd860f8f69ddaf76c5998d117edf4ffef4222f2fbcd90ba9b3e271dd94cb384dbec783985c8be564db4024a7ea934b826e3421f84e3820d8ca942c29894c975d39b10247cc97bf7786c62c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h83f541199a014ecbc3fb12727bfda6173ae0a651b7b0e1e75115ceb2e4986978c95bf5ec8cc457326104bbb08d7e85482a4d02e4b00ede207908c245daf1c1ffe34d2f357174ad986137003cd9ca96b0d5a1c4563301e18617216cabe7b6083f4101af5e231d52c31612179f6b4f4e9d553aa07dd39da5b7e7c7a5a46b56e70cafd80b2d6d6e7f07c62f0bfbc9636e6e65117eacdc3c468453a584ba253d89ec221e835d21b0a5f0a2c359aa4eec9a8b69ee40fdaddf3f74500750defd773f2a0cde796da604b286153eea7e9d949b0feb4e916aa1a097f8cccbcde01dba3526726643596202fa9f182366e7507a018cb08ea212409223c187e9ea446e97b5613908009e5a160a65ce221511496266c9f0b5ae02d58edff77ea1d8f19d6e6117bc4ffa13fe82e8ce0c5f7971c3ca10cf443a9507c47faaf7770da476203e57dadd92160f71c54357665083c49a0280b3ea1f687be11313ca837c49048e670237d10e0d2aa5f5e6ab8a69782cd42a68a2f97cfa92e635e1879267057db9cacf3c608d4543b25320ac626ccb4bd8119d33af35d70b9c40ea48305c379718cc41d58c048a1cb2b9cc9f1f46c3919d24309ed0d60d655061a1cdff0f91ba35133a2d61a1b1828f8f954fd2c2d0d44ae8d9b08f5e99acb424af010d45a6b4c50a004614c8fea470cde8c4c656b2e1700630d65c63a89038c700e56e701932826dd68e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3f0d92ca7771ba9b71cb947fdd51f37ebc66944e9c5ef38af111b3f2bb5560c4e7c59548dc223dc9e352329f395d471e9aa7c931a1fb45b12d45bad9fa8e06dd76196be25f4c815d88e41266b3ccf90cd5cba2528321e2b536c8f265eb810fec084925eac68212eb29ce3dab6aa70ebf62907e96da4959b6c91cf7685cd01652b3c8ea72661f9535fb31f484a1add0d7f580621cfeb73493c61ec6f59bf34c9341c610492af2c2dd00fdd72ebec67893ae66a858a60598978ef584f168afafb86404281a01659cda2c99de1ee841f466068d96441e0e73a97fd43e768db6470c269d6be7f5e769f9bc34fea7fd2c89dd3c58637f155e1b1dc569daa14a521992edbecbd1ff97f633724f42151d3e3b2196df4d64d7a44db983a09b60ab06cc779fdd10ccd05f4de4dfb30721fa8fc2c68d545b120874b68865bfa0318b207bce931c8b8f68a91334e15ccb85098aef57f18522f992aa18c45019e8d01c63a99f610fdf4a2d47ee3a704a4ff5c7209dcb05ece368fdc8e878c84a29b6f707474fe777fa48e5fff4657279b7fbf5ff146661194f7ce9eae38ccdaaeb8db1b62b8f54f03c74990c326fed70a5f2c025062f6db2ccf0a942c27342a9fc75d8a95fb1fdd227934346ebf7a3e7c344347abadb443077a87a5919fb1d1729d0cad2ef9228af8d4ae954617838566b231b2343077d7eefd94ba0194a0b5d46edfc2a03e3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc7a95119b7a7c56ba33b3fe844e4ca22c4ffb0d2aa4fc95268b01d0672465c888d806a8fbbb5ee4e8349d297eb9aa10c4e93287b60a1a21dfa1c8080205cca871df3c8fe2c8f6beac6825c7924e57159bdb6ae00f4c77846e0d0ce044f181d538d3dcac1ab0c9566cc16d34967746fbb33d62f4027465f16308e1960fa736199a98619ca1e9c039bb14ac8624fac9f24f13f202e52d5e76d1bd49699a3e4ac553dd68bc4bcd9841065ab56117f0d5c7bb820438bfb40dd1121c13d0f594c0fa6e4254010debdaeb87ea88b027bc2482ff7345df45686fbcc7a4a1e47c0464fd4bd024cb5431472e12206503090c43bc24ec75a3cdb45071bb9460494f3a56de6528942651c75f65eaa87f5587a18e0fbaef0ea253aaeac1344f7634faa66efd8543877700e345dcaa26cc32429fa65bec5ba9adc550c1ee88316c840bcde2e960a6b024e96fdbdae8152ffdcd1f396dc4a7c2c6c736a3cd993c96ede5cecebc57643748991a76984852b84f52f56f5516a8024b38bf5a2d4ab4bdcaade9f30e9eafb095c32035e885c23b672d8d05944879eb658460f9b80cd3b2d83b7f36d08daddec2c6872658b1024b09c0c0f01adb8f87b20ea1c419560b7c0658dc02c3be1538434e678c0a5acd6128a7842db6ab3ccee5ac56e814642cbd1db022ba7f38754e963c94b4708c0f507ed7f1f0990b1f992551d491b32bdd394d0f2c8785;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc4472d95c65ebca792c69d0f58c2bd6d87820537e86843f7939fcd57e90f22f61a81bc512b0d4699c12d876f2b4c0327c85ec3568ac267ee631e2d3c24c84cf9d25c13120d43d44dc009bb145e9ae36953a45b53dae6a69cdeb94a38d09f01d4586947800313c0ebfc1164d20d5a778ab5e01901df5c19c68420dd29f55472c41286308f4b92ba1e4259a737683b8143b8c51c0e5b301d897454bc317cf23184a396f88ccac25a5c9f8631f06dcb41ce45e13e67f375c51db9af76e7ad19110469e99104c4e3c2c759c9bf9e9729d32e0925d4a26364c89a3cf4d043feecaa178f9c8dde6f9b4b2924411269ff0777b7ec69d97ee51ab2ff2d22d4b17bab84898e9f13605210f049642458135690250470b7b94f13d7e103596c5d584942e3a9ab863ce7858a810730c97d8b34132d63280c48be544bec70480d318911a3a4cf178179671ff0ae8c19c74dba6c1b83ca40b0748fcc3df4b3ec6da754612ba1dac87a97f7387c4f4eecdb4fd8fbadfbd7af6b7ac1ea677bfcdfba0664d613805fc249172ecfc42d71bed27d0a336c0f856aa74f8aa62eb169055dbdb8d4e61a5458a6ad4ef1d92f44b48d47e0d936781092435649ef66310a2064dbc54c5855225070c53bf388874c1e840d6ae537046b2d1f95e8046f98b0cf504fd57a7232f16b56ddcd1f00818cf977aee3a60893bc04733fcc8a0d5c853b870437f9992f74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2ea794fb734a22a2ef5042150bcfa19171552093bf7a83175594292cfc3c0339dfee7bbcd3a27e7a1d5ae119824871345b96813be5e0733b4dd8874944dc7402ea602a3308e4dae0601af353412c9d5bea1a0b8ad187d888173ab07463c8648d668b5664e4d7890f7e70e7347979fe83dd193caab6d64d56d21ac19b084f660dac2750431153d600810278e849bac262a62f999f24a819726ff2543cacb8b31f7c5acbcf2f5cf11d476e8d3311a073394ac98608dfa552509598021719b88a3f7e3c4e54b774370446c8cdf44917d843bca235c8b2db6b020ca7847d3768d28c281b580a3431db201db32ef8333d4f1cc6611203b9a11f02cbe4a552e0183fcf3674271d3ea68b73ac504f5d966e4781c4653e6b2ae8f01b7dc0d690eee2517f0b6e81cf3b5290dfc12ac1549b7eb0fc13bbe2d757097328da0ca206dbad11a34510deb6ea957de51c093b1f62eb545730c893b90ef3f8c48726f6f547fd811c8ea314d4e9d1685dba3f46dd2442f6495fca8b328189b811f271ccfdae16d887845765e36e44cfb20f75d8a36f44404d015930ebd7b948909fd77d77bbf9b876f80cae6744a51a69bd2538eec5eaa1dec33192de39e59ba973fbaee0e770335e14a2b4775ddf563e7b039c91224ad09486ce29d668f8a1a76ce87a75aea2d7912972e7fac79c30332e0745106f01bfbcef4d8aa802b9a6f14a19719ecdb1a12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h952a9b1f430faf41e3e95277498fc4f1e0b56dabd41de5d968896ce3144ad1aab741d282ec9c4e580bcadf3d5545dc77c3e43f9c11f9a7a0d6bac370ecc8e89e7684054e7fbcbc40fff8c04536653dfaeeb82f4061f632e79be3a3ca6c9edec758defeb659182f0172e5b47a405764ed5e9f314b3a9c1f01d81daa410e39e1a0cd474e04391272355012189638fde9090b52748269fa12627897fb9d4052a325c59edc1ca8d95e843ee859e61f0b77d6a62db4ac4872a287d74699bbe69f7a8c3b5ec7c6ae65c755dc056d722401fa9d035fbf0043933a35b2d04ca35db6de009c6dbbd1080e7f76b0c2222f55f0ff9f543251615f3aaf1a0b28d755a30f7be8a0915425a3e5ffc7fb805aa380d85c75f100777c96c268cfcd120f844098021e00fb22ac60756124bafe3285d25bbd8bbb0fb30e004676df0fae08bb207e198f5b51595e0974cd466255771c724baecb36a271696676ad393dccf7a8171a1edf8aee924caeb930292b2b8aa28db752ec8ff2aca50a21e49075239a7b879cc90fc64fdfbe7546761369bac3e792c01a9673c9c65f546971976198a9b120cd7ad6f57435b44a13ed5bbdcb5deb73d5c94b574928a78da3ea0e182ff21360e185ddb8f06623dc6f3fa622f87aa52be0a736cd80845b7f5d387d087539e1ff39711d0e9b476108a103aae1a0092080ca755742919bd043eb16abf9b7099b5190bc04;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he8931dd6465bc7818d8f6807574b607e984617fffad24ea3694b2534ffb6661500b30463ead9707790062fe97220c56b6339bfbda3958924d869f70273265574b704d2367a8e8c36ee7f00699c118d4580cdfcf4e5b4ca462d66d204c8ddd3daffe88f8b79ad3a53f622e60a746ff67acffa6def203bd3b06d649e7744a470ca5d61373ecb112baab50d287b5daa47498001c06297b372ce3bfa2cd46c531c10e19a18b572490a0785d845e03664cf795e0889e057ea49841425a07fe0515cfc4cb5aa524483f6e5cf1fbc3eaa11900545fe300262c5182fbe408843132e21da55cec15e80995db7a840a2b7de549112db6697bd647f96aca16bdd243713cfdc3dc71d34e19fb7e1172c5816a0a4d5e7d00d1eec5cad7f2ec045770461eac9aa299306dd7c3407db4589c1934ac59cecaa12c7d3aec21de0a5b9a7211153cbd236a05f8651d0e7d2c808b875512e7f1c7c73e62e84be425586220cffb51ea69966f9e1517c0103e3e3bd0028491568854e772ce87761d1331f9d2464b245e41bce3494c3d420ae54968fd67a082fe7a8bfdb5bdf5a99d8a90cb6765d9731ad40fa048e9a637b88fcf6251075fdc7189a0cd4e4742d9b8ad5f9aae6451b16e66801f88e1c64a147923ccc5a0993537bf38d4443f52c1d5acd595ca6c677cba5d1e43fe64c4146876d68e81c3542ad8862fc698c244852a7611352408971815c42;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h26485f910f244d7176df4494113042e15430bc45fefa1b76bd34dd53b75b606fef4a07bb1a9e33200745a2871e70086838ef5fe7d1a34da76273b25d8dda45e20b0d2262eceb6712e18c6de39f5f1a027954bec629dab1b40d527ab7315af605fb3cfed8976b9602a15fd56251c09b4184bebb918b294b2f830180ea11bf9e4ff1ed2e30b7b6e34cf884b7bb799ab9aa1fd41f18edca4de1d1e0952beb093c552c6ae5c2ce22ae040f772c8fa8860b74bd76f9d3f0620eff0499523882a116a2fa51fdb1d396df84d306fa33150f765f9b33037aeb93e1f8fd68c49ac3aa2d1fad01a0d969d5e2acb6e09f03f3ec124d28167a7ec38fb1f5b1f07fa84a937f27eb025cf29a56d9b184ecef071ffd6b47599e988395da4690d87fd8f36ccf3b281aa26d2f2e1f39776ed2df6c10c1710e69a83730b63ad0321e1a7bbc730f590ac2e1b1fe8575dce66b7aaa7d26299017428b7e631c4dd07f5075dc97633eb80abb4d02d65e95c5f0c4a32dd888972b95faf6a728f7924cbaa0c66495fdcd9929479c85f3822dd0e211e1f8726b0e5dbdcf4ba2bfb984d8d70e76e584d4538535c7b233f36c1d3c70574f24096fd339c144470230ccab80af7fce7a8e432430cb66a9eb173ecd41b5659b70c75d7121e12a8b475a3aec612eeb0b7853c5835f70d834bb968ab0e91e5d03b564dfb56eab35cfcad4541bf6e38a334b25cc23274;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hce4c68dc27922fdb26c691cc369df1b40769be9361e1bb08ad98b5dd1e169a163be718a2b0b34adc50d0af23f6ff93ab67465739e6e284057cc5bced4b47c69484be352af0c2cab6a37fccbada8da26a6fdb2633e74cc7a931f676fed4cf16b028b94e6f66b6169530801f568b7e68f01753a6fdc0a352ed6e0d37ace753d23546c45a08c8429b83a95197ef4fbce838a6cdf43b7ecce1c1c8d1f016a84dfb0f66da612c15a1cc123c11269186c8540494ebb3825197b1852c80c94c749dedcda87346748a6d7eff92367f7b72380d399098c0d12b9135fdfdd670dad59a4851f129e599950f137f399a05f1d0108e7999528702b24bf79b08d3d164634d1dd14a6bcc2978855d918cd4b1b20fd52ca4244c3e680bed170105277d89f119aa1fda4575d0cd2c03880aeae2706b120e64aa8db1bf4835d19c98fbe59f665ee37386cc610b8ce7da36b4c8c7f6f81fa4dfc7d5db536a7892794929a2faa34143fb76afad86e21d1d0ce06be4473e1b348633d6c813acdc89a65c51feff85ae2d64d00c1ec4a15039ec36336b3cc742c95c231b43c4aa5368cb0d404db6d96c0982b43d8566b5f8f06e2e8d069041a05530c01198e4a2cf593ab25f7945f87ed1cba49d9a7be870172517dfc14613c0a0ed99ad0bd58e12f057efbfe0403725a740e42bcda52f4ddf8aa00b890451bf66ad17ecde235c5b2972277dccc40dfef2b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e15dee49cab7cf699d07cea2155c7a81a54a03abda121e4eb561b8557883d3fd12b13455fb11f1becc72da4d3a52b34eb596a34ce96b914812415883647fc70c187331a788d1bcaa36adffb4eb579b3cbc87fb62340a391933ed0a0da44ce504c97066eb71ddf5e8a4b27c1d1c71d01a0531a99fdcf31b71855ce3ef1aa474267353de3de8de587b796019e6c42fa344167f3d833906377246212bbe8a3d0345949d285fdf2a181d8607b3d7b9f9af5087ce88811d468926ac2eaa7d4364efef00c2cf26dd977387b19ade266eaffda247d20f5921090b41859fac40c2781210ad243f8804732dff213a4cff088fa1734521cd3c2ca25119f76d1d4a2acdb54f2bea3545bfed98be1add8a4fa85f875b5034c17ab93c77287da33d298735eae5382a55709431965a2b29de8513849627b38ffc68737a529e779a41b62d90999acea1a82523ccb9ea6ee2c20047c5ce3fb7079787d755113a9fb1ee8b611b644bb9cf746a73022c0617917486aeaad35fda3bee904bc5f22910261b8406427db3eb472f2c5124be2ea5ad86cc3a50e940727bbddb15c12cbde3d4d49a4f9796484b45d3fe83f2e72c711dff2408d04f6d3184cf03b22243627e60a13b72cb3d5ced882a05e7c4ae9a393ed987d9d027df552bf2041bf9365ddc8ba8293523be5a947b2c2bca8425abe3108740f2fbceaee82e62f351ac52e4580057e9621f400;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8d5e144fb5d3cd79e8307b8b234434772a9b9b854ec248ce67c67a44ad88b7d2ebe7d8d86112dc0201a431e36cb68b541f78e6fdeb293049493966e2d74c30db03d15218a270a10e3e47035c4814f5eba0334cc58d5826172dca5c18d1beb4e30ac3b9012266250d99038cccb0dbfb3194e9f2f40edd1a92036f9f88d03909a45f38e4e2d1d23fb6fb68184e015bcfd1bed4e3da9fc6483ea2ab0df576c5f0c2611e9952793d0ff68ba2d8f194820a5faafd694d7c4e2c5d773c05ca4d2df2d9c09c6988aa9dd27bee7a114288c8a671531cf93c392c21d06d64d20103711f2171d3fe09e061f5509e7c6dbe2c0d93de0ab34223356f47000bbbad39f7011295071bd1264712a6358bc53f9268124cd28349b3316e449803f8db69b3a729c98bc9d509f1b108c146f4cffb68b39b7cc6c5747b2abccd2939be46142e349148832a9ff6dffae4cfb393a628544c3f66f95814198b9a2103022f985320be00ec6301f24af19ebfd99d570ab9011e9b7e6f314311aee10061198abbddb96bef9f5657e2ff2ef7911d435180a652873b9598ba57bc4efd8a348ce88bb171260d78a690978de38955d013c51d4991e38d438d448997bebc5316b3b18e9be7d431be6655bc700eb7f06bb582e195a5707c1073341c9305107b3f95f0c804b0184f9e3d75b5964f62548f33660e218807c5512b112727a806b13d46b103921fba9c03d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc91bc6c9ce7298d30d1c374abe65ec42c3c37b55fd3a68fa6bc5e1cbe7970e36e6785f2499e560ec95f30f2b299b61148dc633efa02d022c9c29f2049b4cc574ac59436d839e551d51483f969951f66fa0183dc152fe2ceda6cbcb4efd7a9af3ce2deac72d3cb882ea19345588bf7d15c13828ef5373b2b180f129c04baf793bd33d03d507b3fe0ee4b0daf6ec93177b017983ac92ca0c78f699c809e3209599a205d7ed6f42e107d01ac0ce7794a78a96a23280a69ae0533ee52c4a6923f3b91ac37861682bcf2ea802e4433b7e635e8d6f614f7908ae76bd0d8d49c786f7e7c8c259efdedad2d0a787b3d688b252dcf7ff448e5c0e63519a129b2aeefc2101ec341ae95a1cf579e12da595a7c04d54eb558b4d12e32cb7cc00f405fa4e3ae7b5e94de414316c35fe168407552a4fce95429d6292816ea58c0c394a57efba9222950cb7809cdee84d00e023454faa065722a7bcfdfafc7fc245693ef407f9a8ad382f5330aad5387c535af5ce9db57d95102d8a6c23ded66bfae614fd65d074b53dfb897ff983bafb86234d9238694ab4ea4b0c9d897c9a7638a8ee86b631293fbe266c65e3b1058d39e77bbbb9aefaa91a837762b330912781effe91c4344475c5e2cfe02fe58f1f5d304cfcc1f258c23355774a9f0d52e08de98cd66cac532e498a2e47cc03fa1fe4d6c23b60b975be06a7c5ac03a22c816894f050524f02;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h644a7212a12289fc63a253137b4a9b43041f63c432dd909d090f8455430783ed1fe4b4828c18584d82cfb4ab08205b6b1f86e1b26c08f8a028472bc39ac36a3708fd690cb2a62d643b95ed2c7d4d86eb693c378a12ec62b6cf3d1027ed7dec38ce86fe6ad52db81521af75700f24e179d53b2f85fc2f9046149ce2d40d6b9cae40aef6ab441673110712597d72453df535accea9573ca4efcf79817c0f9e594bad584d8557e39172a6bd28624d2e5b595d2c4d042066ceaabcfbba75fc43334e6f3d4bae8a752b85c7ecfd286ddb03f81eab5705ff57609f0453af9ef1f46270f10232791c7fb2c0af6c0a119b852c1dc9e311809f6275247db4477296b329237c19e5233cba14337eec9a28e4e2b9f741f775b315d8d2ebd48300d29a93b501871b00d8916fffa0d51b01011ff5a2185c877349943739be7c74495688980f25375991ab87baf5a61a096829a7bf0cb092ced42448ce6cd17e9980c241a6baa0f6e4d3b3270617f1298dd75e0093ef92547541042e6b99aac5ab95a0bd1232b3e91c19ca42f6684d7717e434ce86dc534fbc70af469d071bf891a4b7d18fce7c199a0807461d10b4ae42ccda2fb41d8b9bd7a028ec747d5f6b3ced5d3abaacb9d5b3eaac4fe14d27875cc38cf80062249332e4c021c2b17253e66e7f0fbf4f8070316eeeb990142016d44650ab7ecd9a75ba5bb5ffde535509287c4479e9453f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h487c74c400ca0b1282da6b097f96702c9ef722e876112fd9daf34be62e69b517c955ca5bf327a3dc59e811a293118d372b944be6aad7402bc26e50aadf5a53bc2a795f15170da3a9eb9a53970247b61c01692751bcdfe52484cbdafe5913c796209feff5aa5e171bb8a3125e059535363535e5973cbb8b2b99a8f74c6b79b460e5fa7f332eccedb4acf322da9e3d7fb4254dfa0941cf302b9ec6ee6900d83c4fc9fbbf99e0b5c85e3bd5aa25fb1e4de426241e2fe739e888af8f8f6dc413c7aa71933da52babf8b0a94843bdc4f884dbecabbcafa2f867f26f26d7f805cac83797da04261507f6f0504410a6ba2055908ffcb94ac875432698b380785b0c4cad1c03fc215bb9a26fe77af2dda4b5d5665fb347103408ed11f1833f056d2853148cb68981d96b87893d8ddab7ab74c6392b8aad00edef4bd3c07eb48edcc9dffdff9e7f81023daeb2fbad83084e7709046f4ac3074574a41f336d29442b3b7980e56641f56ce4b7af2ac01d3dda75b991183ffc3dd335a3462ed6c0eb9fc20eb548a9b131be8345672f3632aeac5b3f06509140f2d73363f26b0412e962ee302b67c1e1e25d87558f961c7699a935cfcc149e6e33c979200b589e9d5169f3cc6bc091c0cc8510daee476df17df2df0e82a180475407497fbab4f5387edeac576a1d8094633beec315165db3050bfc9edecb773cb9e06a8f5ca2412bc948ffee71;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd73c3dd225952e72675b9813c8fa8b8b91e9642e43afa7c23539e638e5cac452f32170e08dce5c3ab4499b0346f0ea61435a5e37cfd4bdba10e2d683bbc5e99e9ceb5b7149ece9fef2aaf56bdf37a34a0fa47d50c3808b1aeb3de6755b1403c57445760566413f0ff28bbd18ee892aa25ef985068d830b49373a5cdda8620deae873c0eb0dc0476cd0862141cd4dcdc18167f6d3dd2bc4a53187b779db8a5f2d770d7558405de1c982df0e76418b0698c9e147649377692f28cf69989d67b1664b5fe573a3f0038ddc52e3e327f74713a33b575ff3edbfce14a649d9f2f911674f30b46fc7a0a02828988c5f191abacd0ff4e9a1c4e5f38dc70d8cd5f4d88988f5bac5e1ff31a1fcee246a662b3de6beaeb8c745fd0b39906abc543bdde7f60d04461509abef954f84fd50111a080ad54193c9777840424fea24923865eff1fdb98edb9e13125304a384bc0567b9de193e4c0b9d715896e38ff2bb85f24a0811eef06fc4e3b41a044d5e0989f7e58d4ab499aa8110f419b241bf09fbb1b8e3d80b42126fdafc01f32246b8dae762722dcf677be692bef00a6552fe2d982b0cdc98636ea7109db6d7946cca2c6f66c9160a37a1f59866cdb2cdd3efaefa553327824936d1fc2a9eef69eebfa4c59bcfb7d37cc188bdd3db71afb3ca4a9986dcb845e742b48f405c933130eeb9b9739542411e0e94261cc4a9dd89c555ab096b78;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3bb77bac1c51743936a9fccb1e0b25a8feadfd88231165040cffc4428fc09b440036518eaf8b1710e9409edb0e714920b568182d8a6482f575b7226a15bca0d767c07bf0a8a454935d49bada76379b5de64db03e78d922b3c35be9ded8089807a559aaa0da3d6f0b883c49c4aba297f9ad4070b46cd338d67cc59143a0043d7984f7871184a2cba2d84a418ac29e653ae73b4d8c3dc2e5e736a82351c5ac3c65a1af2058e134e0abc6b83a79d320072b697dd6bd42bfc491b1bdd99def62c8d0071f53eb171ee6f5717230b68e833430b9098a7116a508304dbef22b5f13503e5bdf1d314fd589802f03b52d0f258d34f6ac8b887833901a80dc7e0aad40a98133b3b3a7466572003427884bd13c5a7b7a42138a2f8b833a3d7a83799bb26265eda83e3ee5c1ef410f518f8339439fb2feb5de4704187736bd5f1587a991bd015e003dc3ded6523d045815748545e270687d0231f7b91335f650f1e842df36dfd220e4011637ca98ef5b04b65b8aa91eba3e607fe7988a9b2b4a7937c52328a2293a6922a827411ab0d71dcc690a1c7284c4913d8dbacb1817467afae1237fa87f80706404e0c6deb60da720a175a8b3f340519b712ea1ebcc83ffe9d2a8521c44e52cec6acd9ebd46b62d0223c488c83fce20fa9c8c5c636d92fd8880c7c10e0e40fa9f6fb8c3c835058aa91e0181c50e862543bc4ee0d6a35aa4f075e58388;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h424b2d249288cc45873e42b76f261fe44e192aae85cab6b9c9412fa75a8c3ac850ac215bf236dd1f91729fdb606a99120755554b67a2bcce72d63666000db367c930608ff3c1fd2fc0108fef8de64d23f9a7f3c0f2578a0fbc99f732bd9a57629dc0a3eb59edb4412d51c50f81e782942a46af397d02c71f6d5c51a89a0ab247beac1d891bd9a9840a46c4fa7ff3356405290b55ded9d318e0adb6d9cf2bf37fa6debf5e55f5c082c1e66ee8b309371e4e4525f97d35e7caf64e84901acb047dd631948285f72f9e20a0cb7e72dd746d779091f002b65f6b1e1c429381002512f406ea2b8e48938c73bdf420a63401cf5d4bf789bcf5977145964c85e76edcdc8836003dbf15fdfbad040fbd9b0ca05a426d5c39c32162b3fbe2ac0f4c2032ef420c636f04dc92de72a31558ed9e0b6c2a9dbdab3ce88b42877e1ea8e4ea70640caf8c87940760f17b2c51ae62bcc749e598c99f7e79404d54560a27a7bc936f23e30eff2713ba85806fd09319d9b6e549d09a1a6592960fc6eeae172a2256378624878fb51057d5c96c7480d4b7ab7981cd1076450e59feabc1c5f1c72a152c7c75ca7fc2051ccecef4d6b40d78bdf69703ae089c2f30979789cedd45229b2bf64044a201effbc707103b9a96296edbfef365fc85a7b89a5fcea42dc898e4fcadf7799b5539206e2d211a3ad4d7eb016e11cad75ee2e08dde14906cf56b1058;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha3d37973e478747e33aeeb2f1cd594dcd159a2b84fb8aaa0b4e0d3b181c41a299d7fbc35897e78647a174330b0c4e4c1c0b092739194db9e75b2931e39ab4e314951a7e744278087bd09de975dca77a7b7eeaecd4dc701558fcf13a51bfcf3f1597d4af9d479c117444c8f2e661b52bd6a7b626e1a8ada15f8ba87b2aedbff9e5eaecf10436d0e094b4c51f846855fc64c8846ff6f53cb904cf033e17cf8e49409b52f5ec4de953fc6b6d387b700222788b4f098ea2ddff1a678d8745e418eab7919503813f240f1444cc5f9be6b7bcb64f2c78e0fc8804fbbd62f18c203409986007d6df4b53434d4db6293a70f46b5f93efb892be1197263c17f239dc617ae051afd0a73c89c957f2e77542868d8ca167ae7eb13554c0439477a24a846b8ba88c7dfac37535ebe698189c21216409ce625a10035123ecbb698ec14eb9c383eb620b0e85dec3e287629c544326f9e0dfd96376333f95f55154c5960ae02899c97a480a12bacd1d3ea9c2aebadc35583e999a100d60db7cb1df62e6a9c6c168a9be87cdf57edd6911bb710c4188411d52726ca677202b193a9ff75c94f2f0fa1b9f4d614450a9312f61f9621b7161aafbb9ffee063b04f348bdc7e630eaf08ae39799bfb88145e5e3400069a4964e67b1c19f5b0a4bec002ef49cc57b4aaa0a062b01f6a7a865769c2967c2907f9e2547ccb56fe5c859ec05cd090ad7b294ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffaae5fcddac941ae01587bfb11cab4bb299f120138809aae82113c1b9d90bb99458a9059163cbed6acdfef12784b021f5fb75b79ff096d94443e54091e83b5842a61b797d94daa2ec557c7a82c56a933fa29430e3be2f9e8c184b8e81a9b8b1707d7dd1e0a2c568857df832df2c214600e8048d19f3aa781002c71809d4f258e767ac92f8f131108e9c2e195006887db62141ea4535359cc8c8240b1171a5ba6ac49b5fe96c985280ead592ddf094d302eb3d2d085ff24c42a0c1d802415464fc6550aa0e9753c901a38cc30fef2bcbc2cb4c840859467cc90d843284f2096a5865aaf2e58570e31f57df6897f3dd7e4d8df6b58d1e2f28c6f2f233f7f1df4472bb42d3139179ee0e4e91a2c84903e8f7902e2a7703c9ad4ee0f166b0b2ba0036aa64f64cbeba4dfba29d33f172e7d5b25317ece5470ab733ac2c00211b8608bcf223984596efb2d0f70685450cb0080ca58d845f4d981b92973eb7e4f3b78ea4eee053fc2745440356efa5236e322cf136e8473a1f1788bf0192831f383cae30da4ce693d1d28126c1a25e21c91eee2a673e46b9ab8462108e7684675834d19593228b29513b7e03354a15f890da373fb1b473f58f4fe22b0aa96affdb4a62545c7fcec341af0bf69ec45b6ef8adbb724376a4d6ddf4716ea8ccc37e4b3c37bc80a3e864413eb6b91ac6201688829832b553ab4828af1f0296f18e2cac0eb9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h75bb8df2ae259d95f878207635e51dd5efeace4c347fa435967f139bd2d7158324ae20d2d90063065dcdaa6c264eb9e7d13bf98a734bf478c3a7597e78e2c4ce234f20b2810be109ddc2488b31b2a09f2dd9cc9f62f6d12b636a17abded43f8fab762b70ac2056e5ae2038a5d81c6886d97058d63d02c955abdbb781cdb15af4bdfebd165751a7d7f2b5d528f36c4ed6f07f13ea181c468aceb1f51bb47b58da81a120fbf36ca91880337b0bc9ffb82a90ccd228083997f5b533ebf6d3b85a3c64bafab5c59e8f779ea60ee549b9e820b628159363fb29ea9781a4b06dad90ef7677070d69ab666ac3c68807ea5084e4fda87dff06a3f27a1c14c29b67cc7d3c3a7b7ba9b98cc45c17055bed66bc199a3fdb37aa90ccf5f73a1cc74e3d8186ee7d63769e566ed1ec548cefd3ba20be60d7b1022dae665c3ed772f461b1c7ca6784787f139bb7a465eeaf1de264b004a97f61edb82938f26eaea9e051f1b3cbf4c35cd9a11161bee460357e1a09e725dd5ce9fd28f2d1a673c418211aeb29f627f4aaf999372776c4858fc46f9f0b2edcb5c6f769cab2c74f0c9360c1139bacdd3ebc7f88f3b0db7306915ec40b90d18a044524fd000988b39ed07e03b3d62bdcf33675c5e3699de01c622a77e256cde581b1bf2786edd45fa1343252f543bdb973038f6d787cbb64b25ac29af5eaa2166b2a9b4eac94dc4a2aa002902e6b9b74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14a4c58171ade1fb97349aa94ec89bda6d73718fb3146d68b6cf1d24f2adf00915ae7779adc275f7ec9f826b1820bb7d367d2de9925bb2e912cbac0256b6bfc55988c00c12e88297cf98cd5284c4d03f7b41b6320a48d386bbdfb54cb7ba3d42a80904ec0ccb10cfb3de548820a3047805bcffc02dde0dfedd3d89ff8458528a26d67e137388e90db2e6350835da3a2ace4203aaa4f61f46573d5294dff6840d810eccc03d73426a61165bb418421bad6d73924754ccfeaf8f0876967aed0ea42fa9275caab213aa3f5b5be8d3a22d364df71dc988e4f217aaa76fb43109dbc7f75660f18f8f0fdcf7d543cc870544100da6e6df4106420d858c17d66f5be9400759f3db1a26d6a2504edb9505201cef02c91182c5ca39d2fca13dea4f9e49f1f1153c4389da234ca2f834e4c3fe395eb56193cf44aa1409f610826f2c56a69457e13a658785a356c8e9493e90a85ea86155427de412249a32f058c04ead73a9077b4dd6361c7cc0ae02bc4f69c4c9a1aa615e7420ef471efb4c254451f436e65f49a395407444265be82fa773bbac123bab67d87670605cf0f46396c7c9510878a8975957a2bb1b092392adb58642760d0a4848d259b133015a2b6b4638f3658f1c720d4faa1cb5977292a8f4f2e5ec0d2d71e43554adeba874fc2035dd045ddc793681843003641d49fc41faeae92e90092efcbacfe0246cbf68a3eea3412f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb2e859fa669792185a21fe52d73c4b597ac19e2d39740be777d1c72a7aa688416b3ed52db9f48e8c861883115e4542c73d564c1d5cf45c432435746cf87da09e0734e354a43014914722ef15fccad1954fd7e7d7567e8de96e26458b224db2ae4b6c91107b45e9459e7185fab5249d0513554f7c628ad99ef3206def388cef1dcbf9f7f56a64d0aa817394915c60f6b92416bdf641ab3d43624c18df8afd28611cb79872ae922fbd5b4e716ac48afd6d173aa963705df70c00ef39fbbdbc4df9049ae84960784df9780133e9100943f66158bef5ca9b1a3802d0adc336b9be5aa35869a2ff0133a860ca485828cfcfd78c0a5d736fa8b30ade36a2e101736fd1c3a449428a5361180e48f7f81ba21388243145fae3187714e514b523e7a1591e80118a71c9b9af536b2632ae37f888736c8801c8cbaceecf4fe50ec3071c7719636febf140415ee4621734fd0ed0a69d6d3eb53873219c172977fb6b7076649c33e8c031ceb8ce1ef4691c4692a562a345ed53a7ed6372d4d3e1d8654499c40cbd0007aae5f7c346f845449958de736d410ede163a23e29386511368b87b49635acb3953c246511faeee980afccefd53eae52dc9517d3779921180e31bc0ea9020bba19eb8104addaaa53899163e0460a66053da25fe56818e38bb96109e6a55c1857ab7f3608f9b05207133fc07601548a7f44a6cf4fa4e6518456817c729d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha42eda6fbe37bdd4370efc519011f2a9ddcd49672d4343926709b065f0fb6f284477da01bae645fb56da74ec9b70cd9846dad878acba08a1b0df953455347cf6da54415f3c1a3bf64ab7096c5fba66b897493abf23cf6b0025c378d3049c645aa49a8ec34768b1ef4fbb45274462787b43d4b5447bba9fa4b998ac87ff8e24a723a7a803daa4ed8ec9d3eb88a56985e388923e6e975f4c0f8bd5bc0e30800507949a9912fc581b9558449c6a98b52e40ddf32d65ff732f477c7006378344dff7d552148d203c11e15788a78cb0a08531c7f07bb0211a0b9c33b1bac65b6391f661644323b5dbf217de0bcfa7862c54c52e928a0417daa7a2d03ed55a37303fae307d9e6cec5f3b3211e0066f885e26f7687316a4ab4947acb517697143f470a9a0464afa87ff2f875de9eda997ad590e9939dfe7e5526113bbec1a6ebd6c706d878e45faf6f3e6130ff85e82da2b2aa477a317326897ada58523c0a3d9a96ef0bfcbf094036c63e2ca35e7cb6f79203cfe1804217b01a4a8a9200015348b87ea1d0928aa4c81508451c9d7990dad225fe4235da0e07798d6625e6e5e6051caf50f16ced060fa78c0da019108d5d9429c21078bc18405b0e0709fa2ccd6d68698eeaceeb81d5aa5ecc9f9d22e4297185799589045be11f76006e1c12702370be835df3e7ab58066bb23a6904f7690a1c49f7cddaec661e9f5d703ff7fd816ca0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4c3a1e96254227ad92d17498293bcb5f7f7176a7621a257d30e44670fd8b3d4d3e54017a60a7f77c384fc7d72fb0ecb86f71c01b51d5b59bdde53b62309e34ea01faf046decb20db6f6717ddfc659a87c64c53af287ebe631010c4d020c8a0aa46e8bc69e80545f9c42c3ddf9b5e63625f46874cd2bec567af5a3ddf6e8cd0cf834b3072456ff97acefa578fa66841b42bc65abd6ba117100de9a8c63c9575c0c9175caefb49087ab0d42f2cc1a083a63d409c74ae6ecf4fc57c12514b89c7165d2ae5f3c8c6312dc1cc1362c47e07fca800b5c7ea178e473bb71b42b211cbebadb7083e93d3f36fc5798f083d35655ae6467e1c72191d603ca67bc591375624f8d8a130b3aaf23fe169fc211f7aa2ac2510894b4e6e040c9808b92ed500d532d06ed44f71795b1941bb1791865b5925aac3fc687ed080ca475ac7e59b017a98d9974782d320ceb4cd79b9a772b017f18d52c2c448da082a8cc614adf3db8a45291516fed3da274be352c44b7ce6bc298a76745f789c34c573fa39bd0ca98c40660b6b309948992d83e1564a4b55fdea863e9aad65acaf9ef74a7506eb8749cea9538ef730632bcaba9175a968f1c54f2186c07c5b0b08144c2be05a5c2a51d1b19d26f729707905ff34c71254f5edb06db64bf4aff116290b0a1b845cb5ca00c52c95e08ec7468086be05b27d55ed4b3e9848de5b8d62e0c3349332198e11c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdb2dbc7600885045f1d799155df848379894bd78fdf6f5d684d1a686add6203013f070d2da8f2943c94fd644dba3f8a15013dbe5326607346ff51c054cb1eca8e21620071790c4baeb03451bb78ea3e610a6fc5b311f25d2c1e15d2e61d199a27964820e64a04d57c9dfd9dd2eb147db5383a6c13e54231627082f519be612c655e648ad729d561575e22736e59db629f5f5c8b91391204a55218fbc7846e8b64ad759a56667cc6e21f8afe8534c908053645abf6f52aedd626bc89c82552400d56693d1bba6a91aa36d481eba347aee52eb1b36e9c1e473c33f36989afbbbd7c38143f66c5b1564debf958f5645de09518bd71b0fe17c13a47743bbf67051d65cb4c341ae134a6df40196ee1d45fe288ab302007132a5e81fc3ba38db985876bf98d892eea94f4e13c3b057710b001cdff3a799c2558959dfd7ccdd3d0af1d4781174da31453a3cd91b217148c57ea7369886c23bddad6ac1d01e3db4ee1464d6b5560b3957fc603b1b7b56875b12a91ed19f13f21947a10f38a2cab2de8e14ac4ae3ef1c6b8d9cd38c2115015c25fbafa253c858faecf001e38f17f02dd24b92183b7dbe55b3010148210a765c29bb783a1d37caa259bd6a79a9089a3e659137b71fa56d3b93c8f34f77718f8e2895182d045f32eefea2df04647dc813cb72575564df742a22087959c667d7d380d245ef6314e92163f8541483b715cb0f63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14d26617d6444a86097cbe0b28ebc28b9e32ce46ea5f261b67a90e05a8b8bbc852c83628981aec540ac472ca08dedfba5b05a84ac57e5b36a4d68f030e8f5d53850d87de1ab8d47617551e044367f683c5b637b6dbee9aca10674618bbea9aa4f94652d6e189194a64a8f7768b1a3a11b95687986d374fd0db3fbb538dc02401b2fc68e46fd3fdae1c4858887e5855df1c493929adbd0005501368ad0af893c79e6be9b31f571e20ccfdf4794e02e59a76d32f4218531a7542c8f6bf26b9fddd2be2aa32aa34ad32a53a0015dea7e9f8d694aa1ec6ce891a1129e9f77701e18304c2c259ca04980a7f251317df3416dfdb6f9dcbf968ed579f95d31a753bbc56de06634e7ce9e2e0b86eaf858378374c39a3b1fd1a8e58d779d6091c2e80847f1cbf1d6f6f770f19c7d25df3adec1126921f8bfdae6183a94d911c6110d8a589c47d9a0969bd604d92be9acb73936d9cee539436cb0f81a2d37bf53c7a3c35430a8f8b9ea7dd6e61ff186a3fccdfd7bc984689f2ea8665e6e3ae903d8f6068727c134c594ef134741b873b7f78393126b696042366d77a36c0d925392ef55ad7d1cf149b6465fe637dcc9f922f09512c6aaff7d41925edbaa2edad324e99250cddbed125eab633d62d1ea8a371ed8c752aa113e9fe2c444415d8c23378504f6b1c1c368c1bfef2bbf4d67b1bed650d845d24659611edc4d23205d74106540a1e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb160caffa9bad60ca14dac51efa4f1b8d93435952f2f3ea39561a7b7cb3b7cce40015efe074d993fa7bee0ec0f011afaedb6c9f585e2e40484a03da814d004d8ca0d9b722a32e5d7a808d49d26d57be80423ca1041b4acb10ebf50e8c9f8cc04063833fff3c35bac3c4d60f82a995d7bd9ea2d9783d756e0687a997f04917e87729f208c069865408dcfc090ebd519b2a7b0daeadb17f6f1894ea67f7fb79c3579716311adf8234d3c37ea0ca6f63401026bfc8c07bf23da69bb900c10b4784d4e77cec7810989f70406ded1797e83168522e624299f59483625a652eecdcfe55e266954c2c96fe37bf83041790eaca16a6d1e5ecc28de2e40bad4e10e1e85130d9a1526b6b35a4dc9cd112795096d37ddd3814d96e676f8420318b152cd9165048a6aa80b4d9d4e0fd29267aa4a964553d090f09c1f179e67ed27926665a25ec863fbef89d4e9141a6594a816de6df1d92061f65f276eafea888f0d420c18310fca8546157351caf65bae1859678eededbcbc772e6a4e17d3ef34e8d04d757738ae923a354ef9294ec0a8c5809f5896ae35d301e793838d8555f399047cfd068c42a91ae14f4b4f0d3b73ffce0e7bd454da343ec0ad900436ff8b95d2760bfea2546c8d1f839dff6e2a40621fac88fd1a12e3b6103ecd49f6e0d99ab539218d40c0767e4194d01a0cd9ac04d595ce696f93f8b2ae6a9749c8d2ebd25f36b450;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3bae231b23cd4d1a42ec8a1e1ea0029f2e0168257416b75c250fddb116c12f1a34b264ce22ee31983280777ad417a5a80face049a90b6fea72b36227ea30b31c94fdd38d3580a22294eb7083f7b0997be8f60eb43d7d030aa3d885ffc3b8c6f608871ea38529601c88ea45917b561b27ea431024b9cb37d59ad6a77586a8452ea47abecdf072d2b8d845a716367bfd4eafbd940370b28700894a739868319cd7e092b46ace2ba9c503b4fd6ebd34f6487f2431c7997578413ac5db91db784f27ce33e9c7773538068fdc79ae44c9b47192c9be4bb84b2e104caebd5a7836ff340ab188bd18800487236aabace42171d10aa2f64d7de62a4d96c1a19317bc456adeec622e41929e893a5cb6ffd4c8189b429ec389a1179220f414b6aa28ccdb07eca7c21bb5944818ba6882d78dbbaadf5a5b483511863f0b8906f70c30508e61c5cf8a9e882b7c492094401e16ecb1d4356111a7fc444a8109b492dffa2fdb257cbf422fe3d1cf9a8546de40581488bbe7336b4ecf49643fb994b199584eec5c69545c8392d9b0fcfb1a8a50fbbf4b0cd658c6857bc75cfb12b0a21e80e9cb3da001c8476619be850a1af358129dacb55578ba0636f5e9a1ac72a56a871c3d2fe4e3ad0705ce5b26410026eabcc74ee03363f6730b4360bc603e18621783fb48b3f45ea17ad90d32e9750110c7fb17e24c898024438c945571ad8d7885ab98c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4daa44bd4cdc51d84e0feb50acf5e6531c618fb2d4013126b3f12473ba6fc1e1b3c2053a760bfd3dd0b7870bd6a649e9713e85a58b2fd2aa6db353fb8c4ef7d2e6654fc7dfbda84e39088e6e876984bb12038abe57553b8535d3fda032b9c4cffe44f9e0418cf02635a8fb5c987ccd8bd186c62953978da44dc10b132237e76b1110fa39be57a58f42ed3ba92d4fa06a530c64b81bace7419ca930f44eaecc32030e541daec3aa65674fe25ff2c291abcdeaee57fd41ddd7f50a546fe7a7166128d1382cb19b9b6b65752342c927dad409ba98da011d889f15fe45472da4020024003c7983815926db4ba489634b3d8d3c3399fc0d59a16139d0fade5fcc36ca7a61de5a855f530da30dd399bcd8f5e327f42f4556d642a649502118dfa8be94881dd0c9cc65093919a0469eaa048ebc601f6bce2605937f44e4fa00f5f245c82faf6357de51d3442725c8dd7c99661d406b6263202e8d59ce2a737ed5c0f88e39d312d44aaa25cae0d11339d1f465b73644b9614f45c70bcac391b0233e94329a85dea3342ec037fdf8841a0ddf9d8b20d1c2e002238c2473fe3b0c5f32dfc7399ad2459fadcf1691296c26dca2e5c719e6dc94304f44c8164cf64057db7b17405e0e8d6a0c7989849097ad45871c0a847c684d7eb2a869384bb2f48d202f698dfa67273f8c8deccdf77636bc0a831716d209be052bd46ea27d28661dd1338;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h76909467498511197af0a603109b18cdfdb390f5a245416a0bc128727fa915ae677c4e87a56a4af11a804fa6091b735da294529579bdf81b9a83b0885ad65a6223af19d356e324118f1222696dfc80be8320faa7c4a1fd9aebff4e3757d966a46f9f9dbc646a70345a6552b3e69a23c8c3aa3dcd003b4ed48f6bf8e09c77511edec9bdf79d85d97915bc3495bc094e16ec6f85385e08cc440c0e13ad07c0ad95ab5d03e0fe846db1cf0bcd9e9429c77b6075519b708f7c46157d452c7c690d0917f82ef0a6acd575d3c027da2659e2df29ef696fbd90a631169fffb32d7c5382d1eaeb32609172681686a3219ccd9fc9ffc2cb09ce8281dcd16e35a1ecff6a627d03c66077a1462086b2586a8bd2775d075110596aaf2500c1a2f3900ba288ea9c6b686f576b6ea6813880793fe0cf3cd24d5c8b4af9f2f0b4c2e914fd9397dddf49de57c97718deb18dda6da4696d333ae7d9b965a2f5873636c49c38dec3938cc61f9b6c5cd6cfe5700f80bafe5506ac8e9857fc537763ae6e07a36533f6b967b824a89e4669d278095e362f01e5c9e8eb58c4ae5a438d540aef407cfb4fd3346962ece243934efb71392ea91ae2f5ff9c40f18d1baef705d22318e390dc6c3ee77cc9f91a4977ee4c94680d0e3073902f80f4da7dd930260f034b4802108165fef1bc41fd1ebb455c600848fe08d442643ec8c364cbb1582374ebc4e7d49b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb76e29869f950f6af33903494344f0842dca965519f5f9a2cf752321edf8f98f45281b29dbd89cca99d819cc3fa46ee928e886794ae2186d57c0799b3a6192fc25fa37a4f3dacb0c1ade4c9af77dc2050278dd50c0fad298444359b465dfe9444bdd5a81ce3dba954dd3db56b20c5d103de050631e5d3862a92d5f2903762eec5257c7605cbad63c0ccab2dde383159c4eb82a98cc52752e6003d6f9a900822e13d961511e7a94158ffa50c12210518eecca075237f4798cfa9771c885037eb7007e885d49e92a4291ddda4a37b279b90d2f4a6c515c96e45ecf0649ef42e985b9f155b83812610ba4b6632c5c60350edc5b383368e3e6472ba159c7b1c4b1202b767c334a95b9136e3bb89a8122334f0364b9287552862bd0a44ed213c284880cde0a960a166d1a45271d7710b030aff9c14185e56166563b0f99d6b2b0b14328032ccd9d7bb0ed000df8af4d1cb8bbba36295c6015aec999121eed6071053337dadf2e0248cfe157ad9df038b947b98a27f18fd6634fd1d854fecbcf7d099a31907f7cf422ce19539e671cadb9f95a78164ded18bf9dc6aa8ae9390108fdb27b20872de8d0071b0518f7dbb62f0eb2ccb51e9f05ccf7fd157c264f83e31942e7783ede56d7300f856cd00445c0a4121b198f36124516d11c0c2ea165925cb6d0533bdfe12f0d2d42735485a9b16febb8d0b8da2c71307ace172fd5ed35c383;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h846d1bae0b37ff4c360274f89ac7c4edb796cc2eef6793cf60570a0297ee2e20238d525f1679d671916afc1b70223dd9eeeb3e4754a8b0aa86116321c209c6b44fd40b46404060b494ceabc8d87cba17497218aa70eff8dee9e805d4553022aa7ba5215827a3c70955cbdb9c8e08834c43c31707d198db9ad3c4fb4218c4524cef624dbc406359683dbe9b989eced1de08ab627e5945df1aa7790049fa79435fba2d2c9e02ef718f1b731d1be1f203b6fdb06132ac50606f6f91f15e2c932bb3357e17578ff7893d44b09554af8e923b9cc8f2487902188b3beb5a8da1a16515010d26a636e96f3e384764b2311997cfeaaeb1888d49dd441e2730eb9247e9962d45d739b6fd64f903251558bb85c4c1a203efcdf087f61f3ca149d5f681f74c85f82212b76afb55e8010d38631a80865fa36e53fa67d40dcb44b5536fd92d3954b00289c0743cc75a6ac316303f8eb1bb772c585a4fcf671573e473ff84f6a90498942f9eb2c95e35d3e5b18609cda83939f218b18ec3584a4ef9eae3b4da4e4d1516b3c99395cd07061cddc66627836b68d90fca47e2c237d491fffc923c5b863426da0e468904f8f3937fec7d313544ddb8b365c63feec5b993f35d0961ff6dd98eb38c149ca8c2fc227d2a1bd813cf0694c053735db189ee9c6fafd78dc7be72564d940c2f4b00e03bc4e76a86169db833e126dec182db7a7bca2e254b75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8e9b9aa1af35b0d3e4aec56593601c347a8c102ad4addad74a7381b6060762a326a0b727a5ae33efd86d106cc8834ea9bf257ccf3a33f0d5b9f1f65ee0361dff6deb0ff22465b07b2317477f7f6f5eeb008cecb46493dbea6a320ea07709c7207252037e3b22ece2b87f3565ac2b7c172ae72563839cdb64fc56a53bdd8d38663d975ec1bfca360fa6585016daa137b7d26706c16db793e9a20eab89559ee69590a1fab334650fc931393dff577ad0b3e08c67aca03fe02750b8e3cdda9dcf1806bfdd97b2d4d7f06d94cca65ab39083f8cc32ef328c474d7a24210431a17d113f61423bf74dfabacb7f49fdebe6d965aecfab70b21f5c22d67c78b726bc6a46cc3a680cceada091781c24723e14e514ba2edde9f2c66580f71658de7c088c3ee049546bcdf8a7685356c202bbd6b510e96bddad599d364dbb4bce9b74baa4bb3f1cec4225f770b9aaf28e1129c999ad0acdf8e0bd634c58b889a1258ffb713d4c04b2be3bb2b789820813e39e90845694bc1d4d6fc92bb43f9fc182a1800141d339d1acdec9c466fa85e1d1f2db2553d16dfa8cc95b617d266d202f0757273ddd651f0f52e51404095a54f1521d5b7f1b85dcb3d1ed68e9c0880edb491cdb4546ed164d6cd7e10cf44cc0011ca4bd9fa567015c62ee73f5eae7ee2a8e1f077cff58352891443a92228e3f1b2762a7d992402dd6a23cd0afa1c8445deff0e5bf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h29eb81d6102678c3d20773769fd6263b8ff61514709e38501fa4ce8073eea442bf21454fc1f9c5e6385ff9ebc57a96618d118be7895c0a7c64f26d5e76cab47f1b0b2b9ce2ad742efa0c5eff6153ff572736ea9162e655e30005b40e98d41987e4e0ee783d3b9a6946b28f40ba69f34e286e80012a6e538151234353d91504194f29083b17f7e492dd75b13b47eec26e3a8a766b2cf7987b26073e5759b09952faebaddc319817b875c9b9776c231381c33b8feabf491bba4cb0aac67266d817bedc16cbb96b693af65d8b26dbfed416ac8bcd190e25f51162ce09a510e5290be04bf99033e10b650bd0fb64dd363fb7883d5adc2529ab6e8fe144be666a6d45fce7d79e8f2c7dc61420a5e5a57b93d0aa43d8bca54f5f80e71c8364bb8cb3340d045b81f18397926c412fccfbdba52ca8122e468846ed890f77cd8c8b6d8bc44067c1d8a99731ff556a4a838126bc164885fcab71b51cb8aa0b5545c08374fb33e25805fb436584cc44bb391591afa462d53cc82b494e53b73515acbd72f3328e92e438ca3671cb218216b792688ea4d95a5dfe0d10bb03f02cdd4f2f4d8a37ba1a0f685f5133258f26830b66ae4ddcaa74ebe8e2de3f07162cb0019a7a0cee2f8d91f249abc0afd1165b643fab1b7627b87d2c8aca21ee51662e67bedf965fce0274a8d0a37afd640a62c0f04dda5ecffa61000a59356e1013d4c5bb883305;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h46f682ffa48ae397dbcb9e9cf2c950fbd79d62bdcf37fcc27b84fcd0f75f20c758be5ae71602b77ed7d1fc3e3c86529b26b4b6f7b4fd6fe7d01e6e7b557b722c7caf8ba5241e161c4ce7fbe886e0416ef4c64f384bb49c617e93407bda47711c13a0c42149bccf5a216d0a7c15a82fead9ceefa3f4d691ebece14489cc77feb974c646d50a0fcf608085d3b44fd8bfd212b20e4dcb0737eef34609977f71657c8ae1b83ed443f0e690b589d3ccc27655b434b2bd1948121aa3db7dd63695b317efc972d82f103d70fc35a0bc5e05222b841cdb73b417e98e87204b1731f357482b1685a0d0d8fa81f79012609c7fe5445b7c6ac10643889789367802ea529eb4e0afffb8b097462c9072920c19b8d9cfa02ba016b91d891c69a14703f3330c93586c59e3dd1a598945f1a7888fe040c3f48dfa6acb708ee995a28bc7473718212ac193efd7e33a627c29bb5fdf0dffc709bf3f9771e277f9e7d16bd0ebd5a4790da4553d4f1989419c1bc090551094d561e332166430df2958308a958f2df4805ae93f5952f3ce415f6801267cf01a8a9bb524a5218357b1f9a14abfde83284eb352ab78c62591a2b4cb40da1d8c4b54344ab5b528002934130f6034b59916c4a1174bb7057673c8876c676c808304cbc2159bbb15c65c23ddd05c62f83415378115d1e56d74b84984058f30769c67db95681a5369fc0bcb6890723bea460b86;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3460d142993b6f7bad9b3108f4a99dbeb977341724edbe7d83660606facec3846e6aa427a1ac9dfd7d9e2078fd1b1f67dfe23382e2b974d9c36621f91ea14a3fd4a2b6ee840b5ea98e80c71efcd926edad313b435c1f2fb40b04637b3ce2c7e5170d1e0707d54aeeee7b24b280a8e015096ec68fc857522f78e85cb9e311d6162fa6fe0a5cb214733991055de12de92b35a7810ca6d5164792629cb843286b1f84588f33834b912a56ab5f279a60b040294c8166c484f279cfa99cf67dd71852ee147cbe54cec1e1d6c8d9c36dfdf2dd3f5269974262b3e95163dc916d4f34abba29ec160b74de47eaa942549339eff850bd9c3e1d25bef23f894cbd1d543c77f5a50025b1e112329ff61b8eba7bda6397716f472aa3a8f5928da6994715b28adaec73591190888d71a4f794e2529415ee79980d20676a0d63c1564cbf8186de3bb2f41d2044e66d8a5bed2ea15034e4e0f60d94f5997e7a8f7df8d9956e11fa4357d9c072b7cd640b014d955b1e53c27244008bfaa285986308e1e24814456c50289d9b96900c205ac3896af368cbf5a5b57cffef0ede8ee1fde73a5cd7a851ed379b79dc1c3a4d9d5ee9c6832d603aed166d8a77103278928e7231cef8a986e2e5c601b08b5827345aafab6facee3cc9a3ee085489137425eb679328a3c54167d0dc67c12462a5a6a7628a4e12eb1027c903f61e3696daabaa55a64b36955b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h140b1dc720a343880805cc5840f081921063fdd125fc7f13286f91c0f0c12261685bafa9878e5539fa0635a69b5d2a24e1fb620e45914b61250ffe8a35735839fa8a570aa04a6283fcbcf7c92afd11ad7d06f8c75586bf78026705b1d5a95c3b3d14d8922efb58e4b338125d7c23e6b3987faecc4b00fe5c7cd105ca320cfc9ba658ce587df76e5ed86a7e8d34c0dc16796f4d8c3c1e92e8cd8b64110c3a388211c97ab99b2a20040f9d85045afd176b96296aeb33a8c83b31e5e3d2d2c3cee321faa6e8d587ca58b4c302cffe3ac7c933df70d343d9978eb91ff201e047726b1344c6435ae13992078099ba2b2e2b5dbbb04fd3497c80ecd188e4747ea05f237c0ac8c57f8d0f2c4e8f798d4e9da69f68d106f728ecd64d2f5e4757458666ef1ed18d6dc29445b651a664961d69d018bc2a679d5ee2a9111d15fe53fd9ae3a95fab362919b6fed2cbc5debbadecfc2a0c4ecef6a60588fc441786b57d1358c5f76dc13bc12aecf5bddec570f5c720f166fd2300a4a86eeb51e1706f3ba3a9663b009b682a9622648684ae2ef7f7eff374ae7f1229c04489778a8e2f00235d41f1ff3ec97092bebf9fc597d0e2cfbfe91b58c281825b02c265cead5287d8fef579cf44b68bd0157c13d3c9bc39cc6730b2fdb1d1f4af9afdcc82adb05a365372cb5c85ef99c7bc966bffad51b521f007793c89eca61b7bd2b4e9fbf8c3e8e13c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5dbcb4e7ab0bb4582427575890b5844dd6222ca5b97e4e679c3005be7b1185972848b8fe36d847140bd04ac22f8eccad6d6c6c6240b7b0d4fe50d83d13978542c8de01eb13a9c2e81ea1503e1eaf493400460085001865d58d7798993d1c2959b473ccfc15fda28958075c60f80b0f8a8fb48019ae03ff7539a9daf93640a4e34d9e19eb71a0906ccc537cde56317929eef3a8a7de91960fe4d819e95982c8927363882aaf1325086bb60f5a513a2878a8b05f4fc60af184b1bb092fea7350ee65adfb29a95ad7f0020bd6317a254fa998c07fb1684045a329f6e2972a56b63ac7a4de3909ff63fed04705d321b2bea1fbf54c0b64dc43d08ab8eb3c34b4759840f2ca6054820645dcc4c5cf1654992f35f4a74bcc97978f9f8cf07a26eb9462eda16b77e2709963725ba831c8fa9fda88d813014a831d91adf3efdd1ac9c2bf57749c267218e6941cd3c4fc7f9a13c858898dbdec09681db1c4c102968d7275b0eb895152d97e35850b1493b9d53d6ec5e675bf975b8d665327daf72ae32e915f60e16da4331e7f306cff8e6cc1a1e046694632f3768dab920e3f2b2d49b78f422a57ba968c65172c083ebc7d61224f978cee11557bd747e655db7093fb1cf741e1abc59349cc10cfde6811d6e06746e48c071b817ef9c3b105a7f1448b1dfc23abe22ba3dbadaa301d80a3e11d2c199c0dcf69425382f401938d3c6cf5a309;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd69360a7fbad7d82be6ec37996019f3b2c826e3b0c94d2cddaf8f049edf347cd82a8ab2d493fe41ce3656f0af8b33bb19ad39976ba0f4435be325904f09dc5e80198067317be46e16c7f19bb5e53082a0e5ab75fad276427a2c8f1bdb19de031267f0c2b73f123b8ccf50840fb1e59356c2f12e3a87340cf7e8c8308c916687959f17cdb79ba570148f3a2c262028ea34dd332c9584bfbe85ec3a1b9a43e7699b0d6344b3c829172fdd5ba5b1a1a8bc845e39cd3bfef282164ef17d2eff0a480b6f69b76d89c49076e986c050b1a0a999064b0e797b792b5aa14e742d5b9ea4fbb222d7e1873c22f207d7873fab25882cf4643cc98d9a5ade8cb9005cd98a73173acebc2c0375546a76773075bb5366bd32524d7576c25ebd66b31bdf0d342acf2f81f64298706260ecf967a5f258731fbc6606fd1b7e79d9781ddc47fd9546e15b7607d3d4cd355e5acc048a24a692976f96fbd90b6fc79de1c9c052e6ccbda358a4a72dba930a9713b3fdf3096934de7d300a908a2a5562559bb1acfdb8760eedd44e717f75282acaf55a98679a49311f6da7cb9cf057e5ac0ba21a1eebaeca0566de861dbe36cadc06c70b7d8b56a7e5040060f89f30b6e4e313469fede2326ca33800b7123f1c2c7bc03da920b8509e3ae704cdbe1681c80b370e27906d328313074370d07bf63a1ce3a2c1cd8109eb03e6dd3952900af4ee24626af4ad7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5c914eaf049ca90ab5d84f0e6f55da559fe7ddf8864a2b4278c490f6dce000096e74442844f21cf30c19abdcd21e1976a7ffc02f238a3c388b5811ac57bcad30730c4bcc2027a46b14149723a777ada0dfdd68ee1452e36b3d4940537ea261645ee3ae748ab46021c4ac3874e04df7b490bd876170a507a14542346fd7215184f67cbd49f7ddcdfaf3142704bb2577569d187aad9a936772a322e5a6041f1ae7b62f8a825b9aeb30324ef96a58ce2559021d51eb52c528b87cb5d2217eb012e4a8af3c4aaf27449e35bb2f02145dd0fa98a3d38caf87271bb674f65a8b9b0c3402101ab03608443e893dd2478f23bb2371395a068bf67816d8699bc4fd1b183c74deadf87b75fba279b8e4cd9d93905438c1c3b6692bebdda9ef6b654663a1e2269a755fc66eb6dac902497b2b88b0c5356a74cb6ce5a3e55e9d8a4fb68d4780b7adaac2d4ec50d8113cd1ca1eec8d0aca2a7773da8a954b5ffe8a771d792c074b27ad8564082b3d7cbf46e87c9c6eb83df016b03b2079cebc4345bd7af0248f077b6e5ecde6fb9e40108af7d7a9dd0d5896c69aefd1686c074133a2b786a213f9f8387036890c54c2e306eec571e0e0d426ff08f7e9146226edd7abcdcaeedaef46df446d7e9a469afd8b5280a6d5627c33349feb632e8b83da9458fba9b5300298653dc7beed20d837bae2d0bd8802e5834b0fd501c813245c079de54b4e00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8aaf7149a375d85336a4b8b77b7d6f54ca506c05dc903ed1daabec6fa74b9f662a96e152187ce4ab7b7354077d033c26c7964b32eb1385ca66599312c6a2702e2508d36d31ecb918aa405f0b0e2209e4ce8ef37cda6d30b6649b132b1bb07957ec5c4fb072587d3b9f8168ab320330bc802483919d47ba832e5343e70cf4eadc96773c6b22e33da3d872e2927bd2d8ac31c6e51aab05956d059463a9d69c6639b1407e3087b90b16b761f031e7d39373a2377ec8f35d7ad84c2b1d3af23051027ad03415fd7212e1034ba8e0d37c18c87311398c65426d11f766b648d6b47f5dbc6bbef86167b978086e1eca6cd3a21ac56c0424c190d2053ce10df90b0dcabbda662c5ce4cfb7e351da9f527105a3ad12654cb87e0a5f4a05e0cf5c9e51e1402cc7a3850054ad5b3c73ca161622e505fa4399e8b24c743c70c9e9440429e424d4169f916acee77bb134401767a6309b40c4b28027ac40a3828871caa72dce8b4a6c8003b1540f08ed607e7a3cf533d7f5f3bbaf4f46df6ccb9617445b0769579fd0bf6a40ff6d50e6daf01fe0da03a78ef51258b89ef902f245eea3686578a892b94fcbf21e785e5234f83d1bd2f7b542b37e4fed68b3a2debdff76c02cad4c413abc1b3fb48fdaf5e60dd47379fec86f44ac0c04419bfe6d364088c6e322ad8e50efa9d19153f911becdec2beb59ddb29dd0f96b5dc1ef2244f21b3c336f87;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8e7b4a829fdca14c747cc2651edb89ee90e6d508fe61fd927cbd638e83ded4a6b79ad9acf26dc065b243670294bf3ff120714965b77f3921887cfabe795cf45bb469c0c8be2e571cbd9a779c2d715bb35ce36a07890d26898e78a0eea1187ec25d5b82ddaed3620a479921b72a290e0f66471ec6cb7a9897e57c57926a0b009eb61618beae5a6e0109ba4713657643957ed3bcd1340cc16875e8fe7901dceee3943cc0f0616590c15582cee4b7f321b0d7f48a74156ad0f17cb1f724cc8fb10ceef66088bfbdf95872d39cb5c0360e32b829096025e990ca6f4f655a97c25d9f1d9e494bc5afc1e130ec001a4b99cd58d7e719b77c198b47cbf2a54c892cfd587ee6199107732634ba234fe6c0afe552be495fe57192a4e71b5fab975fd5d24a1614c115f1fc00907264bb7fde53cbeb4c1531bc414b0997709b4ea42be680e3406991a9063dabe7536df491ffe3ebaeab35bc4bd7104402d9c411a6ff4c947e2fe58efc90c4b963537363ac0ac2174c1b61161912c920126f81f7c7ff3f7c3ee8cfb376ba80eaab2a0056a3cf267bc4d4e211c05498744e6aa75f2c87b7eef0c2bbc3d17001bb97f5c5b568cf0a5fd78d12297de5574b1532907dcc7a1dc82c5a799dd8c9a7210e1c9260803f4ef49d486a8064feb4ff662fa0bfffe47e1349b4f693aa2c08287b4d006bbcae249ba9a84fde8ffef8464eac102ac05cca8360;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'had19593e6a53f38a370ed87b175d9760df37258d92849daae18a8426cd0586a0654e8cb990a9806495bdab95cef142165e766a8c6e326ceb00a584b2c0a1a1cd1cde0d624f87a1d089eb48f31d3644cbc84d8660ca0c60e06870713f7aa93f556f8354a877ba88c57d14f89d9dbbfed6490aa7cb01b4a346e58f36f91ecb2480f11c6e7bca5b49ae6da4d0a134270c33f4ee6a2ab264c6aff151c0646330e27665948ca384845a9a29cc563b6bb81ab4d8dff873d9945608c420365cbfcced7eafac21a817db189120d46b6f95bade9552037e5259e93ff72a23958efd8a816f2bf00d05d897d66bb8f557bef3c44ac69505bf14c2f070ebb5d4ae913f75c14b6265cb34e7b57e0a2a134d494ae24e3803540e08f468271364608f5d30d5b2af6d92ad5e17ccd2c4097578e3fcbdd2b5d419fa92056bbf63772f8ede0d5d03a1ae41bbb902f8f42b86524b87aec1e2bf521b5d84e3d2915b27f688387c6da8a0a3940e72fecabf9f8da830f408b933131e1563d8043c65148b3ab7bad68d8f3e88947070cb1ad1fb402ecf1e48a48908df8f7a73bfaf525a5c8350ecc89b8431413d50ad1bd503d8ba3e725d40144761530823ff9c6a109963c559e03f1f163cacaf9d4183a5619dfa3b098339827febe1205c6bf303246034220866c7ee881271296c517d0a271bfa11e2cbfefeaf3bc6e17c2afa64603c71d1d4bef1a2272f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7e24d3d68eb391d1d42304f113ff19fa63d5bcac9acc0487b2a0497041aa9adc406a60efc753e746e00a7f9afd50a255413551f7e9a3791867281715670259ca64097e1fb320820d91edd5e9e7a585e2be34a10392d1d7ac32930cad027b5c3740982b7ebaeb01db1abd6950a9ca790efbecae5d060516a865de6bdd2308e56e0a5ef57028633ac03bf2591b0a34e04d49b205ed2410dde2a70ddd73e31d3c0f2a32d42ca178dd05449f3a02f9a13c376544429f7c85147ce550e6205436bb4227e46ec61d30d6a13e270315187e128ed61c4a1177fb302cbd3aeb2a22178aca80ab7bc72ad00db99738fdd9c6c9f8708ab525478444023fca3aa218e3623e1b0ecefca650d1fa64c77bf84e5d28972dd1214d28088ee855da1a114b51f7b8cb5489e436c4e3ce01f5a7571a1a119a08403c95a54072f2f26f017374b8cfc081bf32aa9bc1944d8b1402e10f642108f0d4b874996a793ad3b83f53212a0eeda0d8bd523bfbdbbc7ee594df84a0564ba1553cf35f8282838b2da20ca46bf6012f28879cbc837f1652e53e2c7d11d8606d512905ff9b1c2678b1ec15fc4488e51c449f23a4c6dc6c5f9d8be1a1dafd28c354ca184ebfe240cfeb5c20bdf0d1fb61961fe1aaf2a21f1ce0907aef128258930aba32c604e73e7fb5f29d136c206e1aa96aebd79bdaf5440c8100ac867f93872851add20b8e8f0ae60fee19e07d4711;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbef32514bffc7551b04b0d4e8c80c81ef4a4e724835fab0a27828c20b3e728c77cc38afccf1837221860f47b78b25abf4e4700fe2b17be4bdacc8315cb68a7f72b9ac26ea86791d5ca9b16183b61c60c16cc9970f16f28aab07d516df65133bd1ab0cda8a83c6c22424434332594ae88a9cd78799e3c9de8ed1cacaf71cda25f492082c981df49905bccf6424a8116a5171ea222b9e192626897162a89f797c45c218dc2dc931ce35d641545aa9522a8fb5fa7122b638628d1d1c7919486b3257e7ec2e73f86d8fc7fd4689dbf0376b07e2daad3d3c9d2fb5f03eb94e5c2caba253c7273ab86b95849c0485e47d0b0b59c0eead32704b1c2d90c0956911dcda5b069bb0f3934b21d89c47150beb84376ea6b3da492b96915d72f080e792fe5a4c5f7b07a5568c8c58dec80277bb1f28645e2e4370740e365fb2423a467cbe2b16a3298b9d0098fe50383bc2c0a49c035eeb81951a1150f98637e008114fc271f307198e8c5e31673359c0f16607e87b6c6d5086aa87eb48367dac151d5af4f98e33001dcbaed280a9c414701f510d2d15655e057357030cdcbe1a6902579bec67fe764f5e228288a3049cb8190e374ab34de178a45262212ef5579a6611a1e25956a64d2421984e6bdc5cb20e3cc6afcdfe1cfbf635ccb4bc6ff2eb65f4a18fdcec07315b90a78a7a102dc419407d4c553a6d7e1324572a13ece925aa30159ed;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h826a39e136a8af8cd0d61064adb7c9a4f5828ba8ffbb41559dfed9b173df5e9402d81a12aa73b4b81bce2d728dbacef6ed95990ee617f4093b0d75034c2dbdced11cda90713bedc2274fca722a8162a6584b700394bcdca770676c95c62571405ee391f866f912f663c9ebaba3c64ed5477e4375488f357f79650105263e4b61564ff52b4c8ecefb598dbc313b5378d10ce588ecff4d619170066abc52e7f9a8df229bd0d26c87c92f28878350d11de6771296e80542adfdbf3a50bf5ec70f70d066155989a701818687f7bc5ba46ca708c8e0de16391337851a834792487dd01bc0a6b47c0f85738eeac6c7272ba01e5729253211d35883cb38667feeb216a1ad534383931929a17b7cb09b29145783761e6be9812a0aa2aa96e571db72f01729e61aa6c2b42a3b9ea48e499c4fc4aeb6323c238722e932c2e31b297bdcfd64ccb65dd059c7cd4619a9eb2e6c8afd313013db7f42df38bc9dc05c0886f5e7b3cb5fad7de01dbd4a4af0e4a9013d2731540c7b59e8add0044b9cb4bc8b5e88fcd880f913e228eb7fe4d462fae21eeb07fc9b2008ed3dd807e3a1b5f798a3a04283e1de9ce7cfb5c89c537438f58df489f93b2acf0ea0723e0c4df1da1fcca6da4825e732215c532bd9bd48ec5b88465c84536d03087d2eddb31c3d6862c9f43b0cad5b8ce1e7040f8df1b25e0bf5998671c69461e1a6bc01724586ff0e7ddb9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb72a339958985d78225c780e9a52a868de09fb114fac15f327e04d10004283110b2f142f0e4f5e5db58442d05f63498d5442e037e9b693f1fd3a4117ce2f139512d2deb31757449da59d999c86fa4025b38c51f5515c3f842a3b64456f15b104c9f128f2bfb09480280124115e87b85f70051bca70e55a86134d96c7e98e280fe3730a328a06467c2179a9f222337cfbe52b13a3674303ee96b064ce4b71656bc29c0fcab76c27fc19492bca1a5c1dcfed7005d9579cd2b06ab14dc5686af9ec065933c23ca736f6a9130a989403a35dda2988380a0289a3344fa7a8f6517a6fbe91706cea891251ba0053224b1178ad7ae3ecc635f0fe374da38796a4bd36bd386fc0498cff8d52b3042fe0cd216fa92afcc152c286f9d52d1e0616900cf2f59d3706054f67d495aedb675829884fa9e1a6c388a7fc43c821a08ce2b9bae4eb747a5669b8af2836ed8aaa94053fbf60744a22467f8cf59e3ee29ae443f2cce3ddfa122cb80317ae2789b0de43d5fed8dbb6f4800fc89835e644d7455944ebb2735d6f5c1a7a0ae5198ef6d31c7a696dc2c89bbb061b598cc25051acae12ac0ef0de8bad39d4cabf11bd6aad32fef0b9e3bcf591b61faceeffe3f8862a1c110694d7a5b43657b394eb75a43f7df977dfe27288bb4e593cc676605100403f2145e859a4024fb658461d38043c7399dd75c841b6751205aa53e27b8c16a806c292;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7ef2618abc1bdbd1feb43821a6d79e606545d8a97600002abf1ce60fc59b7058648e98ed216bb33574740e05e6f306d8edef93617424cf845c21e7aa896b9f1bf0df5fcec3476070003342c1a5a0416bf79be1be95668dc63477b43c5c8e85bb08d09de1d67219462f45a8727e2eda61fdbbf07003b7f386f0e2e21314faa5a7b72e1acd48df2a9a52d00a47d670721b07c31fd54c993fb5c0c6e39a81df5830b0d2a1e3231c2e654a7d2bd303a086942de1d814d75a38bab14dab785c8d8887c0bff357cb0dcee4c838abba3743a25564a0534dbe0eabf2bc3ff17bdbc394e273ac89334535eb11776ef667dccded86a746b1d060134a6664c4c30a581f73d43199c6950fde68c19fd8ff371e6ee89b21d12515e48715fa6227b705263f597e6c5be7c0bad6406536283a5fce5fc5fa39616c8b8936e522d112f55204fb71c6435d57f6fc694dbd8b193730c82be2b217799e4bc0a0b838ade19ab98c508c2c0b2d6070cbda128b5844f4818f2ab821eb383c1afeeffa9b585f7bf8fbc76f4d258653c158eef1eb8c5e59579d0c9c63fd644bd5772ba698893fcfb7c50498dfd53d4ce15ca97ebc15379b5d010653210e6d26729e8777fa27314c5d43093ee2bc41a929c3bfd42df137ea2f4cef12884418229817f1d0189ead45106ffd20fec2c73c77298a0794a8b4ad72b10cae208a25cb43ffd5a666b237f32c19078d2f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4f85bd08b32f8d1c88fd0d48f83951a7d06bf2002163157fae07516b80e1d2f986486cdc5fe64507051ac8e341b4e43e3206d5999d20f533c896fc099a48f28a69ffe062b72261d96820b8629ec8460be7ca4006adcb39542d4ac7f459dc3229491f611eb2185597eea29d62969024278859ca2dc1c7a3ac3ef12e6e37535085de59b0a78a4d73699c1de5c862a15dd970cf8b2447e2296bb0f437855d3ad58bf4dee58c2c5f7a425d7870279937b13ec02da2476b6d7641e0a821578770af4e2b738a3ef5ca66787f00eef64df3a6185f6ce5205a2f4404540d2cbf9f29ef0ef8ed562531e629a6d8ad20cd1fe5bfc441d1a78c84261249906afb96f5a5ba6a705141aedcf321dd4665f7e39b9b2f73bcddd6a94f659f9327c3f12e1fa12a90ad6a5c2ebec853a5bc875b9177258e8a207b48ea1b7d3aa65596de58100da2d7cc921c043c9ce81a37a87148f6e4db488597d8e779a6ea11dab1b10e2c31785149ab458ec8d86b88b9b330804197e2d607c90e741fe442a22449bc488c5a7b2e0fdd0f55a038be40bc252d93aae3d9b9d4a7aa3a40b3de04b127db844699df87b17962d9413bf60577a9f02d279e6175641b738110379242309f037320e2d47a9c06c1e075a0824f75fd48491dcf1e00bacb1ae499c14844ad6a475417f679bfc72c3a8207a12bcc841f3a2932241a0e3c91b30e4b1e50f6111ff468c90da348;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he9a947739add3bc05987e4cfa8288f54aa9c45a333e5d7918a774613c644f562506745ce8e563ad43239a5a1c7b670a7f048fb6303e116b066b047115578d740e86dcb2463d6faf4a59ffed8656c8d2bcd20fa86d0ed2d303f4ebf6c1996bbdf32ed744fb23f96f32a72855cf5af47b20e0e4b569725e9b011bd3019f0b53fae38a5e498b094bdf6b9e195e144e4000f42aaa9fccfc200bf090fe983b000ebd1495b779f5f708c68b98fa478a4ad5d0014f7ec5dc252512d9eca17aa8716089b8f11ff2e9de00510e961266f1bc60f6f65110d086678011506688c3f078b74bb71a09231497472a63a32de83f6e77cd64a0c9b8da9e4c5c734bf7d046c08a9c8ce49ffbfb63dccfc85635242fb977477623a9f6e9c30b1deb0dda44824a179cd9464ca462830978e6a4de14217245ac701c670f904147a20fd3c6107e271b702b66f227da5eb8ab31f6609043837518d5b24058b55b2909955029f59d85ab07fd32e4b9bac6bcf096e1c0a2d8f2477d62971fd7894b77890b188a5e82341585bade00669d09dd2b207232d4a8078634616273e28f6b77b5a8b381541a6cc63648f0f121e01ae12e5ed8a86e963379a80ef8fffe7db3a2bc3066aa260ca638d760a6ea436d1518609afe232ec7dbdfd549b21d28832d29a6c5d3415d94b08c8b00a26aab6c819f0fb7b2e9fa426da70b2b8e794d0f44c489ddf8a61ac89fc7e06;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfa3063be5df14bd9bb3f5ccac31390bb59216b9e69d0bfffd787139460cdf90cd28e907840d93b7d587641eb5a10b614331187b7196cdb1fe15ce58151e94501408ba58edded512540856c6875c4f970c4cb7ad8f4dccc729a65b54fa2954f3e0eab6b80d9f3e04f2822872197965767d75279ee7d6562e0a334fe908fd68732bb4421d7145465417ef16346df2fc01f0d70151705d5ee10b4fc46745be47e5a1d6c9118850449a018b25c3d7ece8782f4509d839181fa25865c8c01ac9b00c4683ce55632bc04ba1aa2b43471521e764dd718101304d851e994becc08a15e4f0fbdc32817e1f180ce386a702d3f63eb70c7f7dd5fab156ab50e16e42f2b7561d448436d2e3d90ec1b3a5dbd18fb520bb5251367f20c2b40b28cb70525f5cda0d5fc340d225b4cc8ed755ff7a6d696a8fe848aa618633511f6126cf273c6c1e385a02c33888a5e6049e896e866fce22119b47654f425effc8be8199795be764e31e3953ec99047fb7380986b26ba52a5fe377e256fb647d35fbe5048c5cc0b262de25727fdd9ab29f145c53d1bf332f0707227da861a6813b4cc8d798b3726be0e479fb431e38e1fbe8ff64a0c9a0bac8736d753ca1f673cf4a3089ce860e06fb9e88d9063f66f40fb09550ceb30df6d661c7adc0249a10153704bcd20dfb067b704f56e4ed7d3e9245e1b29ee894de82d47e7df3c074c57dee950cfcb776c9a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5aad2c9e083feeb845174217329610e1a63ef24f45ec75132805934f08625cd53cd662de8da7406dc7693b0b209b81aa1bcf59ac47343966d299a1d5823b7afd84e46f0cf14b46c4c9595a7ed5fef889372099cc47379b8183aacaded60f1a7415a2a0d966f0341563e1688a337529de2e6d780a9a6795c1dc8dc2a23170007b2e748e2f1b7d32c34731641f569712a7ab22f43801ef1f5cf600c186dae31236c7fe989839a3b386d85a5839f134aab31bf7712c24f4ef857817c6b1fb35385625aba733ccd72bb655d1f642028c9d5152e99f2d022831706bc8fd4b1929eba8d4319cc90fac3b611d4a0e904fbb1cfbbd011765ef0e571f4713016ccac43698a0a9745f311ce9e041b264a55584f381671c81dd555258466eeb61d7b2b69eb78a7398f2cfad2f7209fe6a263edb4de7be6d69515750250c7e4bdd698223c105e74fd62c5718e9eba4409987c9c8978fa9e3a6670f936868aa8e730ad890c066df8a2b399fbfc060ab8a5034d13eeaa5e16c61232e1ccf94377da1b7bb1334c85b0cb91aa4e598550bcc388122df4069864c924a230404c26407a2348abea82a6b56a5657143f6943b97d9619c27c2c08a730450033245182d9339674017329d96cdd332d8a6f8882f01b7633f746346cc6659dbde4478564a3391b58add5a0f6aded384f027ed7aafb764b48f9d88a3b3aefbaa2c5db3d2e6b4bc716adbe6ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h832d21134a832de2e336797785c0be66c969a154b0189e0ec61d441ec3ff141d97b9abda57e65fcdb6bd2e5357dd7fbe2cc6f18be5094360b15205d05ed372776c908d4ad6df85692d4cd64af0c940eb46f989727ca971dcf752f49ded5d944d0c23ed968d83a05fbc7c08fe5eb0bcb34276c179b21bcb19e913a84afb3052691b630014a36da7fa4b4c8ac4d5548214c8bcc159882042bc9a561a3f4c15293fedf15068dae806f58460b2ee17432d83ecdbd8210ad43beeea7797f66e60f44e955f66f767935b7612bd828c5d9ec95fa3350a9cf12d6518b1fa2e8ece04af4e6a7e4a7d42a4ec9f8e7b57104726a045bbc1122f881bb83dac15a0a5fde5fafd6c54e51dec12053bea0f08c396d972fd9a458b0487958988582fd1f5dc9d310385e86e2f49d05f3b4490b18f611e2d2f3cd2b95788813f44e1ca493652a2575056f7e62bb8be9c385781b50f77affe94409fb770af5930c2df8f188487ffda3d27d36e15fb70aec50055712c3d1de74d2b744d796522ac9827397468e1db170de64912f2fc713101f147c5fc12bdf650e36464189676b1741ea28b9108f75dadf1b3d8ed907e469d6daeba6d00a14f4b2cf627327c9d2aeb2c8ca8489d3599d97726f874b5757db93c0b207cc55e967144435f9283573b8219385be86f767c129469d5ad453d602df9342476d187863d4165bb0051b627ef4d481ba92e69dcc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb54a943b136713d7dcf0831ea8a190a8056105ac62b1194a7ae8b68eafd9fd4f16e81b8254272438669b662b7bfd8fc37682a69df4d915c3835d99721257b71573cba6dd6f6b38db430fed1785c23c9757ae3f35dd1835895b44cf95e4282aff349b4ee710f3b96693f8fe4ccda3c722cb8887c170411b859ac39fbee09bd817a37e415023b8c5f488aa8ea20c1bbd94bb777bdfedd900528d748f8c0947dd541636c74a6ca9ad55156dd7c3798b402b9e3f2046742bc89fe4fd66bf5cd4c58a9bc6db2828682f43047b944e75e35a6850e201f037c0878e373ca53de762c352fb514953494ab78f78031754ae711139188a0c7729112bf538755b366b99f7f393e1e54275fa49ee47afca5d1b60078dcd64f7506e1aa53d33f168b3a796221ea7f523fe48b8d3c9079b22d83341f4a9b2672118f3bce9ca2e61ecc65b0ee98c7d0266163b1f53f774a699753dc9155e11e160b7e8efd8c8c78146d35bc37e8fa47103a6701f1015a934028b1fd25b189794841568b154f1f0fbfd1630aa152c321b81b06ae32a1b17c9728c6e0d8c9ec9ad0dd61c97f153f54f8b5c975e56ca54354b1006e7eab51e5819d506cae2eeb5f091150dd420f84230b19048da12009703a064e2ef4ff01056dbbf9e9a3b0500dbfb94279e0e322cd62a2fb7e4d068822e983cbcea226666844e0bce9af71f64c38381f0a3e042631ab82ad864685c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1df9f6c80334aeb9dce0d49687308f9e4aab2d92c11f058905d2ff91205b6e681c91eb728ec1e96e5010b258876437488028aeb115ef1e79e9a67ea0f622d1a7c1828674689ccc596f3ce8f81eb2bf85540eb6589e431b8ba36720348cb500a3bddb85f567cd17211f5e8086acd2082326e4e13b06e661dacc1c242eb4e182e5da70c31de91b3c512fa36f130245743c96841e1d721124e27e0ad6de5087bd2381612c9ecb97f3570c590dc960ae375a0968643e634c6d9dc577bb1dec8658e7f4919428117032def3d1a37a777c834a028abd4956e0a2e5ed9bd01b682a20701b858cc20b570caa2bcc8f07e1b5243f4cebab7549244aeaba5055bc7cdb2c02fb43191c6303af6ed933875402a349165f2ffeb467dad3b2191146dc3b839b55e6834f556c9f4e6a4f3ab66bef915d7aa7f34eae1de502c4a2d1db08cf5182ff18cc69ad45d05c84757d8c44733cd1de8712030132b17b5bf3e15b4e6feae51129004d53fa1b3f42eb53de67a2ee777702a0b0228f1e9e28bf080265ebab065e99e686bdef6fc3b9e0809443d0aec749063f9ea7c5c3012e5105ba9e58c89a366918398810ef49fbca9fdd0f1fa69998a5237f382f24509baff1a545be80cb578ed954a4cfa3df8742645f86cfc51b4e6fc09796ab01d88df61781398ffab79a9ea622154db50ece9f23f56fd2a76cd377a106037d13bf5eb777a1c279aeafee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h24e75de8edfc8a343be4297fec4da09fa55e623ca7206168d2f5213d2dd5c547a6cb37a311bcba6ae5994bc5053be8715e88f26cd8d3f98634921b74489a0c58327ece1b97e6e21592d1554ede289a40b34464de1366e5f7d9beaa4ecd7aaa3e4944330df72b4d0935f1c414759400e5c547297fddc19a77952447a369b09450ecf257d9541aaccdcb06ae90dab1c4e6a0ab82a1a645339a7f5b4f3620d405272805a3d086c38fd156e403961e6e69446f1a6c1f8a260a1ca705223a4b391bdbc03b41b4a2d0e426b8447f7ebb53715840d3dcb525087a01ebbb279a02575a032339c4a36d1f4da8d73dbe6c3df281baf26f931ac2159e14a39e74918de7ec16bf4e2dcc63b4962d27704012968bbb72fd372f24d1ef29ec3bd850ae2db1311427584d6ef948ac209afed8a58d628649edab2c003fddb8f0a9ba1925eff3a78a33774f2bc1ad46ac2699a647689787ab87bb5b18d8870561375c44fa72947b68763736ce8b666a09664a3f6a923eace57e807a5fee11ccc326095cff16fb21ac8fd1273db679a9e24618c7024b678f68e52d0e97083b032c089451483429618ddf5c468c7537ddbcf2c901fdb8dd252fd28b01c106a3a98f468439f97b621ea414ee87c3356eaace414d621424ece8d26c083167334d97bf03bc5f7b9667d9ddae2c9180e30f96b7766995d842f10c0a562a769979253dd7cf01469d1d2a3a9e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h22d4b7966a4933bbbfa57ee8ad6e4d926612527672f64a4a63df9a58711c2725788a631efe2249130aabc40fd1ce091c6551db01f2c2393c06f30fe25abd13a1ec623ca8fddc7b0d0860f97ef72132fa512b5f514103efa447e5931fea7faf260fb28a6ec9e2c2322da298de41cd542eeb955733fbf445ca1f9dc6cd95dc9d4f0e52d51f96b6a0cc469dcded01fbc34e65353cba8a6b9c3fa571ad4794996a4921a5c4cde546619508aa41648232be379bf14b2466c2713bca03ece94985b7299c73dbcf7bb9a55235b2324b2deecb760f1c1b127824d268596a75dbb2bcba13839d0b61148255f49a8688d09809837e8e762d77360043901d211da78c4e5cace3447f80cf608197fec6ceae81b958af86cf8f5e6f8cef68dbea51d6efc0d8fad37b54eb9107100a058f3543d87fcb639f35e94905469485f2bc7e0f92db5b1e79f0c0501a9116b0e72f7cac62b1bcfe9a2cbd79d16019a4bf16cda2120daa5ed219c125f1ba1cc7ea834f28d952373b392c14362018ee0055ae632de5182fdfad9ed6b53713b4543e92b9ef48196db0aa0533afe7f3b24a154dfd1a1d9ba0629c76596bdd7e9e54be89baec08c2f5ba2a667dd6d3b406caa6b8d155a9f29f810dff387a12876ba8d6d61ba67803dd2ec0b36f8499ca2ed100db4b65dd869e9baca5bf5f638e69e620a8ce098927acb2a012a4328946293b35aecc4621a0cb18;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5a0a24b346185ea9ccc7bb5557f03d8f39208c5e2b50bfaefb202c635675feb282b835fc9422ec74ce30de1518b3c52dadeb00407e56ba8ae62f434812b371851bcd94628cb18f892ffbf70e917dc527e86d70d448cab66b3bbf3beb6cc059bc79a1daf08e0876d7888bea67aa2899e091e72119b24f6a84ab2d91288bc1ed9f01c11f5222cc4c6fd7455004207292c4c9ce5e1543dee8cceddca194bd32cf1aa950d7b588ced2010138ed6fc9d3304ce69920839bc660eddbab358920055bf24b5ffa7c1f961d4539891ef98a2f19f5d8846545b473992c541dbe98661b4e9031592f9ff2d8b3e4bd535d9fabc5af2342214ad1caa2f399f55aba219208ecd5362970e860005852575941e5c2725ff7073d40fa8abdc6a82fd50a5653c976019221f96a02a8187bdf80fd50a7dea6c9ee88a4ae3365b9ebfb7f012f6b595f38b0de77f57ebc9692d4a1246c5824f2252f2701a3393cb3371f71859c13ee763071a0743b48bc85b7927254529239c3c2da6487bd47037836467e370c6b423da000a15282279264d84a2559f8cf3b8551f722c03dbc03245b675c76a1452f4500d4b0f6b1600ce7f07912b156b06c00cf80dfaf0b7bca24865cca1385a63ae326bba6d3bc1c668f516bf27616069326393afbd86b94e63fb087c59811cfa80c0f0fd2f2b891cb9532fa919f8b3053db62e45725f0130d50708cd8ebe469ba9a8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14f5bedc6573f7d1a6fbbb5449b15bcf79eeb2fefeed0309419cd5fcf018c1594589182745b69ab6b7362ebc4859e1262b241a09c89cf25ad287ed2c253e728ef564abc948e6c76f5f6f6a6e22d27d00ec6b0c416356dc909c553441e662a145ecdc8791cacb13a9beb06a308b1495848369f5d689e932e0ba7f54a3d98b58cff05e8bf840d461c207653eadbc2dbdee74bab2fded366d45344089f649879efa87a0b0e0836598898c2e0b4bd6cedfb897bd8b9f3fe2e39bcdf798cc25fa0393ba0d1f3a307769d1a2e1c58b998bb827b35884e4a4105c211dccc5632d8fc52b199e169ffc663e14b9acdc449c8eb846328cff8cf3b5badfa9c35e53ee3f8abbbca8731cebd73aa5ac21f54fb76a8b3306faa0bdebc0c61bbe91d32a1f86db7b38143453010850f3ff98615be4de0e7d945dbd33c62b9de01a141180899f95a274d393a9375039d8dad7ecd2e3c7d64a1c21bc6ab8791d7816d1cacb1b9967d2c739f668f38162156bf63470c35c2b07fc729bf96c2b3c77a1fb817dc4f3b7d80f5e7580cb83525e3ca8d87d883ef03cbd8f773df19d6db59b50a702b68769654c3e87c24de6f2f404a6f6e57ba1661465ceb89bf675e3598a448be2a118f0c9e1330b17868b2bae1f0967afa883954c8ea1fbbc0a59c49e6e6a8f906f4db777b519248d29904a680e2386cf30128058862cc3570c3eddcce0cba580f7a52002;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2a8a3c50cf78ee2df8e942ee00158b56af3396a654fdd72a4b91e68269dd0a985ff7ffd6b326bf5e12c5352a6fd1fef2b8cd53269aed523c17adbcd30f4f93cd92f3d591149bd51ab9a092f549905a1b6f484e4cbea08625a901bc1e8373078e2d291366fbac1c3db1b99c63e698fc8b22cc9ee2b89ca03c7bf9d07c6bf30e7df5bfb962c22f8dd2db2ad7c99c5927c2092aa5784b90662058bb235d628222fba88e82bd59aa488c85b9566f310186c56c89baae0dc9cd5ebba51f4a78d281ae0a87e65ff5cc7d31a91cda1e5b0eba117497d47852e45bef36041656dfb74ba2b6b9d5fb896bb87f8f22322005d2b38dfcda90513dd66501a8b78a4d4a6d35050ae3652a4ee07b2d920103f1211b663d4b2a2d45b5798879158c54b118666c8e31f8dff37715b9b9f78d8f14a3f496a9ff14f29ee7776f6c34eeb56d7b860decd0c34b7daa4a10374f62e33c2d697bd9761221680163c1452d8c3f4cfeec181a6b4760703b8875419900cda745b2869bb52291e33d5cf9860df2d32d173d59125f2ab5f05baaa4b60e803d7a61763950f77bb470737f05ea3f5955a645b9829bab218ee8471d0ff5084de1aab387116cc529b38dee88fba2606988bab416d98f70a54bad45e1c67b83cd248207b7dc3c79a4d5c470380a0eb2ac4c312fd844156fa13d44ea51c28463a186523bd068a42a0ecbb191659b985c7a5c79876221b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h54a8b2c2e975f19ab2c5da0b399092d01d2bfa495505b14bbc3cede8d9030e6ee8786a7413b143e5dfebd43a302476cf4a2d4ce50d3cbd371a80bdaa8a3e7a9e21cf89e6b0da9e5b7093da34cb88ee9c3a9a07dcabe173f24761d291093324288d1026707a48070ecaf176f458dd05cca88be7e91a7529b2029c5600a2bbf2ab7ce9250cba8706fcec266947aae5a09cd9878c9c05dff28c19a80ec4b833cc7ccfc2b75686d869d8c49c6086891c393eeebb94abb0ec95450e0c8098d1654fd74b7d17810bdcbf5f847c669933a2dfbde7e3c00dfc15e26536d1edf7a062275adda4275cd78129c846a4fb37b4523ed18438faa4779db6ceca4100a1c6bb14733f99ac6f94d09c628806c707b8cb7a47f00a64fe63c5d8bb5af7d073b7ffa0315202c6ebdbf6548ae052c223968b877f2417826fbe75f035f9c9b5054e85e476860a1d2cd3a272d8a2181d38dffd2733d2b44580626f52a749665d6e9cedebc7a28b345eb646a645cfde999dd8729ff177c36adcadb0f3fc2e3fba602a0ea070a42608c4f60910ec4ce3a68c976b5905d2efa72d9d41adf5067ce3206991e037f744400fc1aef98a413ae6e6f83324a28e78714693766067101817e2f81ebbcf34923e66b5477f13c3e584a1b07cd988112f0796563ebb510143736dbe8efbd5e29c9afce5500c3ca72b48ce05fd4cb9e8ada6c1c932adb1de704fcf75e54933;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcaa9e344320d2ca5066ab15f47e4ffc7f921e1f69e3b73d85b7e448869996ba21924ce7509987e3683f8c34a0dac014d9e7e0b46b9111a49daceeb4c6bd5a02b1cfaa7c3e22debcdde8e2deed54eefc537502518ce181a03c8e415d20b7ac1b0fb86ae10fcc84bac5ad9dd5e00a5f8445ae248e63b8e51c63f858e1fcf943f785a2e15a9ad9ec222155d2b996832851f5c82f7f0340a45efa537838b03b8dfbb1df8e20a233cd0d6f20e6257760b4dbba769285c8dc970316fe5027ed337a783ffdde793ad73b8c1cf97de8ae3b659020b285ecb9df8df5484c5a8a81a914c81f9e2aa9d960ba4d3ab7bd58856870bcca902e9c6acca68590429a4523386a1fd21cce3483e19ea30cdfa7bdb11b505a8721b7d4f685ead03f458665cece8eba2455cb95d986454cb0551402db6b3eb01b5aa8302457f6596b5500442907bb3aa0dc1999b429170778d199697dc509e202f1c3f7cf474f40367e2864bce529c3e314ace2c32f48b97c392d625ac9860d947078adfa9bbd8a59ff49f420d85e6da1f0d3b480fad6df054fd164648154ae1f745b5651e973e46250dd018d760c44c2976f9633778cb6ead67311cffe20b58f13833e7b50b32345f6b0cbe3c3570a1f76282a9a0c41a671368eaf53659f1954fffd46e7c39a54f12f892de9a037885e06047f84f391d0412da7b6b72b13eac9ce3a3b59f48aba0db68306ebf62888b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h994289dd4bbdf9318d1fb22895eef2f2a46a50b0f896275bfdbfeae36f3cad8c1fcb49aea326d7bf1be4d25067260bbd7b44da90e8aadb55d419e9f0e4e61ffabaa482eab191517f01709c1835fdf9b93b73f1387c29dd03eb0c97f924da2f27a309c6d9ecd85273414093c8fb9213eb04bb1802b000c3493bf873c22ffd55a6d943207676ccf548f1ac37bd7b184988654301670ab56bbc941d24206dc2c95f7d8cfe13b77f496896d6f3203baecf8a4f4c39f972cea5441ddfaf6cec662eecd5fcc1ee27cfc4ddb14933bee6070991e313c81812a58e84d83e601792f24565522a4dedcc049b22ed4ecc1039480908d984f734a12ba97c6044cd3f9182b97a9ddcdbb224937175bf8ed625a5d1851d0b8acd203175407b8a9ebc9d2d9342adb0977fe0b5f3eea33efcd2c244c7abe1433db2d53f5829d9f4c7df71644ecee29c53c51b06d510196b7bf785554616e0e0b3398098e7db5a50cb42f85ad84840188bb82ed384fe5b56eb8788bcf5a2633ffc6b452e5816a24fc59ec9e6b039f549a342b4c2f1184515107fc6c8b08ba60c6e68ed195d2a0dc9dfc109bda9aee2f543875b50a01f39901c79bd6be1e09a377ba8a5999b1a9f9621cfc41e82ac917dd9c5e550db6a9209422cd5c3999d43e219afe19dcf7a3ea23c8bfdb3ab89e65cab5b58bb0b5eb896911bb30b0a3a17f095c3105252d4c163d3a24825a4acd;
        #1
        $finish();
    end
endmodule
