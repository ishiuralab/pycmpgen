module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [21:0] src23;
    reg [20:0] src24;
    reg [19:0] src25;
    reg [18:0] src26;
    reg [17:0] src27;
    reg [16:0] src28;
    reg [15:0] src29;
    reg [14:0] src30;
    reg [13:0] src31;
    reg [12:0] src32;
    reg [11:0] src33;
    reg [10:0] src34;
    reg [9:0] src35;
    reg [8:0] src36;
    reg [7:0] src37;
    reg [6:0] src38;
    reg [5:0] src39;
    reg [4:0] src40;
    reg [3:0] src41;
    reg [2:0] src42;
    reg [1:0] src43;
    reg [0:0] src44;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [45:0] srcsum;
    wire [45:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3])<<41) + ((src42[0] + src42[1] + src42[2])<<42) + ((src43[0] + src43[1])<<43) + ((src44[0])<<44);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa3d57a696b05d43fafee2053c831730612ed03af35a3b52dba4f81e38673b0ff4c4e520fd0763169c9465995f6024da5d49fe62d73e8add2ba0987f927316b9f1c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h912c8c4195bc2951de9bd687b188842146e8f1a6ad36747a27bc27570ad2fc921d3a25c1205a2f4e7ce3e64de12f624be0ee64006d188baf4e3b443c3b6578536e15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e9a0d811e9394e64816260dafa141dabd70a490db58ffe8288bdb61b3ece205cae1142ebc55f416bcc67b65456a1717838f43fef599febe7254adc2434032ac069b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12654133aef8366b82c43e533753133af1d2f90397ec4243eea2322e92c85552261622dfdf41ab767936786794c58d8b4449142a582927bed2d5e81b6b469c5097b07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2376e3e473d205d469b8930885773ec694941d9b0003ceb21f7f76320bad0656a4461c82f278c9fc4e658f0c98298a0bc4137a5d6d276270ce23b944446fdf829d06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4c884b1606a78e1eb4e7d2ef1ff40fafbf44e28164738ac2693c4fbbf517aeb83770b31de4c9eceebbc19dc855ed8ab9a66464c6b8c5a3174ee078b57479c53aa7e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87cb1511497ab1d6f6bcca8509c4d961a616d8313cd666d32c18f5f4705565995a8f914d0b7d3a935f949f5932f814005eb5ea65eff10b3802a33048c1b76ba59b38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd5f3ba2f1389d5e503a75d737c2c89c33b18469bb7fd0b2bd2475a38ca4fc319ad34f317a4ccf60792b71405c91680c32f19b6f7563da0399b3190619f8c497a53f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70efa6d1f7793b1e50bcd445dc5046060d70a43e234ffc3944ca37b155e6fbd20687d455c54a71eed24c1695d6f272ec6573cc62a704a2bb10ae451a9df81031f1b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13dbca101a411d0dfe1331545c2401896d285f70a2e29457305b71638e47d7fe5aa0bb07d18264f4b580c82e0cee46b5d1e51ae3946e34c6f21a4974150b08d63d7da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bbf58fd973456798da4608ef4eebcb55b9bb3801d197ee4c5b59fd3f303d1e90ede2887bc6bed058d822765136a34d80e1b011956e5dd29303574c4a98b9a3db262;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef92995066218848005746820323bc62b9c410307299a79c72aae97143bfc9ae6df6a0c8e91d2ae3836873f1d522005ed7108f06df532bb3b8bc79172fc2c9bd3cc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7dc9b4612032376a515189adfac2fed50626dfb284e55c324bb4e0a6fe1260f588b340a22c5394166dc54e58705128b6ce43ad13fedffb0fc701b9b776b78c550cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d3c70afb73960813bf0805cd58ae28885602a618ad38d427d240c63219c70b3a1ec2ed2c55516e3d740adbc0e22a71ce76b86e2b783d2248b32bb54cb6d9ea6b34d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1848bab8e8bce9ed6f099397fa2abc0a3744a1a34e72f516bdb78c38508405251deaf2fe7e3203faceffa82402581533c622d3a2a4b317967e82ad7810b77da33a8c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1048b06609e137352d00f5f3fac7b629b9090ebdd34eec6c20882739f98f63478de42c2c675b5eaa622268bc839389140dcc816a71cf4a538308972193ecfc185a54a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6802383234f5ef0269ba8e7f56053b251ec255cd390898e80ad7af4de57c8bc81bac79fd5e30cb4cdeb4e507d0b1248984b12884a07ccd5649bbe903033dd7672dc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57606c754804d6e2ed7a301c41d6a8a35ca61d371f1911f1d7b4313b5f0d7d550ab5cd6d51b7d13102496cd351915734f6f677b678dd0373e5e737a981a78bbf2f8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb057824517a9c0d32ea3013ce897a6cfe3e0072b5078155d04b1a0bec920908b85e4fa6e9c73b55d46d623a1e48c52edf7ba24b6ed33147b6f657cff64022a4207f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e580562c5281214d74f6d05979c084d889611c9cb520f07103e19bc5c8d7d255844d435a27d77568049c6cb620097790f20a708322e9fe4fc93826f2d857ba70db17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec8b05c31b3b102774562f4261d01c8cc9904f9bec41d377fbbb49a769d71ddb64d34dc2f95c3a506afcd251ac2ad54a50bcfedd70405a1004a976f48251b9fc50ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133632bd45b92c4426119eb7420a20c5dfa2a823dbb5dbf30ce02eb363a00c19bea3b2f7736d48c4f585a7482498e76f89e900fa601684207940167c4cd696bac9f24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f3d30adf534d2230086da2cc392ef5ef1592f29691a5482b3c49852727cf5c6c899f0257544376e376fd0d3392fdfa90c04e1a3b88cec437a1671cc2f241c123495;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a6b86d3ba8c74f4748533cec57b63f55494b1024a88f90fce27f5c70d1e0725a1106004f7251b8bbdfab79c6efb0aad28d01f687b075c7fd32428b8fdb6b7780c91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185bc51411f5a8488aa98e33a47505bb2d7bd4612f3fe9e08faeee97295c1cd53d30bf71b5f60ed0588d4e0895f12fa2e0b88f12d6436fcd5df335c9716a7da7b508a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e2f629bfe36dac044ad7f7f910cf80e2794e60de78e2620af0d89b7b67ea7e9beb387b1f7fba397f5a92c207d174758873d1ecfb17afc47837c341329abdc8af29c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab318671cc100f1aa96a19819b2bf5f919a330d751931a76b3db060b3915b23eeb0c169602e46fea3fc223b69abc36adad640f02b5962fe0bf9dd9469ec876eae176;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb109adfcdcdf5dcd61440394ae7b73049016b1d74d2d3a0bf6ea34eb187e19d9160a763a0533097a89a1a2e386e0c5e2d9c6fe8322708bdafd08a7b40748c3f5d723;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86b670b09adc54a90663f8042236855e4e4cffa9d7f8e2a413c5af3de76e8d0eab238f7475fe492470dbea33510906c566bdb39e1430be4fc4cd44ea0456ae41525b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fc3147436d738c47865db3c3b29d0715e8ee16bed4e60e77d4b19d14ba2260439c834ec57b369bd4e1cd78c68b92e652095cee66dee89010e8dd67b566cbd5e56f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb97ea8695be7969e1ccb18b72129393ab3251d7bc43ed48e9b02b4d45fd659c9eafd3c5eaea27c62793e3d099dd59cb84ad560d01c870c1124bf3912ebe3e185560e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h931a3df4156f19eafc73a676c8feed00c715cdee047a44b14ad3cf0b2c39d03290ee5665c880fc08c4a33b07efa26b065c6c11e5901752bdc168a989ed868be3b8fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h590afc5b1b941dba1e6a126f9c51d31af7f48b48617ddf48af6a60678de819ffb5b97e38985b5b0914e19a33d8e018ace288a76a802fd7522ef950cf5fd36e9481c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b9e5515b748a0cd378ba3c7464652e2eb505855163ccf6d0a41973f77fb56c12226c437cad057b0dd2f3b2140444733f5bf66e42b46fdb322f1f82767ed55353792;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141413bf7ef365dde90f51fd0a30688ab8f6308d4c33e36d084200ec583fcab4cb2c2d87351efcb63fbd269105c52c0e1b6df2691d2d9252f5656792a59c6d2f3db0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44731dde45dc1900ff14b8e63fd7aba7b867350c7131d774768034e9ffb340ac9ce7b4bfe3479c94ccfaed2fd16cdc7f0e2fca000978a8f9fb4097419bb152e723bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135fcac3a9e9c10fa3a5347f69ed62f615bcd1d9be22b26e48b5748eb48f3faad7d11b9f9b8d40c6345654b4e1a5d6bd45374ddb7042928ae986cfc63c6a3de606894;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e26eb194d558a24074801119cb96c93dcead55e7fbc144d7e1c50e671c3465c8b1a3f12b8ba25e4203ef0a310acded68a200dfe9ad2121770294b9c80f128f08f54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16668ef96073ed777fc746eda586ea2290fe995a35f0f108d94f447fdaec066185a36dc647848ae09f22e995cfd9d46bfd669c37176d267b4de404407bcb7d9777baf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134de4689205f5bd645b0b534bebab66684aba9d1a97c8549c0e39a82b0475852bd7e0990e36cbe374dfa2f6d1c6ce1abc0fcdf38af6e743ffabec5bb2c5eea85c143;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h233dd673cfdd2fac4d15a7fdb274623f781883cdedd3d782eea475ccbf066cd81d88c64b2f6fe8e3fa0c1acbf4dc1512d40abb38f762ef647433232366ca894d066f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18414a52dfbe9812b8a611e1b112abc497364f8602ab581d9425ecc3aced15794db59fd9238b3c291f4b5260028cc61618d583ca50c5d526e75afe76079557e810e72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h787b5581e905c96c96ad94570a5bb9148ed6780c7164e6eaa11730daf305339798d0f280c2a570127155eac1c1608bab9f8c037015f085fd4b456185532513562871;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d5b642b5096b80bb11daf170ee7020bac168586b1c3d8887c17f8f759de52298827377fb4663066e78f203a8dd8f589c30710e63303c3e49f4d3f145366bcfbfd73;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42a705cedce3994b7703df1e23d0d6c9b47a29ac27d60f8538b6523daae67d5ccb8582261a8ece05eb44b26ade8777fe92390a34fe5a75e1fe7b27402da8c481c92d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e26a6627b4ff60d6241f01e1f1aa7b5d8f4fd377d42871e3fc0496a90b2abadc64a33929de4feee655455e244a9d3ee44e992a1892ce5adcc06bf9231cc814f61b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3513d0dd94ec0d29e0382074b0e74cf02b313485894dbbbb805f8e8f695d4555223c5daaf3a72aafbd6a57f07910ae851bfc5f1daf627f57cc96f1b22d8077ef95dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106879c520e534fbd7a035419027d33709903fa86e155a34f9e944260624a5985f12d2f4ac50e729892c5cb7edc1821f2f606008eedcfca19d44e3ccd6341d1e983d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3a2f248d5fe922754d657029b13566ce9e9bd78831ec20997494b4d6ba54ce58c9fb4e7cd6aed207d130809ce28d1cc167caf11c3f02a9006ebe5583f6c6aeabe88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118460119ba2ca65c51d843bd2151843824b5182a9c6b0811b39d3fab838ff9b819bc8d997d3a016c4c1ffb60197e2532a2df31efb952ee63acc5909882cf48e4d006;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca1f92c697d4830a73cd9d43cc866db73d82fee93a7619ebeb644e358e867e379c9405417e282d055f08ecf70ff132b0241b1b772459b3b6cc1938c5313094cad134;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8376aeaeb0bda721387af91fde663d90da336da413f86844007f0f74b0306ba4343a7bee195d331956c6483babd0273bab0e2cc6ae98afa9c07a5df45e6663dbda91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bdcc5f642d0acc295e671c5293667c6190ad59ca10daa2fa14300880a20fb81606fd746aa616083bad479031809d162c06df4daf2091f39c852b1823e10630f69c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fac0ca961d62d9991564fd2b5b8cf83393019ce05a48cb9d714394f0d670ae1fdc8cfc6cfd73957272d07e967d920ee4e58883c45b514ec8058089bdcaeb014d384;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19de96af4e7f107aa825da7b8b79bd1de666e8abdf2aa032e1607311c77d22ff7a0b3c68a12559e42ab0e8166348ea4b32390a8fb23c1a829a6ad1f06394f3792b36d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1017640b94580053e42cddc12d6c0fca864bf2e60a94f440e73919c5a67741069afceb593da8513cf06c5ba93397b7c97c635ff976ac35069a87276098cd4dba80e59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17915777bf1fa9cfbd55747dbbe83af0f858c31989c98f004a03f9a1956f6da3e67e61fea73486511fd1aecc722bc6c200b38f6fb5faa06a3c53cab07dfdfdac32572;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e7c73be85f2e32b681f0a7ac1ef69fd2e1057ff159c16f77e41b0163957c07e5b869da5818b2daeb940e75b740b59c5e13a9d74c88917d2af8bbdb4ac11a4573285;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120e656892bea7c5c87d0ba1c2fb3dfa5f8d4b314473e2c453e04514286f139736ae88296c6704bb82dbb5d4c1cc36e2647c5b655bf812df0189ae2a269209332bc6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a30166958b46d341909edfb12354d5e2297e4afcf6e769084b22f39e906b0d9964ab114ab5000f986f9c2c43cbfc307b1f23ce89c3b8f66a9fc2f3212bb16aa21ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f62787781444819392cbe8e688e34e3c181c40a341d3443d1cfe1f03ed99f25b3ca3cf0742cdbea054e0bd5f255e9383ba62599565e6fbd961ad6c7f7d6fb6abce0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164d166f586c1a1c4559b37e49c52942ccbb36d3531bdefe19333bee63cf41270ac9e9a695b07a43c97189d9d80c4b2476dbd3d2969cd98813183d4ec5b07d1efeda1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a7f226063b209065cde40424240b285c349b68ef7e8d8fcbc328815ce4424c729dc4563639e43d026f6e650f6111b160e36f30b89327eaafc4143fd1001b7db6060;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45e758fbabd9e7df10edf1f8f01a3b2d718d96bae91f75c88b016bfbceecfc30ea05cf20ad89f8372aecb5073591fc7433a21e1cb10a90dfb1e0bc076ce43378462d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ec7453e851583ea811def0f71759aa95363632dca882ff6088b4bb4d4335159161ce9469700ead98e8dc4791e4958a34432642c02db610c5a7c2ef45c6ae8be5768;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46ee59de7b024b64791bc9ee0df8d6512300f6c848f5091757d6ac2f2d3d40be653117b92715b53e7f5a8a802ce63427cfee75de966ae488bd0e946683d6911c800e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he77d631ac57f4adc2397bef3018ac0d72f5c0b2fdc8ac07969864e89aca5910a89b4f59f7ead5ce45de0bf4e0680f7a94926b8bd2c81cc825b784b17665b728a609;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171e69d86f56e40f186136c0fabf11b865af293c2a32e262464b5b6a2d1aa7d4388f3f47242595aa6d9127090ee6c7737d87e00412f48bccd083dfbdca4fc284e5552;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156b9b5efd79f8ad1ab27d4f181557583f5a78ccf1341733cc6ea670d5c6191d27cc1668fb42f71804de5ef1276d90425df026ccdf84c114d5e02d4c1c019f7ec091a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183c3c6420be916d52a87a9e32605960389f921d3dd4e6bb88f5d10b380169afd047eb4c5e8cd64c76edcbcecc6e4fe5b4a517d750e769ee5e54fefb89318926311e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he083a926fd44343f17d9d0e5f74a3978fb7d3d8ae41eba3720fff9cd636e9dab0210f369923a1d52571a1392a09287881f82f31dcc455c6f47f089a95acb4fe3f8c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ad6d196f5b290a193d1dee031381d7927e2354f5e31e1c79ec64a6c8fa6a8eb3b1e201e9fa0f2eca30bc1343745f8f930d6e3b7bfb212c0b851db9baa1ca4afaab7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1555882b0e1f8b92301f691d77a005b3cf0fc6c37efe2d287878a76d809c796d15d98beaeabb950811af7121669e5b2465ce499581539f99619bc65e80d7c0c53968b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b646c39545153f44d277512298a2525df14b8258c19e8bdb456adc8b52cb16dbb0ab67410432a3cec4a89975bfcd55dc1b46fe7d85105bbd14e4354421ed72c69841;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12836915391c2804eb20abfeb1501bf260e713e86210fe81a2cd076b373f99a743f5d00a1c9bcd3c4e9cbb630b467307ce75d95e6c91193ffef103e9a1bd3989a97d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e07c2f4e4173b0d6f0aa0c24ec20783647502ab1a3a7cd2fc80f5e474a93fd35432bdeb36aeb5724d2a313875def63f720d59b51e42a635bbc6f3dd70a991b183c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b643ab15cd3629a617de077c44eb1a610667781f06860529e6c5e49cb3a091ecbcd7b46f5c73e9deacc2a7338a1afcbc1310493c3d957ec34a9ddfaf988c5af9e269;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161c5525538f1a46fd2e50f0ddce534b744078338435cc1d56a1f1a89038adfb17917afcc77719a9ac82d27531d7f8c61a0f78e124e14e3f93e83bcb05d0da02da1a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113c5536ae756dbebd4a7d51222254eaf58d663810648fdbd92885f8bc62135c81d4736287a99355c02b47d49e1a4bcf0e9031224f5d4dcf9a124435e23f47c29c896;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef730e9c8c21e64b95ccd9c05be10ba0733ec53ecc0e986e297224159a44a49596045ad527f15061331fc87b635d671c078921c1a47679e21883589aa91b38976126;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160ec885b3553f4300d0c2f367b426f82b7a107676a117d1f467e4437a708219a9e2a409949c9026f3bb62bfa32d4e8a2b01269fa5381913637fd148386d600938bc6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b52fcd9488e8bb61f5c069b4ad5a018107017793074b78e9bf219191b041156842331bbf2b2fbf72ac34f344c5858a7357f8c444640d326257cad6ad02b64767b57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf8321d406c248b606d0f6f92b5eef202df1e5911476a9fe481535701dd9981adfbdae9ab1e69e6521c3edf7a1ea27f695e1b37770d0fbd83b2f66f78cbd034c95b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7934b1b17458795cb2fd435fa11ab5f11c9a1e713cc97357d131917f0f018d26d65d6dea0e9ff0f094bdf859480d0345b81cb689553ed0bf451c268d99cecfd45380;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f05aa096748b3f3d89326407ed0e17ae2c41d63aa4a5dd09a92d513e26fa12ad92785487f51dd38af5ab0237925284fe82c1698f30748e4fbbe45ac320d6f97c70e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59bc9e703f80d3b4610d9e29792b546c96bae9c888f1e093e726003b0495ab815710a9962622baf27425b406e1eedf86f7a2ba2bbf2c5b90e49319ae5dea4bff0be1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1825c30f8f15ee7e0bdb99d61b1be66f6aad43f9de51f4f386be17cdc3e587bbd122c35e34148f7dde6f14f4ba13eea2210f9c4880a6b7d501ca9dda96290ff85866e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdffb78304fedb52fbbaca72fe6bff94fed7c3881d64eb362720248e177486f71ceade92205fe20a9c05eeea820d2912eb383ff1524dfd7a31bdf1206bd6271d13e4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5abc15e3ef7a701045b7090fb0d310e8504a3d8971f8b3f2b9bef685ee39f917b5487755b90f15b8843c71a6ea43f9fca4a0370bb6035550f28a2c767950676cd75e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he08f5fa186f450edf43adc4a211d34aeb40aa9b8e518480d1af8c8a67adcf3941b7e001fab1ecc8a6dc7643a8d9c212746ed2da42dd922036bde4285735117cba4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd6a1ed4d0098d59ddf6ccdd24f53f15a74a32b51b636f9b55dba586e31ec3ccbd92c1938610fe77111187bc6a871a50a8a0ee42b56991f845efe72ccf601c805694;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h830046195c92a298aaad504d3e981d9c140200583bc9a0312fbe85de49b8ee947a17e4394e9ba981a65edb6ec4aa2f963e60a376ab8db0f7d027ab340ae604bccf99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e8eb9550cb7e7fb71f089106b90d1ccdfd09b13c69b43ab16959fa1d43b95858dc6e6ba12843e2059b104cbd004d37bc8ebc29b7188d9ed7b8616a980dfc56034d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe7e4cbbbdb066fa1b4c66a0eceae05bc2bc8e21efb19920b05e383d3b678598fc1720cfcb253226a79a64b3b54b9c37a7846387986aefab68da64aa16a791739da0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1412a05cd509c16abbe0651ea986be97536bc5805d37e7f9817320297e07a7862ee231863b94217460cc265cbd560b30ad79e768ae7ec5d576ff11db3c8a828e82017;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194d28330f3b87ab41981ffc6974aa51c70331ffe8af2b85222fb065d64aeff5a34cd310c50e988b5b9dd3d95aa4a655b91d7fd1c4d647d32ab3cbc6a0f1d11fb63f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe72d8d89c84e0e404ef9e83ae68143ce86640bd5388490e9e14be01925921a4ae0ce547853e6fee6b759672281aa7af5613707c7f4070eb894ec4a9c83dd974cc36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1814f6287bd10cac20ee3b1315d40b571bdcfefda9b31beccda7ce4bcf105b59b820ab6f73faed1360096056233145e09b212ee618c3901215776e326fba7b2a4f036;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd01bce4c8469dd670a64d768fcb40b74f6dafaa2cca2e78298fa42846b629c37e8a9015363029a130234fcf775bf4531ec11f277fbaaeb645883a6179b712dd0132;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e7244cd5b63b61c23f0bce105e01c13c2094f613df7b4c153dd7f6595aab1464e5f82e2523ed999626c07e8e55cb36bbd226d6e2aca678a42ac1617a3be99a012fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd685b53d0cfa833c5c84167abfba40a185e36a3b9c19443f70b3abf48cbccb0d0223acdaa745f97c00ee87a25faa49b63cdc7970d19a4638a54dd2d355e22e6d2c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103f958970f32fd8852d80588e6c6f111c0adcb33b5b75d69260616d7f16da4c0d19c5b1b45a42bfa527186823e10522a341f070f696cf3b707fa2bdf42b678c37435;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1537ece2b56fd29398e6f9d5109bc41bca1b5b3f329e138747f9de72ac453d8c490ab0fc6c2bb1ec551c989ed51dc2844527853c8021a70ba36c5d6a5321d66db1022;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f8902dc1b3ee9dfcdf3157835e124bfdc6c9ddd6364f02b3d69e813fbc175bee5842e33e8d96356270099a82afb0dcd385fe42d8a338343d5ab75fea0474f434e5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb270fbba34f5390bee7f30f7703f0f3b93424de3a7e608418300ea61f1792ef7f7a123dfb3e3ca0c0062dfe61be7121f34dba304b801f79360506a23bb8e040a3b17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a9e1b7b20decdc2260958f5a52cfbe9b94580a9854496b54b4ac5fe116f406f86be739e598cfbb34a199dcdf9a32ca0d29b66f1d27754a1dca4a682c636c0276435;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1e64a74959fecb2579279663b8257438e0d8d43dd98a28f9ded6901dd45d1826ef48143be960ec12ea97726dd56b56f4c82f4c9379e9a66a567591a60d92a129322;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95dd6fc1a20749dba19242ebac53b665df2935ad9074b868dffee499a91bf57339c7e6d02cf0ee4cc081a1ee64577751a8c1befdfada79bef20095f32c7b8c77c832;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14333748f97c3f5386412fd2e6283c5ca1147ccc413dd9c6353af00d3a6fedc17f3e2fe44271b3fe5a17fefb116c9d22420bb6a4ede8274a62e6814b502cbc939e519;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d29c4c5fd14256960cfe26ca7359c204be788e4b6592adee0b169271c73a15155da6b2b7b02fd7377b598a32f53c5487a833b9ae677211d7b8be0f62668f2373e8c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16de3d974a2ebde1a3504c02842cf4545efeeab665bac64fee317200c1ee9c3e63a2293a34233b8cb1a862ebcf28bfe27f18de92e3438872f86e73611dba4a88cc54d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af8be5a62dbb4ac595c3ae9550927a3da88bf1701749929f9611a68173293e8ec342b33cd2af695ad4c18162cb4ad1b5dfe9c7d6af546bd997912dcb12073ecc9215;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc85df5d7683d36d81172a1b547baaa2ba00a35e06f77c496b87c14b4cfc15865a88fbdd275d89cc9fe71ec848447c2cbbb2e7719c0f8a84cec57ee97dee8d52c1530;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b046bcac485f95a1f0adf641ff9cce4756e9a72641438d7bf1386a0ec6df578bb0967dcdae10b157e8c37856d8531373d58bc698a2dd548f9a8d3d76dd8dff5ec0c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8a34456aca16cd07e9bec1a4a4817f8a4ef4fd93470d5d4bc284b7d374bd3f2d9d19816b3110459a7197bf8d6cfd696db95b4870f7cd01cc5f1fd3372c2aea3824e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb68df089ecc0187d87fc2e843c20ad5dccbf9267decc8f8d63f394800c6d67a855ffcdb08455b119a9eee2ff2cd0bf1e6fa9069fbcceb01c4def130fb01441c9268;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb5a66c7753b4c4f444469825c7d0e57c82af317506e13d64b7920dd53dd248da75ba9f362791817c07eb0dbafb2d60f17364f319313aa5c10fca9d89455c9a761ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1812fe163646b2790fdb49bba9de0de62492a7044cdb650703f86c0930cb633c49d13c803986d23dc555bc0c608ac2d354e5ec0e70afbb051ac2d95750bd3435e3af2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e57b4351dcf9f8baa746966814d4c96a4c0ef9baf879be33eeee4b99962e1a46f21f4f72fdcd32835f49bbfda9e804848d95305fd4f4cfa94edb70183c0ead206dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7630028fb0358a5d1a01c3461de3bb9e92208569820e7a86d763d99160ff3bbd8c68d6a39c7a506921927f164da7607ff273e96b8c72a03c0809f6c750f08e0c779;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd04a3ceb867679d39e093e267bc174c781e9bf4fbbd5c5ec276941233575491c7ae7788ec6114bb941deb7515999df1058f6e4dea1848d457087d28a39a84434393;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18df749aebbe39021ea156dc7dc27e972c9a29b7747ecd4ca7fb3a412b7a139e6504466a485ff5cf9095572c71b5c448c85014f7955a7595a467aafb089a434cb59bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150cc571e1dca66f1ef35df8fbc3990ad874b0e4181f4a228da39f48cc5c916261569393753059dbfd35e18c999ea58a99362d41ccba27cb4e2f713ac420f445fba35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74b6c13c636baf46f48ebf67f77f4d06489024442ade850e05fc2ddcd3eb794d645f9a8338db040d63b9c035f500c243ae31804edfd6e93487e484464c4638f31821;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ea9cefc06aa71c4d58711bf409030e88a5c41c7abbc50f9ec9e0fe65b1ca0ea8fb7208777258dba90d4b716e7bf2791a76faf86b5f51fa3d90cc13243137c22f5fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15362815196fe4ea7d6ebac8e3d961ad3e60818df747f9558ff5915af51600504a41e14a971ff2a7b380fdf127c55cfd1049adaaafcbb8f9ba103cf25a82132821519;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f139ee96079a86a7b6407c361be17da71b5db87054fbbe4a846629908ea8a3ed3f1cf3699f1586da053e507ff9a2820da7b6b91c3d6a9ee12edc3e55d900b686665f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5836ba5f9ce6c9f5ecf7e9e4e23ff155e0cf0c24b0967177132df3ef2ee5e3b1407be85c2a8c5b9c49ad299dcdf075b5aaf32568163728ff1ba0129a2c8cdf6984d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1747ca6778a241139bedca94898733fe456a769ea2d0b504f58a3beca386770d1c80d19ecf6eeb6a879dd3c58424d71f84e2d6f6a9e508c6ba1fb4ddf8828f4fdd040;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90ad9c265f9b49b8c34f4547f8cb0a7aeab3e1f229e6396d0177b730d337a15b2d3187713cb141ae142173405edf5e41f117cb8870b8423ef3355db2c9eb0b1267a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135bf3055603df5476aa10b3735bf4c52c3961f6b6a18d927418b2f9f08cb51a9470c332859fbb8f6935348b27944aca49160b71b66317104d5e3d1605f488e2badc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h494d00eaebc877da3c604e69df6b83911de385719d1ef8aa7d9f7700851761fa532f43b2eceba04ac7ecc8f820c3b2869be78853f44ae435a3973bd3357925cdfaa7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60a9c47f4179c4ab29fc2efafb0ebb4d8df622f2737eea03350d4562a0a1336b38154908567f7ead101826c40f368b9020f5eccf77449f1287adc09bfcfe0c7891d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110dd2bbd4a72515b1cda1af524f0bc34a36f238e657e1b17d1ac8f37d6732967ad637981a1d2014e7f6547e8c5eefc20f59bbc9bad8afb4406857e46f2f28e290c7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb556284dacfec4231b754448b5247299819b9e14d82608f5ed2ff710211f9a20731f4edeacc3299bae1464375789a7a72c263d751da55ddd5c83e3b6e8e01cc9f794;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a44c1ba237996e9ca0acd12bed5560c5ee6adc99208c05a08360f3fae728d02e2d9543474b59602b60055560c2acf228f845457a08a08f2246623f5d6c4b17c3c6e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9cd089d4136ab93db5540e8cdcf0498681b908b8a24b400ac6bb5a7c6e0f0d1ad1f1705b30a5c2e6b4f0798b84cbd7fdf22241b1c6830156e9b86c40a92e12fd1a4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1989177e5f8c4fccc9bed1558d974bb516c802895d596173437a5df9636338fdc1e2604610c98f9eef304ad5762df980d54fed6622526760f15aefcfd5962dbbd9b71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf240933d7859959635b39afac1244f69755809e279567ddea3050b7bd3db97f754c6064e19427a536ce4f7cfadceef435b1e50cf5f35cd632b4df40ae38b03d57065;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a98de7f8927a2e285f1df1570b67983d7aa27baae6d43b4afabd1a5f2b74e79c9089d45c088cbb9f901e4ee5ef32107ed42bd647873e0e579353d1a6b977a1fb48a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67d5d8a1a9f516fb4fd9ef329b4d9dea220a008355d0675e67baeb51d9e2f1e5a7bcf2df4b207dde7e32324a8542ba80eae879780c010a80197afbcfc306e6474;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc742f7aa8fad844494f0084f65e99739e721803731861cac9398d0f9658d1758063b49f5f90c4832d76abe58e3354a8423540704d4a3ee040d64838b15eb8cc34397;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dfaaa5bc9b7d0b58b033461ce1280b76621af8bce78de05509f03546646e444c897929a0db26b51399c9c853e8eedb75206072388283ea0fdcad9644018675eb67a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h739edd08dd76d3904508ab470c0ff8867553e74e3e6b8ea7b54b01a54b863a4bb40d139ef1f26ac8c7668823f39782003eead052002b231c7c5e550e3606294d00c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ed83784ed4844ea12a607adc1465bfad149652e7f6d36cb863083480b464db0c45f81edee68777fc1ae2af8c878eb8fc04187b21935e0e5581d78c6ef98de60a0bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1861f2a5d248c87488b9f240c697cdb0605c2bde0b8d797ae0e168fd852baf2953b35af273cd6b25f74132d7a835ff186505be2eeda17cc965a161a68641c5125e7fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h859e92e8469c2f2f147f167bbe46cb02350042d81081286a17743bbfb4d0c173518a8759b9a8d80016b7bc9b8148b187639533021f0e484f7293375b9a574cea30f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ab0b834899da75faf757201d06f03eefa62e10aaa7e1c486e58a11cb91614b312bda4d3bc7d780b8b9b009bc4f3e7b0a63ff41d5db06cd419bbe6dfe97f17cdb2da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdcc6fe6645d39a203cb66a030ea8b8916207ef1c39b51b10337c9f2a0318b2af912bc25506e5540cff84b73924f890a9149bd689274d40c534eea22ef84422bbdbbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a4793d92e0629859828ad98e38c43226c6dfe7320af050706074c34535b862ffa6b1e54de2f5b68856ebfb5815cc4d0fc30061882e3b1e308833d33229fa8bd8b9e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19435fdea1ecd3efbf36ba2a10f76843521fa8f1b6dea3566cb5ebbd58dab3e48e5bc9da43a199de607694547bb0ec5122d43f947c56c742b9b99ae6b03c752290306;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h33d55751f722a46e9abcf63527d81f8846b5975991c238fbe4c91aa579614a5ab86620095218cab6265afca072127cecce14f256ecc5ff16eb1698c2234a14f1cbb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7364c007d4696aebe485e4c84dde251b1c9c6b34073388181cad54bc400029d13701fe930fac54b0f06ab4319567f2f6038457d22e2316ccd03d3a0b603a0176f945;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f785f0e7912881cb6571bf4d3591da4c0e5a8b3bd1ecebef1a6063053fe507ca1785d1344e2f45e70060061a96241c4b0cd6432c22a0cc50b1565abf598393f4f5f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17392f27e5fe6e1c5e93ea4ffaf3ff9a88c032b836bc773156f08ef2f097a906b1a559f30e86233029f8ecad968be3ecc6b8191b23a436c61360124efbd4f7f61bcde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haede9a9a8d746a3d0893ccd56f137451680d1162cbd5c6ab70cb957fefbd7608b59e8240d3816fa1fd891e706a4856a90cf758cf62ff57498c47bebb55482a2ceb86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfaac6fcd82ae1b924107a976e9770ce9568a62c5b6a842acfb9e571e4742b777fe3463a33e3c62ab2635c6edd9eef201c4ca4acc7756ff8a8b802249eed9544986f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfa0bda5544f61743614c061aa94e974192010639023343776edda2d0213e4f3c1003e6b3500dd3212960cd7b9c7dc902e00f1fbe8d0618f225c4403e9b463e1f7e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bf95c95208b2cc1d2110defc4fae0133ce9a3a742a9478f7c19f959f8449b7acfb624db2f5f0c8a726a49c126426989ddb6563d6dfd819b07bb20dfde6e06393ed1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf6bccb8062706c514b6646cedf25618106435a225791febaf8fdf750e8bc6f144884f2f73295a5740eea1dc5fd27de108f0c2092fb22cfe005167381f21b9ca8156;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12af0e4662aedd73f7ecdba7bd3a279b9dc3d7ccfb3f588e5acfe4a30140dde74c1f34263fa7054b414f024fa87680244ffbdda2c8a78353568a3bb9b524e9d70dc76;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haae1bd82964a357e16bab48f3679a54c63bde85b74ef2e1c479aeb822429a1b59cb8b3ae3deca09a446b401f4a6e21e66082da05c58d26a9891eee3f1ebb46c5b427;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1321730add14e3d95697c05b5969a60579b98cd17dc54cc9f5c35446877212fa1423f672044aa9ade7ee396a76e4272cfc1aa57c7f571d166fc0ba043065986bdd5bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10edaa910910799dbf4f3148a94aefd82b835d781a312a3a5fa4bea2828c2fc4917a8c06f924bd2e079bdddca4998f091c2aa79a773c9141eb186707995711c983e0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ed90d3d1fa7c79d75a1db5480fc4d383ccfb6c28ceca51890442a11efe624c4bc1c4ff4ce05e5db507b7d8367344da23308d8caf68e8d2266af7830fa270971cc8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5afeaca5f58033779d7ee42ff02dbb29d9b4ee30d4d3dc0d70ad4e6c8ac7453659217f741ff14272285102f2a32fe0c6691d87e0dd5e5e912cc53bc9b1f43e2ba917;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3f6f41c82abc423d0aeb60cc3983cd7585aa22d9d465d27332ac8ffd90bd7114020ff65024796e68eafce552e8b250d27f7f2ba8c683cc44d886d1a0fe0f40daa21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149ba9d573a6b453580d90f27455b26cea23fa02a689634cb4bf6ff4c4ea5123f6748030bef51b977f094383a9bfd8ddcc574c9f2c69011431f13d453f18b4bfe4e42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154ec4b5aa6580038b4e6ce4d85eba69f64125f0a9965b0df234aa0949de5e27faa9da82b229ca1ddcecfbd70b243cdd6e3128e9bc35f7ef7a74845c7d04234f4c1b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cc3c33d6a753889243c886190c731115aa55acc60870e9ac50fd405782998c051bf8f123535dca7eda0d530873875291e23f3295b883974a4b61c06b45f6b3491c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dd0a191036f50509995e3f158725f0867ced622aadbc819a88e8d451b17fb94200e48d7ce51db07c45e887e558feb182c1c5c215ab0124054665ec3fa1666532c71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac84e5accad685de61a246531577155e87ae816b55134fad77e4732e10f0c509f17d11da4a8226bd596124c9d8e1e407bda0f0fd93192d4d61b4ee4d56218fb77b6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habcd046fc466e109a5a27bd77e97218280824ca7962072a66587471663abbc34494409e6434bbab7839430ac4a93ee618fc42b1a33e122fd6ab7336a8375549f68cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba868336f72edc311ce0f82cdadf6ed45e20d53798320fc25bc8ad48060957f37bdf018b8917b7e3a5c211a5b55ff8a8c8e15d92a912bdc06322b39b77da75308d12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a553d68fe33c8018f7f25c2adc5a99608cbe28a42cfed14c0f44f4da6e6be57e370097c1ce549cefbf8d883f317bdaef089e7bd3e65d24744b0120f370bbe034c3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146a60a315c9c2e75bf48da9219b79c98d3ed043ed95a2ea5ea3b36c98aca1cd27d80c62b6d18d8f8f69edb28e6290aefca3460df817f188306ffd178d7c23a341de3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1478c9fff12baee3c628ce983a81bb000214dd59cdaaf5ed1f2201cbe4802b7193db20eb0a18d137a93c940a41dfd54e149102a032b70ec3cf6d90f444033a962bcd8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b0ecc94cb2c36b0ed03c5e99cca344cb5e16c5357357bdd64b72453a2ea019b2c3e475fd67b8dbdb2fb5b1722247b66aa0b56a501915d103a909813a6f708bd65f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149770e42673bd27922c7a8d99779feb838f0620c11dea7028f2cc47038e35d1564b1762ae647134d1ad81cc4ff58bf114952c04eaefc24ad1cc75bb5145f82f3afcd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d56fa17ddc18b1f79f29c575c0203440b0a2c3cc5606d6714eacd0d5795eb873ff4e89d530ca5747b163c60e7ea11e6bdea5cc220731d9f84adf1becf62d16b6df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a65c101402ce1a376f46cea82af86052a8ffdae756b0dcb7c7bf12c2388d6f2e7a0ab3e071a239c0589f2a5b364859041db093ef5470d7dfa6c3b7d0ad77486b0025;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3c7e17830f4ef532266a2c623e22f87158ec4b37389a3dfca5a15267a6389dc3a97bc8d787b046258f80460c00b866ee7a8b0fd7bb23a00a1c8231b3c2e8e61a1f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177864279a647e6ef1027665aee3fed84423e69d89d11ca12466e55de8415399fb5fa54217195481baeb614fce5683f97258c04886e51b48663515a44e9e72f2f5781;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73960617a1f11bb8e91fdbea43ddf13e0a44ff1ed59aa33d55abedc1228f7f8d6516d3f2f838d52cf1a905f7b1bd2bb2c2ec71c6fe2f0b2a73c819baa5bfcb5eaf0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1965a87e0bb91557298942bb67dfc112dcad6c424290f6d9df97a98810a6a179b1d93aa8e0c3e050ebdff09fa75fe9b7453b9b2c20dd62c786ef7a7c7fa9936712333;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e25a05cee9be3b05bc7385ec955d13bd9820a326e0ffb6928d96b255edc2215c9965c2f16750d7c2512e7b40014f5f066ed106fee4dffca1089d72274cdce5952cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bfc55bc599c0aa1a886a61fd2ee1dc26d4249bd8bcee9c4534f0954154e82005702712b2e5cb9cb8aa90a13ef2470fbc39f43c6e9ac950891af9dc80dbee857338a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107d07869fc91dc2f0f57acf2f669560d172bdd3071e47f4cf9a88d46163645f33e359bcbe0c3c26dc9bdc85d65ebe8e71a0a8747513d4267ca32d50463531c7d2b18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c378c3e85f0f84e8a0934d93ddf2d4d51601797b7c4db506ec6faebe86d9765fa2388c23973d844be0d6cc7d748de7ed3d6fef9c7f28acdca59cf04092f4e453cd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0df1a96a24005fedcc4ed9379378128ff77f2f11ba9e6492a367e153319cf508ebd5b5c10307c91fa5573a071aacd1628f5de5ffb849e8a3aa1040aa04ef00604c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180f222ba57e0dccff3f872bc9aa10ca66a55abb43dd4009aaca8a8df9be9ff09f1ce4cad59b40f29abec18b3d796eeb099e7315740c7bb8c40bb4eb84c33992b4606;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfe272eb96e488b103e8b4d718c3bdcccabe5bd30a340e034ed1185b593140d06fbe6150b875bd6d6b519543be9b1b175beb5f21e34110453c09a944518b45e95840;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8793508f31ccb8d29d518d707a80e6971b0b7847ac23d0747f2665aa50e680423770db048ceb91243855e85abb3c168d0800eaa6f9b73837ec2662d27a30bb641894;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9146b96f5ccc6ae935829a6d36da196fd6512546debcae31f16124e7bdbb6285662e8e6d5a07fabc830b26d3062a71084704bde8100be2e06f6049f0c61de97edbbb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c305a499039b346fbe947475905535571df50b159a79dad279da2882c4d6606376aa7fd8ba7c73cfcca3115fe848febc82a8e47d081e67d831be845559a7ff98809c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8bdde10f82c9a173d42f5efcf626139e5581ca568da8e86870e820b46c1922af502a8fdf7938697e99f7508c8555835a2b5f45c471125a5e32eb2b1e7b76b02436d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a549624c997b3a5af886a716c153b3c4ebbb477a1770950ff5201406308e744a350191282126ea16b4b42bed7b37fbd7b55535981b20849af0f6891f87d8529b273e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7b48745039774eb227dc097e9fca0e85e6030499aa62b95cabc056ad1a41006d4637e368bc3c615f5f0249039286600a6b3fe56d967f58991aa1a3de8daf3470943;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15607acc4e13f6b94c930c106fb5153ac01560fc2c4a094dd8398fe0c3947eb2b14fde162d50346e0457a677b128733d8deb43af8003225a6c3ef5831b753ba1dad0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h556589fa77c2742fc067660bba0ec8aa434cc695f8d19a3643cc96090f6acfdfac8f1cb32d253f0ddbe9f6371c624a86d4fb85c26772624b094abac4cf72abd3ea52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2754df5a02f0b7b53642bece9c85cae455b931cebd27279aa3288585bdbe2874f67409ef31378879d6349546ed147f2d4572cd43a46dcb0dfbd81964ce5fc14a65b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e1c445df0f02c23151f8b0440484f03eb0a43cc46dc9d11629371585daaa2805c870ff51d413a70e0d720b66f10c1e8f8acac9f7fcc4732757004ff55f6b37efa91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h527dace89a510f8d4e6c19a49f189cb4cc2a51997473a19924150a30859359a871aa0b5bbc217f3603de05eb8bb9868761acf630a87cdf446e5399f5eb93b9c551dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b4e7ca13d7f19315932328ddd6033ebf6d4911b859cb5ca70bf1016a40b4ac62e887e90f342df9c201aaa772a8781fd37e31ef8a39fdef80b1f4c70f9c4186a2641;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0a453eb2ccaf3528939802d60b7109ee2d9fa948614eb5216da50c5a24a3c2e3d76dfd718ebe58d3dbce1cabce36a4482987728ae13cd254b9dad0cc26ceb9e7d37;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ede14c2d30e6be5a0311019e14b14fe509a965381679e06a0c2e7f209ded103d97e6c62fc869aaeaf7f03a7e9af750bebc8d438722faa694203c9e5035b204d07da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5b710e4a1ffc04f8bbf9e0e5fb5eda8758efd2e264e74ce77635462a55f61a5ccd8a76f1836561a5d44f562113aa10cba011a7cc1f25da4d6c0b175b6f55eae95df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21e4bffaa23ee79a6d4e217af78c14458fd38ffe7d0fe5078299a28df0ba91563611af6280cd7d14ce361d153b58f45199351e68754dca68229b6245133f244f2de5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169ac7250d3e9cef65309a74c1ffd24fcf487dcf31792ed00afd32f257852a301adb751d00eca10a42ab040c267a503ad95fcd721c843a2cfd5130dab5f5c413e6ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198a01d97f3cb4a03f21a56a17a05abf5486647a39a3fd7ad5a7f4d770896628646894e9640c957bd35806f59ca08fafcecc2084097be5311ce08a693ecf6d214469c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc13a56d097fb7d64e52a16258a55fd4f8184a4e584d8b2173713c4d1547db66d9a1e72c387f1b01841e7057b46c83eefe0bc8fd6ef2551002ffd2bfa6036bf78193;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1468796d9b7e66a46dcac6fbc6f0500cf8beaaaddc2b02949e77989e12d3750d00f79f74f958c9139b8e2ddcec5d7367ecb333d37efad4a84b89fc502af81e1f950b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2226291088253f2b0884bd2b2f4933f497e6babca3718ed19ba9e7d8d9f01b354c31e706f75861d09f035793084e4089d26a324d8e2021bc6c30ee1659a099e6491;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a6a26e3c9461333c8026111704abe9f3861a98a9fee58fd996fea1a54bedc4555a1c41ea915dc5a2c9166955484d62d074325a5e62907d6b9f9e7910e19397b888a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h752d0fcb6621d123e51e580eaad5f093784b8a22389f600bdeace4276918689cedc3966012cd9bf6c7fd31481af1ca82f87377657e7d537686c4ba46d1064b04df43;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9704b7e2f3c79b2c1d53dd7217d3dbf1c978a5bc7d4e77f511c397078ab848ddc080eb95fce8ba1640faec3a3cccb784f2af8e6d58394b8fa3530210d634a466e146;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c376457825d8cf925373b92434b784e9aa4f2e30a111f70c53f07135b9e076dd4310c905214945252a9805d671fcfac9c2a7688ffbf63bf6f24b170e4e7667252e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aeb51e3b70bd2cbcd2d748c4d803e4b36c1f18cb21e4c9be8bbc02e3b1afcb91eddc69f1c259005ce4095844bf8befbd1bba89f9ef9d673f1f9cb5a3d79f4a4c68e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f26d96acb4c5dce8e74d7218c31f8a84908e200c135f252596722700680f2cd7303d0f02966be34f4c10d5073b2da5bf9b64d9b38835f53c501565fd575909a8b4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b813505942f99f23574743ecb3b6956bad85bfdb00bb29715c0676c3a193fde7a1ab88ae5cb17a5f88ee0ea46a5fde6a8fc213cb4bfb4338ef0af61532d5b899dd4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c46ed3e421cf924380f8f5ea5813bccb38d719222858175ef0e7b90796bc5eb2573ab595f96d13fc8bf86026a82aaf8a73fcee7b68d1c74990503e7357cf123525f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2761319631ebd8e0243c3ae94d6222504c347af96059e300c4c71755a2f28d4b4b0bed200e2489e353d858cbb32dc601d56ec813658a3ff8a544c445fa5525006957;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17eb6c532583982a7c6873d27e6dc8ae87fa68aec8467ce541d453347a4691ab1452e42e5fcf58be698c9f72520c7f4c1487a77f50fdb156f3c79f367fb07f6922af7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176e9599bc4dea2707ff774c08132462c69dd991438981b4eef00a7cc761c4e7ef77b4b640e218ce1d2834382834d2381f768d61db9134422ff870e34d4b3033b847d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae4eaf10de87237ae45f58df259d28e8b9829546024c0916458ca2176accec27b843ee2b03417d324274201b89f01383e2986da6dd0af989a365de5e1ba7c2cf4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163f5e116e39331e8badb204f689c993424f05f6143b042bcdeadf17bb3d2e0c94cba005da7ce0d2ab1fa96289f0b6ffc0965ff67f64b989bcc5bd73e59984271a452;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a24c51509aea47a8a20aa93470c0d9e49e19ed7c5a8d6737ed52c18bf5e2c15fa1e0017b0958c98071a7794cd98281f3e066cf444793a91f36406f0d9e6910fd479;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaa50fffb300adc38ba7aa5dfa9a071a38f3a06680ac338954d2dd2264c1ff1cb8ea732976afcf98737eb430cf5b7948c516bf6f1585e2ffbd45ca4c1d45e4782c53;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1220b27a37f84ea0390071dadaa9f8e6da0a7d046b59c398d3f0a54652b53eae1ec36007d91f1984a32b49be1fca991df57ce1c6e6eb5062c814b749948591820fd4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fda400b2be7051a21ca4ee9391b16c021f04c51a8bb8be33561bcc82f176a403959c71b2408f685080443feae3079149b837bd6ee2493a0c338e40bb936f2cf0282b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1555a137b8dc3994db6f964059877cf9b4b00a55860052da2ad78322dd6cccfd39aef57053bf6502dc7cb7c36dae73027393565112368076534e9e7f927ec0c936249;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153a250efd54e27e7e906f5704b6c9aa63c0d41b4f2beba2d75b621219c2fff7ee097789a306843dd8ea5df5605334325d07738bf80a661e0a39d9d15c70bd8a17405;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d1fe62341d6395ac4344b55ec231e9e02033d3851b126d4b463a7fee9def08a61c4b4c794752814d7f1eac871eab37fca5853e52eb4c8994c2a936803d47924ff9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77a3f23a6372555314cd586be9450c17f6669509c7b07d548f7b7f3e9e34e940c28e33ebe34faef09c4d5490ad5221ce776dd64071b6a32f946c0c6d6eb44bb3c2d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80b091a913b507083e001caf233796c8437432f6ced9285b0a3e63af40adaddc913a62e059f33dac636fcfdc639c8b48758ade7f8facf4219cac4b1c8670cb4966b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f2c73ca1dd43ec58ce5f00879fd9f34a504b6eb5dcb00b1d872ff5e293e42c24d3b90c9a4a15b20e7dfd0aec9dea11cc77b59100cc0d6e9b092108b7ea11c377f68;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habaf9eea9a46a32dc1fc791b8a2dffc7432a17f891dfd1d374aef80fb13b82eabaa12d900984791929b2c9e184dcb828ae4744a196ba0e02ba7c6e247f93cb1be253;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2865ea801869d8e21b12fe174a103d94b131a202ee77493d3ac420d8a3859d724c8c1cf78b6b647ee3d74f66fc7b5c4031913ca1ba2a515b972241216317cfab5fcb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f087072a9f12b5001264fc5ed04ae8a1870ecb165ae0b3588612f07546623a6034c7bc5e2a96c73cae7ca09a7a78e72eee530e39112d71b10ab54b6d9926789a1078;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8da5df2f3512802f644b6d8154b0e95490b0549bb9c998209f9aa07f26a9a2c10d3b55baa5168aac550a3e80179a1ab35ebfdf287495a837738bdbc1e233126cdce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156edcb21b5e7f20ae99704e84bbf2afd4c47d768f124c86ac6042072a848c4163e04ac8c02687d7a8b2ac2899aa4210ff8927a5e8a34bd4d8eb9e19df9015b78d040;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd65552384d340e7c902fd2efa78b1ba14a8822c4be4cc83f53448ccc1ae9bdb903f62d8de66ac2e870005ae6d6bc9a65b3f451b51717583cbc55a821eb29dbf058e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h747a9aaf6d3e007afbbf480b868b59b62f63f9b42d3117934f00c6b268d5d48bb5d2c9b926e63c53e21765e5cbf860a3b9a023bbebd99ad9f28ef6c676f19854be0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b88bc50f5c48da8fe8731753e9c25eaafe43c37822388e1f333a1ed6ea7de4338e45f146e28362792e098f9f6647daa69027a7bb40084ea875ec65fd0c67296e62d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12fb7ef4f41bd19d88d1c2fdaff9300e6d71120141365fd098afe497fb819dec04c4f45437cc5aa063a15cdc9ac3faa62c50cde78f489f324ef9f443d8fff09c67d37;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c470c2118f01bc071aacf43e22771a196ac24dfd9fc218f301e6d7584c7ec8be54a637173db932d50ea235f12f57afc62767194514c2f7b82e967cd39e370596d38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cec827d5776d1d4bc0e93a8ffc23084372952dc57d2f1260fa5fc2c37900639487338cce3828d158d138223d771d5ea7f825ca20ee4ea8a53f9d988a4791d0e45f12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6a5a031f3c345e90261b72874a46142303a7af3db4164b2d72b562f1ad0dc14b9b87c783e6e91745646b0053e55ef30f9cb6893ecc1af59cce3f043c20bb9e220f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde280614dfbf3e72a482d6c37e11dee076ba3e13d174ca689d73b6bf1e5c3a3afcef65e03fa48c88998f8d842e3a02923543d6b39336eda4eba87040080db7fe4910;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a769c87e4bb319c00e9eaf289a6b85cdce469e96f947de3bbf6c5a16e5447062d8c2e3c9baf47646f4542d2115f3607d34f4835ddae3b7c7415e773edddd3eb36854;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c2061c95a4c6c6c00031de26787604417c9b302d0189ce44edf0657c5c6a2bfd9d8c350392c863cad4bef2376ce1ee67991f9024a44ae3a75c0f3d1b48d77682d55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17287bc58f219ea85ada37fa82839f35333da827c1c383f6193a7509f65541ac0be552d6ce81ef3517c5774b85319b421db9ab11c8501fbebf775aa5e6ff15139c048;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcca8e17ede4eaf3ec036f4c43c90b878dea91fbbee521c3ce482c063fe535183697bdc6ab2fc1cce44c627018a0bee3b6075ed56710f1d0d30ddd8b2a41df26cc7b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cda043e1214d6e3a3e637280d3f030e0acb8b0d64e6041c7b95fa97ec322e53fa2f655d2921bb1bc5226497bf372038d328bdbe7e8f1d46e90271b045461f570cb7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf891b1e7976fdaf14edac4c732f2008394a2c2e840781c62c4e6bd2126b7c97db8dd846c415f23c7fab787501a94591067b9b84b4b2c8721e513e8167a9a00ff2dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61940f47c29125868748588f217298b210e4a4b73f55a3470cc08701d5a4de36f689400d5b383a8a3d7516bc6148c1a4292e76af5b97e81e479424482417ab03b9d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150cc5cac76a5021e1e2b7b7bb06e9d1d8aa1d5a8fd9cec4f5b8eee7dc20ec7501e54f4b21fc31aca381a06cc6cdf92c4f2628d526699f4fee144962bc66b412cdf20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42257c2f560b1119b37025860dd44371cb23545ecdf5fc9f65b666614b5e7d40e09fbc2e04a5243e3e4ca6fc56438d3aba9111f356431a4fee35ab4f0bfeb6c94bb1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1457fe9f7393b3ffdffeefa9c8a7a576b01017607d2d803e3577f4a264097d02054ec80eb0931e36dfa320f422d646d8e7bb70d70c959fbde307a502446fde98f35ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79fb061588febbcbcedf64e9886bceb0d5016da2d3458c005dc5e7f2d4b1394df89dafc667faaf5d6e74e3c7d63f5169ad876ee81d8775b17a59761273e9d38af0b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd21ce738ebd871176cf284e63412d8a97bab21738875461db65dac42da782a40b6cefc6cee8e8a38756d43019d0829e1d1ac3e57a4f3c52f76774fa7eaf6315d6ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6047a9f5d2fb12fb2749d7ecc33a922c81e7a9fa140cc36e3a761d06b8b57b95ded15c5e270568c0efd1602fc832e127d0cca188e1aa64e05e65fabbc845074bb1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b02cc0f9725e00572f28c8285e68568439ca09951726b5020df3ff28705618daf46771554baaf5ad3047af8ca9405f87e36a558d58cdbabca475c3a305705d189bdc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e796cab3c5992305246d1f1d073822931797771490a19f65e3c8490772e88352973ebb69d6fdf5ccc34127398a26f282028cec10d29451f0c280f9ee25f7229785a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1201c7a5c2085cc0118cbf45523d1e4c2f4e0a0f42b7288ab3c4083c08a919516dd38bbcd294ff56b13658846881eace2f3f2211c04da4998e6b49e9cde373688349e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91a7d3899086290c1eaa63def71a13e226bb1b5ccbdc14aabcd6b548a06d807b9bec38d5bfab3aae60b92a48fc2a5aa2a73344ad71d666cd714000b5e6eef890b17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8650d2529aea375fd99dd60c01a882604a75125614a57c40f86fc41235b556d2aa88a28c5b14c752fb8d067fd73e9367f7093615eb95f058d481fbb48a755334e9e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8026f908e478f35f812afd6617b86c0f847d45a037fd1773c9d0e5f42d47cc31898d27c23b4a9992ec9093eebdfd645bc11ff96ffda7420c2df150f2cb31c2f9553;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3afe3397c25f1a14f69a09424ca49cd2418da48035f3ad19f572b1336c7da4af259b23f9771822ac01aecc1158eb8b46ffdcd8a4dc94bbb2d51b490a4367da72ec9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1998e26bc87ba286bc3ca75a931d0e111a66ade4ba90b4c188dbdeabbbcc697cddeade915b0292bc2d9e009a300e9640a0481de5993b8e8dd7d12a6243f367bf0c278;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc90774254f908384f79a3a7ed960a11f0b7ad1a9ecefc66646e6fa01c5844a826e3047168a4002d243743c94a66dcaed2d89657e9dd336bd0aea5ffde7c9e5429fd2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24ecfbaadb30bb75ad58f81ad5e1aea972a3ce8c1910d4d9e4c13dc681f98e8f466ceb757d6c4f259365edff775c39fba2b94ae40a4215898f37a9100d26c6d79da9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c6580d65aea8b7b8e5d4d6dd5fe9ec2fb03113a991a036137e205fc418280b24a104e31e9eeea0c8ddc7d4b84c6186d1e2da4ee1e434cae0682912887fafdfe6364;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5b16cbd16a37a9ab590fc5fdca2da5d873a0495d8cdd8af4e9540325fd41892115afb9e2727760fe1e1761d63118464bc564b20d23cbb7feba500e4ea34f64f3585;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4fb730cf5a4ae81300ee4733799339ea67b76972606fb60c56ebb4981d87d4a76745798744013a027e285f5f2431915d52ec381149e35c465d686de807328b5eba46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9fbeee05c4790ce6da1b9b2d7af4c2c38262b67a9b54a1db4c8ce40984c19412ee1761befe5438daa113bf0e23af10bf8b1440787e942b8fd7561130162558dc76ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8aed80e3c9b9bf8c9c6aa6bc12254e003118fc6d9650eb8b0f09ec4baef5c834e333254a10f7601774beadb1a047648f953ca9069bb7965886c6a6b08ab6e65582f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea528b89c633f98ac088a451e869beef051f50f88dfde7404d31d6d3b452e26fe396b4b69235bb84c38759fb3e92ab2b4aec25f4fee9bc69a1f6975df760516cb9d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39bbf3753bfb2eee402a173f49ed66af9771dccf0cbb9a2c36a9dddae85b6ac3ce5de13ff3ec90fcb488b0787f32a14102531a406368ac7955baa2d40471eb33848a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9794e833886bc9af0ef7ec3056cc953503f548b674d013eb6e023305a987245addf6634cd41237e91e469497cfa040e1fb256b04486f0fd1d3f861fab0256cd0058;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68a4e5298c17533fcce67f9677c814fdd2d8cccf2f68ad89132d063d868a2d0e247d460c426d034f815cf6a8d062b4b7a34f9d73b7fd903583bd474e4718bea9fc68;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1550fc6bc88a26f919fcf6190d9a4df425fb0d6838291655833b1dd723328d2ffc1907c039ef779c965bacb6785df00a9550d2a0f15d5ef9425bc66489ba28f934db3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185c38e6d01bb8f1cc74e828261e444f70cb25f5b99be25142910b8af2649e2464abbb0aa3672cc0f6d50bfce91cfc0c724b48456a3c61e1f2ea6c631b69f738f0946;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4b1aa8ebc55f45cb31601ba53389e1e07705d31fabc4fb15554835693e6fb7ee5541d1e51a9d1113091ebf3b000da24687e34dfe4d0a292bab50aaddcd7baa0c54c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h989ede5380b916fc820c96c3efed7a0cfdf07282f806b14260e09c55d64b4248ea9537f705ab78d56ccae0312d5c6b8c854689cb430304beeab008d6611faa9c3eae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17dcdc194b208db3b1a57e08be85fc5d53af55de3f5420c0c85aeb16ec83814e2e1d493f2ea11b226ec9d3586b14858b779f7fe499bb37a30a0025779464dce8f82a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14938609393fa7458d05b9655056e6959253c826f92fa384d477b31dad7498909640b4ea8440d55c707249e87ea1e5eeee1873e3e1b0c82327133871692a0ceeb3c71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f27a714c497195606c9918f379af18793fc273ed209f44a696e9df5073b054a86b81d3ed6cde9550131c6d602de65efb97fe1c5c6e855d10fcb48ac3e27fa43579d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11862171e390b8c46e7e134930f8a1789aa3086a60697dfa59377536992a34806b4f1620915d4e05d8aa4b8b1c6954bc6713c7992b1414d2cd5f8f53ef31590774764;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h814db307b6cf05599d4f4d213cc589d9f33a2df8c7f2561f1ef15ee09a58ff392163063288f6485b781b35a4bb8f1f53ea56f9bbdc9009af32d0050985ed2e4a6d86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9f350b36c19704ab29e1bb4fb3491844fffe1c36fd9066213f78a3c8499958a98a6b4a8ac62cdbd648a2c36f1f1eda727aff1e73cb7368367940a273f7a14fe38d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108117129d835b67ee777437df975a6b599585286a0d96da6ab0ddadde376097665fa61aec406d6a84ac4cca3742d27920cc70d8995476fba3a5cf9fd8b81d9266fb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30bf7c506e8e263036d590771a839708f36becf741cb2d43ba398c82077844ebad72720bd6c79d747025b3ab8e4d885f9c72b284e4463dd4a26fc97f0299fafc557e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1708fe67d30bbabe8960140527ce32ed3ad01ed90f1b6094ec26ab51b9b23b7d8a817fc81fc5f847caf81a8be97d6d42f6932f8fd8e047e8247cdf55e010109a4f32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13597307c66585c994ca15957beb4122682c43b27e2c852993d4a0e45663237858ea7cad4dadea21abd824732fd9863fd2d492437198808416388cea5b77cb4282b9b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d0e45f3970ac4e14c6e91d8222f17f0388fddff596e6c82a43ca8381aa045fb2a3c240c54db4d8591f3340bb2186ae0444a7633cd2f7ea8c355a83b28084f8bef36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c0fca0e01bfcef98d815f0e22d4f80b212d633972553cf638917eba1a7c3d3a4d5824e0630ec13986f67e4b6c50e42f9aa1d9502d00d9f11cb33618c9a3879f480b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71583543e95dd08b0c24f96477171f8611cca30bf6d5ebd63dd097920504c18d172272d3dfd1a4bf75d0011c746597ab11c2a6b1bba0a2244b9aefc5f884364be150;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf56f98402dcdc09875e36c01e723d8d26aea681eddfee0b969cf3c2d337f8d18c823a217a866deb4d8eff7dcebb68735bd4ebcd97024342634a3c82fae6366822a26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3daaf431dae4774742f8d9de5d7d423c5506f2f897ae74910b32c54299a51d7eb74a1d146e97e6cefc03940fc69026a83cf2094c4ce41bb709935b4f2421ff7a8582;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0e9227f9e174942f7834d6f7af7148f226f8fa1fc96ee3f01a4932b64f6e37ea37e4608bc0fa62f634731841346bf32e0440c6468307e1d6cbd3d2672751447d3e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eeb63077a4e89a789f07b4801fd40a0d395232ff56c9a00b09b2876ef427ff73a88e733aec7185cc7e9976b17d38de45aee4180268bd62fa85656104a106994defe5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113ffc5bbb9b48a0db25d7204345b7da42fffb61a7e61988232bd0ceb577a8ea962fd1a4b7ea6f7e7e022788572ffb6f3dc92bd2f5309eef073b2bad62f41f8ddef5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5ca1fdd96c59145322d7c11eadb0ed01d0c8cd56101d1d2b9c73e35ee744052fca01c27820010732cf50d224e625ac8fa81875584bdf5030d3720f80e2288196141;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193d12f4cd569f82d1fca16bd26dbbbe8ee64d189ce516a9200b26b20ebfd3a825f2846011b0f2d84e7d3ed7f34dc4dce645a0c3953f71d3261338e3c2c47d74d6d33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5597b9765717662ef7008ecf239080cfc606ef4b45aa3988e5742cc463685d08fe2ee51b03da82ed88d29ec9166cbac8fbb79002abcc6c1c8e35ef84c6a79f9f7a9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102dde7d8b592b3d1856b6a7449df0cf48fcfe243a3f9e7c432c1499e7b1383a13aed7fb4950965326e878b6acba3cdc51d2be85ade96f643a0a4d5d0b495e0de3e25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ecb098729d4157fcdfdd3bb32386d4ec9f2b27dc8f38c7b76177abfc40c93d657debe0806aa8542e805a01c94e0670e96da67571ba27d4fbd9830c9489d71fc1a47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b263d50e81fe8b2a1235465d4b9ce9d497fccc6cf8f1d51db125bdcbe64071918a1f670587e9c2c18cb4b7406103a1541306ebc631a0e6f04b0857c6fb37acdfafa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h847faf65cd1e52fd2b1796bec71de482cf29f9f53b492c62a136a8cca703deee1b090a9c074aff64717d7786f306615f085be7ee4b3870bc13bc6cad92190871a1cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b7f394ec98bd8e28684d3a2caa27a5f5995ce67cb70c4f3305727ef683d89573329232b43da73b3cacc80d39df27ff7a92332b6c922883574f20ebf4209ddd76119;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f9678283a507dc6c16e6f15f7e8f6dd27b859fbe84f5307d54f135b53af76ac79f3505f9b789863dd0d623d1af80e601d22461b42804355e7ec63692bb91ef172f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1255bb12ea5825058451f10f0b5f95440c813536e9a20d37c9bd07a0aff44013bc74d89c2d3586cd777a9aa5c8f52f96a86f307841b964744310ad76659b92585a714;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37fb57556b7f70f376b79f2463e69f8e28ca3c7a294523684d28eedd6d5e3cd38a698a04cc2ceb2adaa507c222fc151afbf4cee73906643c6ec693db909fa55c902b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5aac0974204e190bee1b08ee64180e021026a94fc2743da44b08f1c4849e48ba4a57749042591d08a67154a360d57f2a92530f5c65e1692ced421955e47fa9f1b034;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h517ec46800b2f8e77f883f86fd51e5280f8103c5a44f42be9ff1b4d3312cc1ce6ec4a6061cbaff0dae00bc211c1262c600a1b7a3c35a89b732d012760c4c8cc1d40f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1348586737a7f6676fa6f2697cd3f829401e170bda7a04495643f31dcb87950e5ede38000380336b970602055035569b5e2ef2d23f3bd77bc49ba7e1e290f46c99d74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h355a3230cba0405507bb0c4641a311f83eeeb2bc120c5de025d0075001e608806a0bd6003e8aa5d7f91b236951f65d81a098451cf7fde8ab41fcda905193518ef47b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fc415ce545eef74361d0d5e18e7f4b17b94a8ea2b47a295db23480a1ff60fa9d5a8d3c7ef4c24412464ae357726a4b8d73f53a696fbe652597ae6c8026e7390dd96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f1fc73fa35992a83419e7ad7a5b557317d04068060c91f2581f05f6c9b1c47f342f21a98826f001022d0ec6b2396b98d199aafbed2bcc1172bbb816e3e3a4ce9b0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a27f9d3e2c5f8601d8907b37b16a9def6bebc223f89fbe300af13e8abf68e1ecc026fb708f4a04eaeba172f5ba78ba731ff2c5acd899f7b885c36a3db0d3a178bdc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18895e572b063e13576e8cd2f890e597658ae2515e79e230b2d0e421b14f7839a3ff7a5c7a17df3da6414dd136207be4b7e0e25a6661b7fb472f7a5509f88a3a274e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15723d6f18b7440bb9a5e58d718289cf0801b47a81757192e799f5e114fccd0f018047a76b747826af3b956be817d52a1a73e10c694c86ce83205d83c259c881a41ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c62234e7e54b51bf763bb3c7c789262a46c4a3c48fd5ea389c5be073f5145cb42f9eaf376998a5d4db0821c93f57e89b3188b14d694c53f19856515209ec8aa0809;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2d555a38fb00ddb1a9271aa17947eb74054795fcc969f054727400db44d79c925107464d7f12b4557bc6cd3cbb8cb55939070c0df915dcf822b1d09a2dd4312d5b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb18101278427476a61e51db86039e3939030856608d43fbae91b9e412775cc9a93fde2ada2c0ae044157f21b8bdab2ce8e566e1b977cff9019e7fc67161e02a984b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13142965e7b92c15c98016489151a615ef0aefb921c0925c28e37102ef57e63a095f78ca77d1ce961310c745159ea8b640f78f21fca32d3514e887098adaa571a8190;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c87c3fe9b612ddca6f25562149c7793a168ddf978ce376c6ef091be5d1ae07b78ddb2d3996e7015c39e351f54343689b49390e0fb358efbeb5dedb9e8c8bc8e246f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91845f5fef24e74f2d4b7bda6c0d919d1136038d27cd3fcc62a8e74c80057b3f0b1deb84958ad4f5f8ee408926bccf821dd38c3a472b70e5575a8d825791672f56bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h676719520dc57264b83eec58f9681837375ab13fb923e41a8ab1a83a350a831a216e3d75ab2fc75852d42d94608ea9f8675490214264e3c3cb9833caed1e260fa84c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d2f39c714f5a7e012ac090a42e99e86f9b9a8457f82cf2744f6fad0f43b37684f93a1fddd059940ead7f55153908efe34e40eac06830445e6b2690f64a48ed04b75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5000c8f6167554631e90aa5a914646a60beb65ecd45c42f2a13c2317f4eb88c03de252bfbdb9e155b7e3e10a9147e38c655d07349225c1b2190979f7e290ff997506;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188ef1991c3752f107cb316d2cc114bed50f0f975baeee8d9929aa2e8ff1978bab029dcd8ba5c3f03356b74fa13ef1ed81706e920ae4035c10831addeee2137418256;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab6174e67fda7348b479468387b2ce62372e16dbb59e50c8d8f6cf007ad3c0e8d82f53e272bd8a8963e3e02e51d55377f5485e26ca614ba005391eaacae3c08305cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18acc19e6366d44835bfd88887f12490657f23339c236f2a11aebd0060119a68361a7b16f499a71d188f6bbc5fa02ac902599afe9be2851c6d7d6ca821dc6448dd37f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21aec40ffa606d62841efc3e580fbf6f691af0f27eaeb11593ff4f3f9f394e917b6b7ab3de81e9b47e960d3033c9b1dd899d5c9fb520b6fb62b6fcbdc7d2f4d64239;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1239765405d1ce92d7e6ad9b59be86894c480ac207cda05c1072ce2685c23595298b9fe78a5331820849126d3638d9d50e5b2f22d120f1ae15d2005aec91f065e31f2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h157bc891a0ff09b807bbdde89fd6c2482f7b5b4c465b803e6928fb38796cd05802d69633ad3eeaf49e1707033e3b629174541e759e3821066266b80cda1214f0d978e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8a4fe55574109141c9093209ac2cf89fed374878f10e8293da418f8aaebf10d0c0a5c2aeacc26c2b786d120cb280502adf0d5846912b06b3f43e44e38db47d678e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161fc788ee6f53e19f9f14f74d158266cf377c3191f7cdf60bfab20ba4502a22c5f08634247bbbedeb4341b6730dc0bbdc38fb6f1fb7f9c771b4a3200f35a8d68ca75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ceabaab6422da5e3ccd3d321a4b4934bbb884192e1279b8d57f232c2cb459cefb32d1b2851e03ee61eddaf1b3a5c7261e096b93cbb4cf229ea073dce659739f1fa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f07491ef943c1b4fb4957d0d631107770a4c22b90215544fcb708b6abaf0a39f6b9eb9dea18d84d7646a4bee7cf3d436932713cea729f36af50ed54524fe30dcee9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbded16ea38d223efe440497787d3325932965baf8820b9dcc304e4c07757cf8a39594dfabcc3fa7de1fb9923bb068ea96fa9b88fb6b95a0244ab784571c3872ba3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cdb21b6b24165dd3fb1709f90abb347a114392ee5042ddeb08e30ffa88cc148368d0c710624d9174c37d115e602c9ac607f7a445847de128f4dde6c35cb06decd3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7e6886c68d1df8fa4d1a3f31e23f9197fdac845ccdeaf794dcac0785ae8ee19e4678cb0203eb280659f35d299c565e3674a30c1bdc533e44cda23a543bb4c8fa881;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9396fccb6da0d6c6d1ece5ca5824e7f3793c4c4ece39a8bbe6b4290d5106ae91c158dfb1797f771f04d041e0cfb95ad710e1643e417ba6ebab917ed191da8f8ed8a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108b8ca04d847944763e71f6d0dd2ac3f5c96e46109ca6861b340b78af820d74d0f8b8767d03cc136f192155a3dedb491ad9fb9f716105b8f05933494e6e5baa959c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9d0ff61077e826a009787dc12f3456ed6506b5752c794959381459ac91b227c45873e48dc6bde7cfd7d24dd48264d213304d9a847322bce29dac8bf67e616445607;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b1bcead455ec22789118fed74a8fea38213acb83259975d1c22c44e02d6e49a12f33408833aec3a2d67cb8a6d98f79cd4c5c5b4e0ceb95b5d71fd2c08bf1cfac364;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34ccedc0bab270a0ca0ada7dc838f7ce5b118b728ab2180735f5fd197b8802c9ba07766648ce94a42303c459be02bdbb0bf3c17e384d4736eb3b1caf70f14a2220e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143282dc58ab9ef55ed117938cff0ecdef11e2b647a3a39f7546e9afa583dee5a42330d00eeaa0ba6231c6113398a158057e1c326ea41d91f4ddb44e2a57430d2826e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7816bba7ae0276f85165ee81cc78989abe36917985130a47e081f428acb1aa06a2c51240fa61d1d830125ffd3d5629e9936b82491b8bdde419a76280b46f08f9feb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1526b95f5a16fd739615b3e14bc4ccf0ab1afbf9b040967fe4bc0732ab8465305ca7fdd7476baa842fe8c9ba394354194d8844b49c1a9f43f8fd3d06177e68d9ed801;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd06fb00d7fe42a1e51b48a4dc6ffcf1f9cb1eb6aee97804348dc0303345aeb4e48f7f4dc2757f30023c93d43fa54b8a59c871de4d6b1f8564d3472e43d65e5e524f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f903cf0968c7fbb11b189ef4bc7ede419671e72266051ca48db5e35804ec0adab97ec3dc0562eb93d7144234837f88685c92b150ec413381b9d4a13ed4732f10bd0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167e3f0e52b57e1d2c34d557e587546eae85ba4f9eb59183ece63b6452e28dbd576cf113149dbf818928dca64161cea67309fca45248315dd1319d11c2f10d203078b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2beb02d49506826b6fe9db9d385d4badad287b0e9acdf774c20cfa12fd7dc6f0c9aa24a8e06f9b144e5e76e9e57da9635d4331d36a8a33f29342328f313fbd046444;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a75e0d1963f09ed2b295a0ea4cc384c654cdd003386f709f58995c6b8d87d27d0bfadc9a2c189580888ac18877967c80e17fa992a68ed88a60b717c7533d99547ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5c8eb37d12e1e829d1df1e13f650d4777d196c97e10e7bd6e5c7d335f0e6c2b6e3a438f68cb2db058a2b90f1a762ed123d0855e146279213d06f16b597f2115e40f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd773cfcc2fcfe8b2ca7ab90f1106d10cebb28feb59397398f97b7d85a9e1b4f5e38db988f73b03c7a65231ed26c6ffab81e6fc7dfafcf6d17c4ff851cb55fe37f0cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a64701d9deda6e5cd32c0ec8955cbe4ab104ececd71a084c70dda261831874902773fc8be166750bfb00324170b3e6a2a2a02cec41f11c3b6607204ac438b2d4da26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d8821e50c479f3a3860c3df90f896c839c9bca98d403b4d908a24e965afb66bd7dc343b023b6d55111871e22455caf509a5cfe4aaaa3e2252972aec92d7537d1c37;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18856c8d00921ce061574b9262ea59cc6e9493c61b992466d408a1810ba4a85ef11dda03b0bdfe4b3c5eb2110c4ffc22a4e7b6bfbb489edc4f139ae1de6c72eb96ec5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57cde8e9140a39d59170737b9dbcdc4b39ac708d050da55ad366197e93ced817098fdaa0b882acbdcd17618ef372b5bdb9602b4f4e7048c3df6c0606a5973fccff0d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187f976379152dfd432fa47c4bc6157f043d29343f351f7b2edda2dd7b38954e771191dc4d2360e447fbb8b22c8edc46062b135f58284829bdc34ca9d3892aa722236;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h507104a65ef1b37fc27ecbec3bf1b2f339acccfbba6776c1c3f93429a87368756aa078296680be60e39bf7042bec1a93f11a93c5373de2d3946ebfbd9a54bc998f12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fdc371f7243efe05ad857617373c5cb94a3fe82f717cb9c5fe202b0342b01ef777b9c444ee29fb365f778ed7bab3a04df59515ab68d70072aabaf3b97d4a4cf98fc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb92f4fdd5b71d08318d1b49a5dd0259931a2fd159d26a470422510a6bfd0b2e1bd27e714b3592d3c3cc102fb17a2e7b67a697d17ab61de04806cd8fba2151fbb836;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fd519a195c5989e3f39e24102c3ffde1c0292d102846dde78357658bc8cc9cb6e40a081a9cff43449a6d481808436043d002f1585f4df8a6a1f3516c7a8b4c9e09c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a970f2136fe373509daf060fa2c757f0f521641939d008aa2f39b3219167dfe8ac2fb11d8c44134a9272f9394bc3ef56b526e20af4568b0b74709be124cd1f93cf74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9cca9434e1398fdfc903627d9b2865419e2c0b762076d59a37d851010ad3056711738d5b3e0023e3f58e3537f43f4747496f4bbd32c00b49d74f76020f8e08dfede7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47745d25e701b4e15f7dc9577098900977c28829d812922ea5e5685c86012fc1f401aad5d4064eb07e13418d43febdd9e0c42fe7e119c48bc1618d8fe8a112e8a009;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cd3b2a25f80b8c583392ce27c3c98f989c0ee2a47d36048b1c716f499842f3a5856279f0a76fad99b23962655ffb47844461d88da73597f33ec671236d701628587;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19799245667998fb42f07a4d49f9bfa1b573234218a04f55549228fda2fd371fe70578066b4d4f7ddb80d15d6141e5030d6812c2e7f93cef280e791c52d5e2ca9791a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1885cb9f8aef3c278372a1eeb0459c62487e2afea32282dade4e064b2fad38712cc47843daacb036eff9dc8ba033c22705d281829340eb1f2a9cfbcb3e1f33cb0b463;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b1e52c85abfc024740b044aa58ea5328acf89012cc202521f2a26c23efce84c69c819c2c890ee527f8b983fe319be67ffb0fd6dafcd73b72c177ba0b4b5dbb7fce7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28929e3ede796273afb3db7b6a435495c6a1059cace13d068a38b33152f9ff8635ddc9f523e84ed4fc2ba64829d214460c9f89eb6dc0d339fb4ba136b744e57fd41a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed6ad3a811734732173e0ab9c4bf76ed117b68cf839b19102bcb404433ebe3aca90254e4faef10b55b317aa08e6b30ef290d4d38820e334686d4efb7049efc1ce7d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a378e5c417516e4109334ac5a3e75ba700057b824a108297c2c58aedd81ebdba8d1d08458010f74effdfde89636b2921776d90f3788b5686edd2aa61f1ece08967e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1cb0ba08987d1d989a2b5955777765553f8e7ed8e0213b50fd90ea6e973cf931f51dc25f38ab570b1af153a5a8cb9b756a267c5a5366800c0cff287d99e1c7ac20c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da9d0a2a2e049af5f9823a3c7ca411e3b2480810ae136239eb14593014ef3bf91b4a2163a7f80f29793c0ccc4fee8dffb20ffb1b8f50e14f75d357b009d74d218d6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b056287514b13335fdcdff054c015a624c5e1ebbd858bc5f25d8c231a214e3da5de2066a2e960fe33d0bd196efa25f20ef064a3d997fc477f040db8dae1ae0311d92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha756e1a5f76d539899ae42a1f821de6df3fbc487e850d5d676dc044a493e7f97a1ea212e0592352d22239725b98284e9c8587d4ad20ec0cb802c34b18e2ae91d2074;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1252b61968c491f73db5e1a0684da516453d0f56e642b73de7cf9551596ccd3cf6c94f395e44f7dda6afef60d4d9c5ef0ddff0c358a7105c9fd76fe244c8a66c6d53a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd665a78c3153f39a1956f3c813dc7160d30e22bb7752d33ddf6b718e6504a28fed854a1db9c55b92a0d111852cc2231df5f6d301f6905bdb151a91f131950bad887;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199b9998ba210026cf90e69ee52aa69804a872b250c98df1095e8e348c384840ba9d0288e45400e46f892fc50fdd664c3d13c3f829fe96af8b7b07ebb3e1e9557e80e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a997593996127266f062a7b62f5980f59b6014662003a3d45d8fd3d7db52a125d49e9b7e1b698995a2bf2ed367c39f586ec41aed5da3514bda4e030989d697a6121;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ba8dde9c54a5b2557e70781760643977ee5ad727133ee4fb8c96df4af89f8e04624ec83f4737447cdeafb7968ab559229641f705e90dac6d846942e976a35bb0bb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec49484255fdd7be8daf4d8db6a74c5afa504213cb48e58534a73cf9321f5748152395fb2916d9589128c0f3fcf7166849072975204320a8886f4efaa083d6c59635;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99eeaa70f2acab4d21de8c63a922643fc0ddfa428ec7cbe8d8efb1ec259194d64577a0cd27904013457c7d4b13ef5696e12cbc2436a8184fec34a10f82d9b65b9bd4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef26f9c3a1709d38a7821c87b352ad791cba9f6627f2279bb6ce5f01f46fcdf74d0b394e80308757afedfaf45b5201413f49b3c43dee12fd3e113344fcc3f05cc50e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4774047c43662b58af77fb7019632088cf3d7bbd7d06b961749fe8e9c93c284060e13ab89e94d6c8dd07869d7f20d9d71a687848ee8907d8ced83e74e843d02d18cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6dca746603f98b5dbac5773dd5f49f1aaf257c95bf64b1d7baf8070cbb6d2c221eeec6d916f9cbcb3deece5fb1c5a551b13004c35fcbac30e8a9235434272f8de20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148b9dd8164491ae39477074bf91df8e45809b3b5d2c4457b52479ff385764561548d72be5fccf746977052944302a96b6daad7dcaf430e2c5c4eda0fc2bf81502d16;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56270455bd99001610d5aa24beba2057d4f0047befbb505f78574e9d40a136589e6d64804a4703fd147edec834b27f01cec4c282c025fe0e128ae2e3b4d9bd4329a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15eb4326f783b410b85953d33b1ab0ba8b27f7dcf79caa2062882613d5c18460e03870b03165f8b0f902b13aa76da8c2badfcfaa81d7317428496b961cefd28388ac3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdf9d5347d742b1a0cbf69f874e62a50aca13c5f2fbd083f26de8d475185dbd17f84ee8ab213d80da0bb5aa6a7fbaefb2ded7918474f8c277f25f222a2aeee46347;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdaeb026f3faf9595af083a1db9ea7d28ae1181fa60fd66c8e6c69679b2b39b582b7b2fc9f2700aca82ec9661023e0ba0b90222d80eee2b7760346cf029b7b3c2e2b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf30a1ec5a5eff0382a7ac1d4ad9faed1875123987ed3738753679c6f0a73a7996debcb4fae01feea8d9c71c8b50fd33385a407887a9ea5e7eda0feaef7e8941d92b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc89f36eb46da0d3c106c9668883f1868549193f9a879c4fd46d67a6deb5575a8dee47bd32ad3cef21ae30b6dc2cdd04e045e3c8b1afe1466bf82cc5564c9995a6b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110172f288add343825fb40a61d9a3d8d182df70561e2b91906c67c8c74dad4a7593cd09f106f236475184f258547b28af1eb9226e10df49c57677447f319d3def94a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127b24116337e394e028d28395d0a941c35c940cc857249fa6ff6474a32711e94532bd713516a79f8181621244c488709e6e5e19675ca1e845eaaf1f7ac584818797c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd23d1643bc3b3c57d55700e0a861f9164b2d9df0be2a94a96d73cf48c734377fe39f136916165da30fa1f47a0cc1bbb5723fb5e7ade0e53af466287751af77126a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102eb5a14ca8dc506e1d18fdbd93cd58e10e386ca33a82fdaeb0ed3b898d09ced9d4fb6a6e5d60fcf2e51755b76103bda098dc0e46f356fba262e7a868c0126f5a157;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7693db8cb9117ac5b1844d4faa8b5ca1392f11b28f3f0c97dfb6b8701086aa86ede88231e3b959ef53c94778b2a1fa5843cc9a814b2a2f1515e0912e7feb183b4c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29fbff57af7f7e98906f0bb472503fbbd0bf0618d49583d66f28a2142c229d8429fc75ba1258967fd26b44346755a1f6c8158860545b84c3f047072a8f6d13baf8cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h711481d9cde5e8a6e86e4108bbfb27950892742bdc0c69714e032d7e0f09d0cf201c9a5a3c038ffb78b87bed79e0283ca88f205d7405f230153d53e427f7f46f32af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11890e0bc55a77277e052ad71abb773cb12ec8495c0550d7c7b44818d52fddbc5b01785186f22cdae6f9c83afd561b1b95a078ee05442e897c9435424e18db72a4727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebbf19b6e5c65ddf6d61989102ba57e447998bc9f3c57e1c6b47e7bfaaf921a568e85db6b760b4a177e1e01ca4df0f89dae362eb18649f7dda8515084d7d245b9d3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1330f8a544378ba07cb2c7270293558cf37a5a1259896def18f2dd733b4c1d089baf6b6506c5cce49ee51f43a571bf0e4669da0a73da1d0ea4e3cab03e4ef8a042c06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he314b63563c791968737d4733cea34be4d71db942f785788e11b9f767ff6f42158800a5b584930f4d06e246fe9f56db2bfa8a41690952ca0396c638c17fe20d0fe1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16747c8937f93ecf0c58577d77d38820aaea71766aa302402b0368a42748a73a1447887e18b6168dbfd7b8910b8be7b3619ebb850283e5a5a5ebcbcc728c03da104f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da36d5d203d9055c99b4cf8875007f1c0a1428053896a4697281c45a5a2947f80f5069681fab88040d2474db2ca9337cffb9116b2289315683de43a4bdab1e47edf6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb840700b494aa5d744fea36051661e8276d5b6808c0d7200beecfc1e12c5ba6b99f16ad4da939471c902d4de31678db1a77456101f0f6ba1d289c3a056b1bc900f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87437a8e915372197a4252f660bf82b713e71dfce5039cacd155a31b35e3c7c60aa97abe60ddaedc05521c2391212dcf47eaac244d8ecfa8d09c7c9bba2eeeae75ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bf8178ae86bfc115dd0013664855dd14bb6366e19fa5a6619ca91450e80b8553a6eb9f9d5d1eceb582304df864424eb21e56456200e1777f6e6ec84ea4b6eb6954e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5c98a866710622e27435c4cd04d18d0decb45dee8da5dfbbde0d4cb3c7bb296696c3beeb640ad6900c01ef079c9c921ceca93d80b9ff0f1db7fc56cf84621c3ba2f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f95c91309693601df86a0f9bdf64f23388c762e4c810ab8e6ac45d1c4a2de8dcf3f120e90249577ccea8fff722eded9f8b28eee2dd1b9fac4e8ed15f77fcf87f71c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5efc7c0d4e3d0a5d0f2027f6191421d460ad3e93a960fe261025f479af19ee4e115cd794d469e81bbcb7b1cec868c523578a17f97bcc89c39252b1fd5564bc1258e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f10974ffd4c3965de26bcab569051499ce0932d533cb6d14edb9da64c63a959e464262c712983af2fe59ba586d66adfbae1f425a1bb1ff4ddce562ff3e7c1387151;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc92311f1ba45476cc33f2fab2cad577899e15d001fa2c3914ff581d2b83d5b4bfd5fceb9c7993b9fb650b93edabaf15a3ccee23566eea296573255866a8849fbd60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1045d32bb0ec881d1ce631915072d46d41c9431d5468aa7318fb94696b4bb24ac4d85e9c652d5dd54679b5c1937ee495c34bcbb719171e71602c422ebedcd2126659f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c43737c4973bf3c55323f9e9aa87ea7c8a92a60b457fe0f4689150d8a5c3fbc3d06412acb22572b7f02e3980bafe7a0e91a6e9db80ddf5958efaf18d253bb3d6c3c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c682e414a4e6fde18894216ba1d97abbfe20696c75f6996b5fd1177f91fbed61451a2cdcda868e2b365cfcc0eb0a53e3b50da13dc44d9f67832b9b6523e463e42780;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ce67ecc806db9c46b3f257a70b41aa4559be62b835e73d22d131be2fa794e3f32a5c82c377dabcc9754e96cdae793d8aeff1e7c8fe756edf57461611e7ab4a3a59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h308098a5095368363b23bb105a3300da1d5d63f1aa36e4df9b20798643b80209512c9906d58a4a1c91024982d8c50448a7a9a5430922d0ab881dd40e593591944cc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heec5695e71eea1a0e5adfd593c260c35528d2a2a1cba2c4a3fc01399db093b0cdc90814d83784497a5502f20a285aab26ddc4c8001bd421dcaeadfc3b748390b8596;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde9af27727018bbdb9710faa30aa239957132077ef4bc1a2f2065e4d5339aff8524af9d95743952238f718a9eb7a174083c13fdd06ba453374b3dc243c4c1612802a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf14d457081c8753d34b013949d8098e807e28b6b50d48ea4493ecfbaf478901e3b17a3529de18083200f10a18649b23dad8bc4b92a6402440c5d1e02675d14c50583;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bf5affd44dc6d34e8b3b9a567fb552659b01980de98a84257f296559356add643b98b3e6b5091e5e9ea994538ce941cf8893c79902e062b3bfac68758597f4c889e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f22bdde87d4f0cf3f7de06fccd5b13b7ca33ad5ddaaf053d24775fe68e959b3a6270f360ab48ede37e32e4badf29fb94f250617ad96d8c9d0201dcced4dd7617628;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h605a23a77b03097f89ed095b4224221b732764319057315d5b344b74580fa1b19851b1fb48c196f01f3d724400307a79b0ab463dae222ab9f70a86137bc50c62f556;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd253591cf0e1b49b6611e8707f1284cfae08b774dffd826380545865b2f78e70fdd5f3541165a304699ec4bd531d55319dc8a45044c1bbbec07e64d50d9c0cddf330;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17478395165467426e0cc1c8a59ac614a3a0380519dfc1d840ec23bea81504e04593f905c06ca0a186a94f7ee7a9d9523dd31ae89f4144c07f7507f4c095595d6855a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cde5ef49dd0bae8e8aef0e33855f32dcd041ccdeb029d0aa5170dabeb3f2842611bc1f5dcc81ff49a06c6dd830f4ffc2f96209a817a72526c84313a031e8061b261;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6be381baf50c8c35cb66df06dfe2e7d7b1b3cb8e19719324e5625e901d958e747e9ee519d15ce6ddd9626c74f80448b5b5fabe026d3ee6e11f4725f5d73ab2ba87c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c92b00d6b619a71f20abcb53d95f61103b26df5d672479db381b30a64854d2f5aa768c327f1418c35fe0920369a114059c477e8536c5f09202e9711ac01f19257fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf02324e6d9661e8f813c00f557e9fa54f14be1aee4090d12c11ba18551b34bd9345779b79242debaf68831f9aa0452d193a2b0b752032a7f0118f6e91c241e772ddf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1270788fb7a833169150d015e4c83055e97d8fb89959078797a1375f20afc35db138064465b257c4b3a3cf168bd8c41fccc18ea05d008fe461d2ec5dd28cb227f3007;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3925481bb2c5cb588968e47c9c79762b4e344487ef0d4623dbcdb02ec70a35dcd798f7ee461ad8713a5e604c835a6162772d8a8532fa4ff332a0ea01ea672e908659;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha68f5cbac86231f749bc436c4921733f99856c0f7477c36d7b74111ef7f37944bb8e42b686c6e8b48bb5157550c3e506bb49ddb998926cad763ffd4a9061a684a74c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14842b81bdb67bd683912d34241b2ea7e9ca7ce31cf23d9077a2db30b9cb7b7cc896182f87df10e408d4aa3184873b0babb05ea10483d44f12f91bb1e55aa12dde3eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ba529678abcb68e295044bb0aefec92352354121e46f0f24e64bc9854b09118ff08373630a5b7ec31894261add5dc79a773527187245d7dccc71a4140d87c750115;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0fa1ecf304cbe426a7212e6ed0e6ff1d23d683a9e366482436c1519cc914fe9928bd2acee5eee738125382563d2dfc18d8bdf5916c21b577d13d7dcf4c1da37c781;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b9efc19219cd5bb3360fadb5da65cb3a2e8b7be758b04ce96e4c08dbefe642f6c048832fee3c5d9b9e44b698a92a3d7885eef2891e3e1150f2f284130f30b1fe420;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d4b964f1dea00569b74a8d5fd3d1861039173d0b5b12acd035bec7929cff197d1c1434a5fb4c9c43b033f32a7133b41b3af88e6e86cd148e6472a4aabc7428ec74f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1027dfa0c8d319aad797d5c8e35597460790cfca025f588ad62f729c03f0a364c5785b2ffba5f86fdee3046f5ea8dc547286dc2fd2fd8fd8e1371347649b11a562be7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb8bc0ebd637e5310f8a28f021d12515622255dc635d4666e799d2b9cf5dd13a1613a29c15af9f2a6bd333076624cde1cc478516fd0d56460f0761d2e6c81a589edc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h291eda0d2a4e91495f9b56576d755abdd621289247f7c065a591b5f23663ffcdc6a0ed7a51dacaada88d73eee844e83fac4a779c465f5105322c8297565ef66ffcba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148f48d3aae1bddb5a9c35a3f4379976e3a8112555fb24efd5f0bc4ec654dbe1aa49ebfab29de70ad43821f5d3285b4c9f40e8ca4875103239b885bc99cf0958f2045;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7303f0e645c453807eba7ec5355c90ced8cc0667192a93dc2436484a734b9e365025caf4438cb3ff4f1ab695d692256257c05f7668cb4aad3f3ac140b5eea93b4ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19614da52c756479fe8a1d99adf8566b95eb2bf387139f288c7e3c9ed223b86487ac4ef4412b0ca9679c4686407687b97337548963866cdc8e75af7571f1f530e18c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13548af65916e27711beff4981ece1fdb3a44554679446835897a9e7d7e14a755e0b439cf57305d6a231325258683f60b4191d294dfdca03cfbf51308340dc8a30814;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1641f2980f08811da1ea40e66ed6bb702f870bcd6351b7e0d3201f9325b8e1209954f7596960c3f30ac0e9241d947a23fd511bfe480ef262a0b65a6b29f485c61e8f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40ca244a762b5c91f8081af19edf3c7862339b4ddeb74635c0c2ad065bfe880fc7ce7d16eb761b5868ac446cf0617580f597f83f6f4aeef23a9f6b8285530f3b363;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a341313c4fb3a3b9af39672cf9507d27b47524275989fb807f3a245122cc5758233aeac8d407e8c4111b64ea138164e83c9aa522c5ce582f8b5f6bf438510e4acbc4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36b0f1927004ec22883c5489cf884f46cefe49f4f8f6c5415ed671698753460c56895962fb6e73836c40963d2dbfbdfa47fd936ced07001c0322d03f6714e3b70c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7d68f6e55ebdd36e0bd2216b4f7da77f453c66463d239e679514fa11997373dd27eb23deae87647fa1b2300d342794d08acca4fe9d2ee1e0713a0365b010e07f02a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12015bf8970779de0176017f2bb061e2e30b8ef326ab4e74af4a8fe7f1d5e61ce8e209895bf76645bab95a971c819d80886eb16cf4d2b1516cbfe89c0bffb8fe52705;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34f4770bab2f043c152b06f125c60e79b34fa2f70a5b3b03c056d5564fa007caa6398165696097de298aedefee037dad545fe314e30ef41d197f60754fc5fde3fa82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfebb1c1f13ca30f3e5602166af38a1b8129a0c1a6de579bc87a39c26ce623360f3f553b380cd2c48949347876cee02d9b4c86de37e56d0a1952264235f4598365076;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb7e2b150baa28e6129f7ecf7ebd89e367bd5e724e5fb526a8a696b2a74faa104fcce38f870513edff6fba9e284ddb2a74e77fdb041f37a5fbf0f206b5cf319cc8cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h328b42dc501dd00fff694c3c0acd415317fb6dc183df56503fa049970a082c10bf3a0af30d24d5612f338eb14cab8355a3ea030c9d292ae7aa30eef9f629b13268d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13beb4d8fe9f52513bf51cf5dd0caf5032faefdcbb32a6f488b438b74f1689dd5d6d30f7e6a47a7027afb9b4fb978bc0489e96a347567a856f3b2584a72bc598c419e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb33757df71932ea196c265e20e2205628699d0f67c11d4bc0cb6374d2110555fb55f4a3311d6063a7be3e451ed1e09afeadd8cc3920248ed010d777fb91d51e22cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37ed911ee2e193ce47eec4ddc666b7c9a5ef9c2dab2d254161efa7fb317397302395c180c0ecc081b12f7030b5b543d8132dfa8a2a017e5dd787abc872bed40ac385;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87e014af30d0456ee9244df7c31a2acb6993e71bed6bf54cf4be6193116374605e2612653b23eac605695afb12af1d0d8dcc3c57405652df483a0227c6963b8c7a07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1541654687b046553783512dc7655cf7e0554b51533fc7d84498b94f90d3d0c2c13c548639964c5e5aeffa858e2ef13d14e2aa54f22fde4524ab0f8e88ad42de95744;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0f895546e3bbcaaaf59ca373aa9fb63ec6edc7f29d17b031548713d3bff9a047548516bc8820a60b2d852073d64dda1fd5c245adb0884f77ca5737c5442bf4d24d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c54e35c897e143ee8e79d968f555a3a20ae9d734266b08f085a40feb3b561a52a40f1cf30b354270bf6ca650ec597dcbe159c92b39003756bcf33aed90fc894360b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9bfdca982bc8b67e15f7d314115c2315a91091f82de4bd7ffb35f7d7c6652342968c1bc1a891236b7aec6d439892c76db8ddcfc8983988b9262b36f450535d72c8aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198d856b391a0123de1e13f388e7a47fb17ace6aed5173fb4b2343ef62523d1d201737128e6541e1683e9ae62dbea7d3379631714b52d777f284f59f9b4c52be289c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb728bdb3e6830a890b4115674e0453091e257f251d35b11fb97f459845d9a459a081485fe6606da3c63e10d536046f93ed5f979b17086ad333cb859c295341eb0aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h863d9cc3eb4d91ddd9095f97178dda6eb782ccbd44a2513f12d8ce215e8d030c359f16f3f7aca40d55cb8c68b255adbaf4ebbf8c4c284c12362821c4faef314378ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cddf97351e76ba11e9b0a3a88850b4731608ae724afac89023714eaca9596f2c2296e7ca43ea9dba31b23253a749146209554b4fd91371b662a6e6d3c53d2c2dcc5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48e22bc447a60ba3fe2712fb7494902b219e28077b830a73cf24d9d09af845d640f32253970b9a9c25a7e9d024119fd5d3502ab2bfda8db1c76a8026ad209c84d4c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2037ebc0bd1c821e98241b9ae38e643a975b9d1b10f3b086d9f39a3fee945a4eaa004c581a3aff3379268b4c07389c4705c03db252fdba2fd9ee391b07ae214d77aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1118b31e49c5e0080b7ee49e68cada26d820b099a89b05c4835122440937ca088e8e4bfe288ccb6f844f36546edffa8f4c16bb0f28b76007d24cda5eaef08ddc7138f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f4f1304a632ed46aef0feae819550d7622d884c06539e923e0ea218567a836efe371e070c06b4aebeecc891d66b7f87719e12db14c42205e4d5c8098a94210b0393;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16241bde31179df69a5f414da5ec9658e925a210d0c15dd9a0eaa5841439676c5836b8fdec2ab3843931bd724bc95aae4fedebc8d672b06f2564bc73e865344c80603;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f6dd607ce681350008489a3df62e9f83ca05ff3f5a2f8c4883f3fecab967ea362519c6d853736e0649129f3e2e32ecd84ccdaefd7f578a49c86c593cb510b231ec5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187c121e36db72dffebfa77b8635d7d321a683d9cdc99720d0a1d19c364df9cca5f863136e2379a11495a8f67aa1db52f4b1d919b2f2aefd3844fe1dd99f9e5885592;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6e55f24c045592985e2114ce2f2c40026997545ec46910f4904d27c9534fd264bd846589f60b8a6aeffe6da9ba0a51bdd8e98fd57f6ace0b9378575a8c613a90166;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d168ddd3d0c3b75f202f0fd9c888acf7da0e068928ce320c87c07019a6c67e87a291609dd9918a0a001b96a7dd4331f581977d285193962765aac4ff1edebfbc53c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149e98958fd9c294bf38ab162dbbec9dd38cd77e54ac8f40d3e03b9f7300d49d5df2629ef126dd03a3df0bed3699c0d6acbe8e9aef38ba4a745192ca30fc163e01df8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfae4d9cc3e2b36bb72577048a9664c50604fcc5715f46ae036be12739c85d48fa2d48eba5e1a316dbfd4f50761a589af0b00e0960b409e575e0825a8c585332a9b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2eb931d2a70a652835e29b9aefecaa41ab825e42b946dfd072d238227343753443a7e72fdb09c6330af8e8dd9b757330c316693c70b59d417a481c3917006fa643a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd208d7441cd5e20eb481e7dc6c3f56d63d30510c05d2a99ab69b7d15367d2250064929b45f8192762538746d1cbb2b04ca031b5589c73d156b93e88ff3180077a07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e58602bf3f95fa6df2d0c6e5fffafcf4a0ecdfff7bfa86379bf439d3efd2fa5d7dff16206d78c21f533a42c8908f41b9d59cf11335ddfab9e170bc0c732f71dc192;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198c24cea27b55eff5a176476775fd413a7c359d0bce2694cc44961701713e6e3c07868fc73f71cffbe2dd8c23d8af12992cb1eba2d959d6f82c07f42ad956bce35bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9964ffcb4cabbac8c80d852944aca55cad5557208f1d0f5490e91bdd8c0b7714dd980cd65b2dda0e1c7d688aa71502ea598ff2365c8c26a2350b4addc45f8ef54514;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103cec03023c9f26e40d785871404fee7fda79b2ce4896a45dc5ee0eeabd586c0fa310cdd77eefff49e5b1e8832371ef47ea3f0315cf1240ca6ac62a57bf8edd1e04b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c30bf7eb1af17e1592590cacd055ad12aca9d1f4d3592e8747a8a2f4ec59814d0c44b75666e80d8fd422d1562ec301a9d3a695183c1ae49fe2a24c5d112717c1255a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1140d7199c943daaeb839d599cecbd10c2f0c35fd0280b60fb89871ba0550eedba917c75290a5c080423073f9a7cdbcce705fdd6de3171a8477907fe3977e1029e455;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ba94dec875f7af5a0ffcafb0d11d9f6fc367761e2ecf705ff6a681a1703b14b8cd3f32be8b2a11c624a2ff7ee0299e28cfa80cb27b97cbc1e33c33921bd85d8ddfc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb174a9d4cb0e6440de2e04092027cd167261fccc7de70d1f68594fd88d8a64cc432c31dda950ebc7be4cb8b20949318e26eff16a356abcc91e1a439dca207df3837b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d87785a07e0b83249a006b6141694b6c7714858aee22265eb3a15c9004f09866073be6c92d4930e89bef008c63a6471401d739c66dd3c8e2eefd639452f0075d83d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac3516e40dedd1c1991d1c5e4ada0de2b6d0de5b25c017e40079fffec8c56666dc24e8907dcad6b6e53732fad9b0689931882a4dc9c6d64f44f8a787b47eeea901c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hece069be7820599c3b9f6a79c2bed73853c864bc09c1cf9745aa611e71e60dac1b8fcce15a446e400dd5dd36b35278a8f8561a19540692e55a922ccb9107e998f95b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e98b040e70010d108ed5016d693c449335d801bdadb48c8f5b268ff6ac3176a38de07d1866a96062cfa73421781c4bf34aa15bc0055923a54dc1fa415e23e0c5c56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha09646ecfe316196b5d26a60de5b1a6d72a68e419d44617c1e1da61f22056b20516f008c0fb20c11b6e40db3885dfef93105f97004a2fe5df71e0fbf38d1dc248ca7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3223dd40221e43ee4c11bac0d4ebf1aec70d807bbd1dcd2a03a36b27509fd0f83aad4ef78990dcf759dfdc83841f4de5660a667ac90f98787b07ea8162f947e4ea8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9732720d920488127e9eb172d2e15875eebe5e57259fbe35dd3a5253a1eda00f6d1b988683bb4cb2ed8f179a943c598118c8b5584b1aa992b7646df47895b84e0491;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b735e51f333843108213946c0387b020a271df53ccf95c22169be6a9f3f7c9c0866c9206a2d0fbd153581d888dc828fe5e968d3c3694f8535ce92495e1384baf781;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h238c990e65c94aaf3c71d18ddb28704f1138402139cb073b837e265422e00e61b2f978b9ac24445867b1f885cf9fe6ebd61f0823ccdddb14f441729233b754c14a02;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h571c88426a262707881bf05bdd4dd3bae52cbc2e9295d971bac9f7b2d994235bdbe061ae9ef7fc4527ac0a6dc88674ffe0f899d72f473381c3b0017ce5e05fe50bda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6cd90687f00c2005d202d16d74185e20074b8fde2d5723fc2bc6f612536d13e86693439585dfb5f259303ff875a46a9ad548d995b795a23b7338c21ad68980dbc13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98ec05ff2ce213af291bc7be79c14ca4e0eca74b4009b842d0a183be0674a82c7fa0d371759c9b00aa14184bdfc7d6bfd9891460e7fa5ae3310dc580caa779e6b743;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eb2e644dbaf763d6635d7584a12c5122297136212f3a7d62d90821b76179fc1bd053d2ad70e43875bd157a5bc6fa2b0346327b23b5f2eea49feabaa7e09449e2b29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8313ddbf27b48a0b1180b92eba567763fbd8957bd6ebfa35ce7c6087f0e08b8bf5621c50860fb02cff9f8cc19ce88f0d300de0892178c0401de30b02e6d00b89b8c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109c895861942151cb337ba8518f01b3db1f30e9cad64b0e1f3f6e6e962f13116fefc175dbb7e030ac5eea62d4bd3f6eb61051f89ee3d22477100492140d8d9b5d18d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2affe4b1319ace212ad52679ac2b6853f5c4191d829ef3bd8700b0a410d4e3a0e8ed899846306ced23af8f3301242061901fb79655d8b7fa30bb5697db1baa0e07e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h752ad1acb754d146552b8af4343711994047df93f7553d8bad5643eca3d2819f02a6f98e8e100dc784bcd85a3acffddf7b954ab74535d91b8e74d7575f8ce3eee281;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10db06120077b855ad8afe7428e07d3526b99eb18f1f2732088f1c7636956f00c31263d0cf6470f4fdc4d3d604ef6606d7f486fdb79e39ec0bc82221a59759dacc16e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f505c17eaf4795c29b5b3c71ec25d69bff74a6d3c96723cc350a9512f1bda43029611f6cd590af7770cefa00b4158c970fef56c41bfda33044155d8a30ecbd80162;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e199bfbf62875461a5ebf697577578dd599316c5a54877698ec6097d072a009c3bf9870e50e64c84e356f72d5c28e4530667ef311f2c225b798b06f30b5ba8ead90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc17109badf9042b73cbff4a06659a058edebbf3740f71b0e67b113dbe7ec161e34f8560480e6b35a0f07ada1b01c0efcaf030e95f0b16f18ab715ca248f0613d8fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc3ac7e5c7d1fb859d292e4b5916c641037cd851d46d0fa74bcba4d7f67b55efb9b6c794f118cac61acc5822496487aef613a654d093f5eb8bb28851d6dc8913246a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee8f5eae52638192f7e9adcf66fbac5e955e785ec7a49c9271917e016e5fde27a676e43c1ae2adcc39e79236f72881eb57de4bdbd570ee6fcb9dd99191410a8760c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5894471e88a8725eda323bd162d47b11a188c5951dc684b4d18fc11e8126b9e5f8149e70674e7df4401a20b1d3fda61821f8775458b531f9dbab3d1244f2b783561e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41de008c551b534b70cd0ea8dcc76545acdcf507a170a9f28037d18b9e3c99f254273c4cc68001fa4fcebbcf6a5147967a2c1c9470b65612f3bc63768c9d57ce4d9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199fcad540f24de3fb46efa74661753783bfddbef06eccacde36af5b833f18f758a05ed70a5204cbcd36c4e16843d93f3a509edc178bfad2fc81380ff7ff714848489;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84c56f12c897cd51f1db9dda8566db43a454e1ef04ae44a2791fcce8e3784f77c270372bd25722f0428339a4588f6055affa43238df752dcb5c7e8dfea3eba792aa2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13893f15b8b675fb0d40ea07464f36f008cb25080ccf11083bcaa7474eaeb06906979270364429f01fe9d7eda40a433e4d02b6e58e3db55640080976cb6266d0f51ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74a25bdb1255f070c868577ce982f9a2f71cb7eccb55673282d4a0ed8de9ff21b2a12e968cec52cf4fee36696f2436634a01582b4d1e688de3dc48433ae8cb873226;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1462fe13005a3af0263407c4fd6c34818d9c73c57a444b23e619af93f0fe51df522367ef2712a4c860d03d2ce9009ec520e3615e0c88c218c2bb5dc9cb6cc61547b32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce2106b2e7f485942901a84001e9761eb65545e8660ecd83d7d45255e0554d7135cbdcea45ecc93978178e4c3bb74b64b0c4f5ef54d63b36b2d786a8368d2a5f1ae5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181cec86c040e0b31ba4a318938b522300210bbc3d73985e24d8eefd04eea6685bdc1263e2c66b13f3b793ef5b71d9f6c965f9f4401bae98269d58d52ec10f3679621;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d5a1ab9de9cf6f59362b37d975e265826ba52de166f4f8133cde40c0de719d35eeaaf71b1060741534df6fdc62c195e73586bdd4f616712dd4543e118709d397b5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd022537379db39f07c247cff776d0dbb8e1606d32f1bd48351278fe314799e445d7e97aa66d9264d602332c07ca8abd285762f723015dd3923504c244d94381a691e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88a50a1ec4610b9896cabac5b476212cb5746c9a7df4147b228df64123d5893c6e4944470252df11b07f6428685122ae3871a5dcf3e867551b5e0b749062d4d16cfa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdf876655a3974f1b2c9ef2840fe37410aed6764b5375fd70ecc93886ea0d973e27cdda44cdedb608df91d30a57885cf9b3a2a7f8aec59308ba9dd4b1e3de9a0ad71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f14d1552545a4f7f9a942d3bd1e73978f3d0cd6da8e3ba2e43963ba8ae06049a6b0c5ca1e9156398b936e44ce5b50c657f1c6dc0ad082174069f4733190e5e15fa1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee493f208972cd98019c1d20a031c04188c7ba0630284c69ec16fab11fbdcfd4b9173026ccd1a7cb7dc473b5e238319cedb5162b3dff010f48e1bb7b1126f09a5267;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183f71e7d9f241af56705e7ab6e0f66e8967bbd9df2b3c97abd514c74e89d27f8380cc0dd5b6542dd46f283347df3d01f1788259579f14bdba9a3f05ff15568bb00ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9672b5c8db23648a7cbfd01445bbd061ace171bd6d6b5f0e705eadc82a82a1b745cc95a37cfb9344992a627c04c229db64a80f914a3ab15c94cb87d74a42c16639ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14186d64345404d49d19a0b182d3115ba352bc82573c3b03c73e5156ac412389f95f776e0b76ef7d569979b26ce0749c3cd4e5fcc5beac4c1154c9047d2cf019e775d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc229daad2444fb5840330ef469a303a6622f39aeb2b041069bbb484fb0d744ab46a772004d29bc797bd49167ff853c6465edaee0191fb9960798ea728132771f27e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19bcad27b7c3b20ef13337bd4f7cf3f0b3b3fc007ab943d5007bf9425e4b565191404ab486d135e1cce399db8489a3a2f9cb713e7d4ca6f2ce276de4d1594220780f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42883851d4e9114f9f9f27e983b5d173a0ecac810377ebfb7c1a87e19a03d5a1262ef591aafc399c70968525c7fcde117fbd29a7831226dfa6995f3f5beee2ef6e4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138ed348c60fdae96287412eab503bf2f8b1492da8e3f6a7d09011c03110671ce169cd1d1c1e43e97eac1a34a84a1f7dd7989afd7ec24b201c5912784608dc5e2e10b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a15671058e92addcb2e6f07ce31d3b945c4bf4d0d143207d9e35e5a8e70dd6ea1586ec798861b017bbd6a242f2f77d80bf4751593eb468ccf5db31949ea36328930f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa180fa714894557c1c13363138f62c4e979170172676904b4af6228546a79ed70f5d7de912eb6a2e133f7203b68f4c4db77d44df55a7f231a9d575876637d016ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50ae37c0db7a07efabe05ceac957e3e3db28631382e87ec68ff504d99adf3bf33bfbcd77166f298f266f7b3cb16ac1c68338d894879911ebb2f7a606d6e894c40b7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19981cfc8cd9d088bff33461c17ec811b9439209d7387e4b20c09b64670b6be6d7da6ec5ad0eb856822d1479b970d978a0837a4d0f3a727b3b59c1e24f26ba6bc4287;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101d5b2819179135d5a73d7ee3f74909d32b4ec5b8049733163263bb6a42f8ca03221b268760aba81b309869e2c7dc60b2bf2531acb40b6626837327dbc49ef11e601;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac02d9a216351f46e7c32fbba330f13a8435035918711f459b483fec75b73de8d77306ec3fff2a614110afba87a4262d8e15390ed3f3c88a58ca486cd5b58a00613b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0a09df919b58a94de71cc4123aed8746ff2ff072cf26c22351a9cd24f53366aecb052c114930aab87d49017183460528d62a8dc027ac99803e22a4b0258177240df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16277920fa82612ea658aa818d43b7c4d209d77cf2af71477f1378f156c7b251f520482544e0d0a392ac8e46b684fe94baac1f770cf6658263bc1e66f9254ae1c48ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4a05bd0455e7c6a03399e99b2665910f861655f7dda327074828d685c0fc7c99294cb22f936ab81e9891a5d32c1d12ad7556fe6510aca74dba9d9d170f64d0e69f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9f73efc1faec55fa34d6e52bf5d1d9ceff978aa4da2098a1ed24f69e812954b740e7bd40a2edc8f4e3c5ae8a6b04a4069fed2a27fc0fa5f9d14444286a385b87c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf55980bca38950712cc7bb75e5fba97c9d5db517298e371c911b35f7942defa0878c7260200324821d52c909fd6050159783555ac486a33e4e72ea19fc5df192ceb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e0c10d2bf7f8dd644ca2f3c24e69bf65557796e267e1a4b5ac70f623383ff5421f7088fd9311ccb2e62c7f808f0fde549ddba770dd42a95e0f99ecdbd4419ca4a39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1198df431a6edf03dc24d898e9e1d97eb64e95ad8be58ed2d62dd55ff25eefb92d68e949c4acfd198bd3c5c0a7ddf4b648076f52a90f7fff2874937c74dd9a8ebd608;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165400df7a7fac6a93e717e09d923da9d5e7e2fb09761a110090fe7d74cb7a22a251d707a230ff67399376fd27bb2c1c4f2da2301c6280ddb0a31d7107743d18a6e7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed1156e566321bfb35a0de512f37efdcea3061c42d23562bed48e58a6e11ef33e5705a05acc53b2602f7ec3449e7f60504bebb829fa4e2125f138c364c3dfb1f0167;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ba6b0cd77a6fc153cbd801e6bade6c5e2072b34a3e55a3979bc3db9fc0e2611bbfec904fa5a3b6e75c6b849c0e851d24731eef5d6fc5e4d1b3cb64c69bdccb9eb43;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100def668e264f54d1631e9663ff7a675bd8b9d995b23e1dd733818c1f90abee224346a98fb8ff57845cc8189a121b4b784bc2e4ebcf45b6be43812b0d16e66f38cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9ff52fca70061e75a16bbb1dba97d57dffa969c0f06ad0b4d9c892004ae6c9a7fe0a2bb7e73dacd44d575a1755ff4e4aa1d98f4ea6588535398b38a89d23b21dfc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb5e4a6584ecc03ed70a5300971ec7aebe14389b999f66c3d3202509cdad30c172d8f00025dd30f7e04dac7814f2e5a91a1ea0da259720e8c3583ab7a2f835d3daa6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1460f201537e4ce7b9af290ef0d540f7565206180a8852045bc45605fc05876bdcc85f289dc1f8fdd07e72b62d673414bec5c5e92eb4c4116b6051b7eca37642bb757;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a220799faa1d3aea7e8582a279f2b7c11f5cc9467d19e4df894a0514a074ec5a5e092b4f16bdbaade3fe153ebba3f366ff31404dff309f6f7556c80bcb09f887373;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he27653493becb318802ada20436431400661e2a4448c37bda89b7ef4aa139757b0e15a97524d62fae409ddaf1fa25e20513d55e1f66f7377428729c49012941a4c47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h716c269b4e9d465e3a15efd0496c5d52ea4d5ec5f1e4a5962f67fa451ddd098fa9ab7b490aa7174cedc797ce202c386180dce8529e99ececa220d9b835ec2c146e43;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15742208f8b81c2a55f96306243bd7a3b266d93550df8af117c57faabd4e66e8ea8bb682ecfd37f3888b61d89b8780d118890969b6b439baa9a94c2e62117f98966e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5d242da460b196a99564cea3f8073d6203e54c8e9729b5417d35d8d8d9a1517def5fef959e99ae4ffecb9c6d0f43cf97b2734f2ae10eaf3251113ced305e4e7eb9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71f2a5ea59f62cf6001e662b67f70d27418b2b3b2fff3d95e4f7b24c8bb692c48955349d910bc1a53b42a87f17c95928b074f21b45e0a7778e3d92a7d293e3a904a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9bef25805eef4994878208f8720aeb6c53e073b9ee4c18d630d2ca9c16779418673e97fd233353df734822b4e02b0ecda9191bfc442414380c3a011010ddbb5436c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de024a05a124c79cc144d61559242489cce862954eeb69ca9e071335ddd83806870c52e1f24af0559bd4ef83e0c44b9b2c530fdefe8041bf568547c2a95e46999e2e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e6d1838470518c12c4f7a58c57afc7f0ff07e1e7c92041640414e7f74eb188aa42eb90b79e655d17074c98875ae716292ba25c398bddc011016a9da48a333be72ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf869f6d134c6ccdd7977d93e528d4903ce74dd63e3d48939e3c37294b8c72c16d635cc66bb8c8817df22ee4ade3e7af762751b187e78f42c95eaa24eba283d2f9ce9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46dfe07c0e10aa68c0ea798df4708bbb22f1d61a7d4d09750585db5f04469aac63234db473a37657cd0a43d128819c0ebd11d9b4a5e9004de3bd887c86afa8c259c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fdb4e22dacf4489407b8198ea27fe4029a20a373e5a789e567e6e61dcb3be539ef515935bf04e4e409bd4bae998d098a751d087bbdf1dfc368fd88bd5457a7a95a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f84be1e41edc69989e1cc98db0006a96249a12609851cd80deceac086b275cbef36e78ca3d2fc557f494130d4d087f31c321321803bd1247c56019cb997e0a90817;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h798efd869d2a6736ab3ce2ea036412213f95e13642296f37140c141a9095e452958a7c9fee896fdcc0c188f980e5d93c4bed9e8b45ea6fb46607150a7fed6abffb24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5667b02d01d05bb2275da736ba48cef568e60d84d505716d94ee27d62d510eaa83a96ba460961da7a79921575732e9177fdaa9a8d4da5ae18b61eba2aa074dc2f282;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180df3dd6348edc8f0a7bae482d8703f0b15f6e6444a9b643f7ce9153207209484b18e1818527cdfbe639c5e303abff2713c6b1dd37564e930596e4f360ce534e7b31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdc9688814f2872abf97c0590df83781d051514fff259726ab23ad189fa6d0d67f4a26339307682099394f19eb540088cca08f25b054833eb85b0949e9316982b318;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3cfcf064a4b69ab51292b7cae298df3a28c15fc70710d36fb708f2debdc94634c8d204856c8e94539c7387e4fae3e0c2d8df1b52daa4b50aafaf50bb1baced79146;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8bcb3a24760d7e28265282acd1f2c6ea84b9591b5ae06a8ea8ad5e6cc2ecceeaebae4fad60a1ee12268e7909e11e48eed4d2649e7dd10557dcd65139e3c03449edc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37946b24b7044b73526d4db8403af1a29ce87d1bb8f468a0b65eb3962d5ec340b3aaf90e31f8b2d0cbeb0a9a2918483e0a67c28152d5cec62917f260bd06c3719af2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a356b8f640c1edfc3735e82a7abc64d242135226943230093f9843c51bebc22df549631671d47af8b17bb28675f458e656a01c2b09941b6585e30f092c1055b63db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbbc3e0063a98124fed568b7fc904a23a3456708d7c78403d781f7ec6374cb3bc642df0154a9daa1e4c5d51e4ebf8f7af0b0675a48672db088e3e97e4bb2466437d07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93fe94677a3db7099ec20925a602657f099dfb55ba0d68105f1295d056faece73835c282590df880681bfba770f8732433050d37b379a290b73570b3d80475a6f470;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1febcd7cbc996bfc7e8706678eccd86e5443546dd0d39ded37af13ed86b4fdcbe27937569e4a8a724cd1548733c5a5fa02b6ceb6440ba1c56aefa5258a6493a9b4441;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbddad33cf8a0fdc8c49762c085b11ecebd903674c8432068dae34834c3b9747c338a197f59c31f331ee852ed6578db9c45dce872e82a889b99fba68922e14cea54a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f7c8ca3030de4aa4a3c8003eedf02e2fab152660f462ef67398c1a90f5caed5d1bb90d95e671400b4ecb20f592e146fc64e4be6c720de020ae3bd053c17086f22c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17caf4e64bc68ebc44269bb86942e2add9216a23deb55eb28c820d13cae0bd293d9a35b08ea83a1a42b4aecd2b4743c32d95b8a575ec2497458c811692e90fe6966a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143fa055c02f526da05614cdd14a392edd5d75cee306eb88ca78ce9fa4be154771c20f29e9d8d683e72bf51e84e9d1fff641e7379589af3705f5c9e7c05e10a68eab4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117343f645c15b6b6b2aea78dcb987e977e7f5aca4e20c93ff6d813133185ab99f1323eb7990b982db9087727b6cb1eb7a67d4f0bb9bf08d48ff868b6a7eee6ee8b0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1752296b57fcf98ee88db454458aa72283de7d6a791923b36c053558812cd5efbba91c23aa8e5ba58818e053e8d8b433613e67e465ef254d6c26f71dc89c1f71682e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habbd03ae946a353d5d1b83fcd3fe509013a82d82490852262134099306fc828ffa0a59a66f6754a904fd738965edc52957d36df4a70e047b5c87ce878c679bd28538;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8df1733a2c211775fa8085507c6ab84c9448f85b53f82960141928d768f519d1ba78f0c8df8fcbbbf82be975529762d12c42552c8cc95b49e7d6f1680b1c101806ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d9f9f74e43851adfcb3aa169ea990c254862f95d783ee8527a52fa55a767e9181d23078d2d06dfd7bd1b99b4183d5dceebc363caf16a63506f96c06da5a33d62483;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130d2a6f58813d2796a26f19b44d67e9ae4e35415c968326b54678b821bd43e5bb5f1919833783fd3da5275262754abf11538c24e61167a4a45139ec34ac560cdc162;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca4ff2abd162f812088769a3017e346033ec873aee5c24e57b0281197c03f48cc9af7a3e675e23ec463e6f22392bb7988ed9dfdb2c8f8b5faeef685e7335a4681a97;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b79d5a22153d47b34c396dfc889cde44b0faf11bf0fd47611c0254ca6f343ed7ce80593ad7c84193efbe4886b4ca0c1e032f39393578967f47b92b36b394a98a7753;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3973d8ae691bd4bd1fbd893d7c0ba81b23fc0d4047a19575cf73d965f604fef3317baffbba10c0cc5f9e408d33ebbee7609b4af26c85276d46ce23ce9b748014b28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cfbb8f89edcdfad67e5af997b563653406b2a338cfcd61fe69d060a10024f9bbba1c053c1e9176c3d14b024e83f0a95458d1f4fa369bd739b13f3179efecb7917ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110b5a09636ec60b365ae20ece3cf9568b3d6f2f10fcd89bf81dd710d64d1c74ec54fb47fec76bc3838b3aa30fa0b8af4bfed4bf552372a86c541231367fca6eb0880;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3265101fc083927d22c6489d9d0eeb3bea8b13956afe21ea639a15fe7da10958ade10a11662dd8072f5a0864fd6650b62fcd7ccaf0b0ae8266ffb04baa468e74e7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b6791f5cb4c1487d11b8fd1f8d78ccd3fdeec4fb9b7bff7db07b529ef13064765ff0ea58b661b0605897afc9ed4ba9e21ee9080b7ddba0d376369c11105e09c8435;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1f35fafd8782f8639b178eebcd717b5fdb005b1ee824d0e9adcb78bb16ce0f56c9b8101b62bdfbb0f2904295b4b4a95568566c1b50e652cd4e47ba038dadda9fe20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f61d75f26612b2ce221583ab6bf9b5ae67949db05cc32955653115eac6607ad86d68d36de3f4f052016b69f03f22aa5a1ed3176059c8fe23a4b0fc23b5b10f57305;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he26139b05b51742f0d476f9d159dac0633ba0984095efeaa90ae8f44ed88a629a8bf22d69124d8ef63c726398d57462f15214567e28fe1ede2aaf75e7b55952da743;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha36f53bf6f99a0de97f4e58e3f364733f11904f50a8040defaf47b664a96b1f47ad9e9ad57911b72be77da576e7bd0979481eba0344b1e09f65bd34c3de239851ae8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa39aad26f3ee67bc6527ebc9bd71765d73b4cb2f244f2f1c0bba6a3904c4ab57064b014246577c1d266f909b005ff5eae6a293bd144c652cf04ea81a91fce92f647;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5298aab55cc06ad7cf61e8a289e7885ccfa3159d8acaa26e1d210940ea7b3815d124cfda94b3eb423739e9a9a947eabfe9fdcaab613633d0fc9ca931d352a7f0700;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f13481ee67ab8c29072e9d9feb3968ce94688419987b79b18a5fa15d8e0fd92a602a5d664fcd1da49eb274801abcbaadf9422a2402c057fc50804336f5ed3ba85a0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h654e43c5ac10552a6e290915414f41b85df0b93666c1dacbf6725448c7581cf43840ac78a3dab6b417bddd5a71c1fa2dfe01ae8fcd2c3f2f899b6c1202b14cf2088b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h781ef82dd564f59f98c1d7d493e2959e767b3501f858f33391293d03887dbac73a29bfe7222b27926b0abd1c381810fe68795f2c15752345ef88965442eb6c0bd424;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae5edc962bbf68a6ff5d4954d9d923a5c54f12b819a6c9e1cc474b7a1b4bea985c5fb35b8b24ee52a00b184405da662e19714b69d62d69bd9c3a546992352f5c0127;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8b8a5029756fcab185b4fedc5e5fc1527e15163fa7717508c87e5c9754d407ee8bd22a9556b120052a027a3e92f8da71aa806824c42323f111ebb0094f78a58c3c26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114ae72cc2068645d75cf43e58bfabccac0ce7254962defff7a83ddfd5ff21bdcfedd45a49815424744584e9bf5445b6151a7682469745ab0796ed2096211dc123e6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff6ae2566792d965125f0c52c2e216c9d4c899e7cc490013769c61107988e049cb0e3a0187978847d9feb3399b1d042da223154112d540bd2aed169cfd67fe442c74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habf61f7f02275e5e2d2f4c1cf1036a7af2532a30b31b333ce7794ca890c67bf3cf2dd1bcbf6429aadead48ce70985009a512c6b0abdffea68e96fafe05640f889cb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d1b584c239df169ba937f8d9f568dc89ff7f25b68f715dcadc1fe7b7dd7d677cdc8efe8c71a984ec578f4135462d91d16bfab4f248be2c027d195125fd1a5602089;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hecf0c5ec899fb2219cb2cd585b0bfd123e7505cb119cf50da8daac761053cb104eaefbad1539da3e0c02f6c3399ffb94f56049a7e10ecde57c5c5bcf258fad79a182;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5994e64944ddf3b46238abee2145c057b9490895ce90c740f226b25415d8972c4afa3595f54dfdac42118b665ac1d1caae33c7f6eb87f15e5f3082c81a27990803f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2eda107d614ca29c5316ec347550281ee55f75d9723b2281d7f3fb6430451013d21f8079d84614f3f30eff3a57dc0a644c7f8653a64d5773a9b0eed9a94cb97ad5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9a708b65850f14792f34d2fdb5ee14316c971892857b6f1708e62cf845cae8e1a0c882b76a2da36eb7a7786c41c3b3584efb609e094a98a90a9b28af4487c28066a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d4858446d751dd3648d81c0b697dfcfe2c9251fb7c0baa15c310b6d75af7b328d897be3b729d99adebc2ee40af1a64dec2835e4803fcc0beadb15b514c799c50eaf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0375d1b4cb6c90f36c4a4fe7bed585b0f2708f75651d52268e237c65defa515463ba210ceec4025e519f0be40a9e3ca0fe5ab8d962c717082e4a056619bb6d6811b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cab5c226b274c078c97a6c82f4b61c6e4456aaa8673de9ec5656a9a5fd899abe8f2886c3c52552f03b0c1ba792c46c3b77acb93771b0ac4bc09c8a7d05120162485c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10993265d2d9fde045d19c9b9bcc47795edf35000b6858b83f067b62da877afc99d31beb5f01c1f7b255bbbf40fd1500bb6c7e8174d26e0b089c9f4d94f6aaa7ca8de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5f73eb67b78d935ee03f790ef702733562bc01d83eb00c6fc88eec4e5617fc1e62a32f9b7d877c3a1df88fb0b54e0057c1e6d28ec824108a86a69e07e650453ae21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h252f7c23dbc8e7329eedfe58c93847b9c3a44386d792aaa306f342607fed785a0c21cee0adc5edd3ee075b4b9f5db533d2aed119d3862fa861e2d3580ce1121f2360;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a9e2079ceb1bdf9cbf253a9f2fa6cb9b7a9b4b401c920f8c9e1d6d6de927b6d1b718df14c1421d8027cb16992bf5c7f5feb23c6796df7cd98245f4c1eeae81449e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16753becab621f46df53d4069157c42baed3a0b1a84312e3da096868a549269adde5fa143de52f2fbfbe979d28d400e2c95434aaa01dc6487e79154d39f598b1c4f8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ab9ac2c8e614bdbbfe9f7e4949a39ffc33d16f3b4526dabe0569617580bbd27c989ddc63d25b80973f4f5ed70184928402775182ea0af7ee774de2873c174263963;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a8dc329c154ab84e276cdc008dd4e3b6ba1a5d48e7cb3956cab84f27e6987eb43ce903c6507184f5fc50b7581497dd2aada10c89345b5b7f91e38721456bb8c960;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f585a4a60e54a2a1d4700478d5973c788fc70842d1fc5a33cbf0a8e0a77fdf26d8bbe05fbf51885f288ae57a4d4a29e7abd1b7b446a7cb9d1e5425805e61bce2a591;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8179654bff200e889384cfff292fb712b04481ca571dd7e00cb4f28ec90f30438134b0e3bbdae01f3e1657ce726034ab5949d1a4903533e9bfb2d39f484a221b90e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177b8864537d1b073ad07780d22c7147a3d2e26d5d09203e6711571d0c4f3459d08ce33c320bb15846e9811f60627475a5ebf73f42be5ddeb990f2d7366aa30471984;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131217190068894c075a07397681646250a74955dbe9557c9968f2391023fbee68c03778fd9c0a7fb051ffaee6dd5060569d3938f12a6eb5bd05bddd87605ef41f5d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6818329ca3fb80424a85802860b2ee36bcfd613d30dfa015b223a6cda2092319a93d79b7f4b0a92c69121fbb1bceecf3731f98098ea99cec32d7a11165aafe97da0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193baf53fa5faa25291054a705dad4784e92c4d9655263c9e7116f90cb515c99f54c13afe715dc44ed81c59fa2e09be01b1699c27106e74c3c26aee9cddff1bba3ea6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11da0f3785988adcbbbf0a75ebb6faf8e22e01a6cca0157e32609cf38569629e76d7ddfcd95e2f8ed8480e941d207db1c7bd286e5829332beaa714a1f5f6cb29535b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f593305fad2b9bfd63ed653df3708623d99d47035ae43fb972687843c2c25b231d6d2c04764504543feccfb1e2f8dd480b1b2a22283ad572eb95a1a08340e4c141a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fe6cb669594c7b96251b6ff15da83ebe144814abbb8fbc146dfab869ad32a43e19bab1b5cc414ac24de09b2441274c28741bc9de00c29cf3351220708f0a049bb13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfba67e0bd3657c3a1d057a0c8bc440fb9c63da0da5fc7bc9cbe56876005848f11e85e0c76c7413fbdb1eb48d84f6b9877e961ddd8a7e4ecff1b04f9596e7bf06a77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20e2ac9f3d013ff0c27e9d2aa507d807c13d479d2e5b37f33ae588aee87c61a627508176de8c7ce634a8992a65c6ee5bb2b163032e075bd934657c295dc0cafea00f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f82dd3a22256aaa9ca6efc69022fca47bbf5e992e847fc31aa6d97683d90a02d65b5ce7d31185c7935002fd28d6a9adb26ba1f28ede2d3f922959ceb0753c39e2b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1041e59df59d7a2c1d3d86fffeca8cbbe2737ee7cfa4f48fbe9bb126143390ab7ac77dbf0fffc0a0a809c3bd7846e730fbea2ef68b903971ae8fe013eb85df2e7912b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a703473e5e9578339ace8f94d2814742dc2f345359fac73e17a04a215d97a4ff61bec91882d93f15a15ee164d788819ac0f6ca0b231e77a789761204dae2915246c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c399d82af66aa6aed98454c704fc19f76d027769da12a20efe2291cb3b37b24e48906aebd1c6b5ff215c3161474271030d88356afd607c0f6be0e75f52463b9384f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1501d4e467dd4beed17b9df7460e3270007c30a1dad7eac931049de2fc885e5112c227119b31ee8704c5d1f90a6d698d0611fbcaeb58eef39e9fe630936c8c7ecaf94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e0c1fa9158b8b02b68a9ed089103274b494c18e56e3f4e0522b495569b5e8ed58682db33578c01e99c1b978c696373cce9891528248aa16601ead88685ddfd3d1ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed2ebe113be5322d94447cd955693902eca0c4d68494539eddb2a236908824e9547c6762d15082ce41b586238ebebc3e85bbf91976c2ed58cc3020213a60cb772a7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd49924c19dbc47d3471caf09f2e88f7a441291dd73e261111d71591e9eab349fa61936294ca0c4ea2a892fbe6ff74981b07c1e92149be09edc688426ae9ec48790f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c1304d7aae1491add1832c8cf20117966e15217bc84042e2570466ece1a85ea6ca1e74a03f73d69ffd2fa12ad6ebcbf3e667bb984f9e8e7d4e94f4dd3ee4ee5d01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72d713d0dc83ec3afcf2dd2c5be9de3c89bfeecc7a1fe35e50f97c732599dff784623a23e427e7a0ef3c2cec04f90f08347b45c1db1f65bc70afa12bf17fe578c61f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1435db4b05a52c8a526420483301b28edfeb8134014a6d6b1ce39c457f79274e2e08b89007217257dac524a2c7ba9fcd51ab290c453e28d3fbde7d1d6cae635b04ece;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efa29740270c2f1de0e4bcb30f3cc36406cc67d8e669065ffcae7decbe2636ab0124d715df0ef59af8f56a4b4e90e778ca26a4fbedf606f5ae5b2cce4f3e44530f97;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1600ff4bbcaa708bc1374b507291f47ab60dfa6944c6dfa656716266ed0d2b9cfb3488282e36861c9a0db51748d7c2bf0f781834e4caca2062da866982282792283;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c50d447a594fdb28d1b8debbe9f2816c2f07b209e92cc17950f3e66cb7f077a40d015de9753d956e09584882dde32a817632c26d902a581e564d0e398b2dc212b9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10061a0daba35ad3b723f227befa1d3aa316533386ea5e24174382b948be69acf77ff163e6071f3c8d1bbdb41985bd228bdfb4c29eb149869f9ff1132f94fc5f41e75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c42a8c9310be6313280a10fdb7a5feba78756265b6db89e9f2f00f98e0cc4f408ad5f3fe06b21fb0fa32e0c2515c6eb8bf5a88e20540d983946300cf96581158ee21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f09efb5edd12ba3727d7bd35e43cb8dbb0df7dedc4c4e81b154308d170337d13d0ca107aaaeabbece3a3336ba242db8b4bf09f66b35c0d5f1653989e634d1c592b64;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad38a13279107303b5db3241d1ba44cfc41bb586fec8591e5e412face39ad713f0f169d66d3213500e6868db6e15546db8e8a7a526e86dcc5867b1edef140145a2bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160f04263872478996e357c5d1a2be1bb56177df10f6da7bdff620c84ca9b64f2b544ea20d822b55ee57f543ea330ad7aa093d0583645d8b1061a8f02bbce4e82a4e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a045098979470f1d88c928dac0fc7fefb81e6fe8fa4d0d87cc7a42d469b97635277b018a4c000b94b4c762566debba266b6ca9ab1190310ef75d9cefe5596eeecfa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6a50d762039becbf14150eef61f75e3f03f5eb8debaa8f424b5d53223979d01c58bbc9f1ce41a1935ab6ecec239219c4510b460643af37fad3d2c78e49ff03b012b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h396b2fda3ebbebb4465d4989d74c00b329f114a5a05187bce372337a90f9560890c26bde4cefb963a85d4011b1c55786060365210f8f34516f9fddfcbf981d9e6662;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he58942dca80e1978421159d49e1c535ac9a7c77cff578b21ed3e1133e6a01c45082b3c5acec56ae92d8b852213d085eb4d20c9c82c531d98ee079b11a2c0e1f99a60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1e90851084982bc6a63fe386600aafc66d392330f875fca985198dd2641f5e2daf81123a08abfbf3e72f194bf6752c34b640b47dc04155f2d74c8dbd009edab5e44;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1775706ba0ac0a2c2e91644b9abb3c00481e4e70ed635acac5c56d0919695cb5f09b06d96d14e1ce3622c95b53392a36f8a2259f7d7fc61205d6217707b969c46584;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h555657cf9bc8069d862559d9bca61560e2a3b57e0fc0e30d8a5cac90036c0a21f28500d4275edbe5e98b5d570f4a39895be4be93eeb85a441f69dc1b4d0171d300ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105a1fd67b83fcfc2c0464e47fa89b4af0efcb491ff0ce7b626575cfb67b9025a9f6f0474b26bc776a3fbd135b48f6bc28e776f2ac5b0f2054dc3d5b1b9d48ad9a246;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he309578aac7ffd6a2f53f62b03089cfbd0a1b8526079c32ec4a6fca755896c7a7d68698b677d8e0252f7a05bd23264268a6c9e9520bc010d7bd3c13067e2c95c78c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75ee16f7fd04fe2547b4b220d29f511080c6751f234ed3490d37cebc43d117ef559eae270dd08e97f62bccb9b6493f4a73d85a3aacbce439ed7c297f078f6e091abe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f06435410b6cf66360784426529f8f8a49f677b302f6bd84adafc15a039dca5c40360e0529bf25d6e30fbc76b8b66ebf0d0319320df1bb9e3af8175a8151f14e66af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbf8dafd5e649b0f247ca0a99e438b0330650a1e13a25656c77f0c921103d08767cf7675336d5e7547a0950885a7f0895bbccfd14ef2bb97457288aea6e5febca762;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a3c487bdc6e733e90c428e0df3b45034c434b01d8694daae4c76439ca76afeef86515773adc74c32d4fb8c3c6843337f1838ddc2b594918742268dbb4818771257c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c92e2d4ffb8441b45f93029f7c5548d7e10493eae7211ba35d90fa9477b86c78f4938c1cd73bfce7d3737f53c23d00e96d88b4486c51840e05c9518018386be3ffc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b53356a3d2440faf2dead471742117f3a22b47f4c6aca664dc3f0a7543d423a7afbad414d897d66a5fb1b88ce575558bbd749b06c0c6a611d795f63834d0b8ff72a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1349e26aa3ae5a3c2204b12433398d7b3a7cc402719a7b2ca72ebbf8d54191ea7fdab61383f90ede7ccf2fcd747d5f7e110af1c3183ab09a24084282234403f0e93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha793c14c6cb915999604e5df2b82aeb6339be80e3269caff11f7ae873ef8fc6ab6164f528a2f4700e8af4e8ed3099e440ac88e3537b0a560bde7e96c82b71dd84eb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3f695f150219ea151ee85846be8c1726732d4f09ff04bd30bcb74366b1ea8e18e6a6e0039124b0e3fe2e72085be963c2dfc3fdd3fb21793a160823afe6f821fe399;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1388d34a40ba8a4f74f3a90689f712580c19310a1afecbc433bd2921e4ce9d0b244c4d3583c81ed7f8a802dbe5b2f1df6a49fc025de85a513b25cff4c51bb49698dca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha44e10b2af91011076bc229b7780b1105aa0d7eaef6ad30d59c5a7bcb998eb8e541a0bac14fa7c92615f9a7470c2b387fb3643011dda6d7d5d49bf784d247385ee91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b327967e6e18d136728dcfda837fb2a6d89ad34076d3d6dd06338d6052fad4f5afe7959d8d4e8c5e296ce0a2551d72a948dab42b7d70e86b14a95c9bd31e3c778c2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1410de3ea774acb5d74830a26adf30e5410a086624b0694ca3b900ca1cdeff43eb9f810c0da37ce4dda8e4630a5e3887c9ab059cfdf06879038a5d6c94bcc3caaf269;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c669c16ba6cdc54bff448493b5c07feaa11d29675d31955598cebbe43ef1bd2d31a0747a65c6d5999e51bff0d294ba65801569ff41b8c49b198ccf350ded867a657;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1cdcd46f42c2dd4a918b28d8e4612d4da4a93a5a88eb4489ae49339623d13c867ee94ca862e265d59f61ad54fc011085e392f5eedfd4c7ec73b448ef2cfb2280a31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6811424736d3c4eda75e9d39f96dab91bb253bdca2a46e5433b48436a3cde9dabccb2aeacb30b894a9a351b8b4091e688e4039fd665d79f5e2a91e4f6e4b38276f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haee632a78c440d9525811ef6bca69b5ce8ee6eaede09c280511dfe850bd748f798601ca9ad32d070b359e2e688031f6fddd5482aa56074ceaa5797ba866853250c34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16525cca56951aef25c060344733b5ca6abecd5ee07c9f30915362b5ef58ff90c50e1af6ef2717b15c4f948b079d9087c91f03f0e15c79a3199b6f348e161fc4cc95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155abe2bedb075bf0b6937c7203e8ca621dbaeca373abb66958aa68d520b42af5530a68b139a6f0fe0b5038c156c13c517b87705f5a5472781118760b8de3d4728b74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he78c75e11da2d25f3bafca0cc26a9249887cc2a1157044943058a8d83ec8a9a76749ee827d2bc075d19da1914ef24fa0a353a554af27eff4ff015d2a2cbeecedfcb5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e3f8afe9b0067f5036ce7ed29a091d8d5843136d9894c1a5c0c2dfe447a4b9e29c4bb03c80122dffd8aed304259d4bdbcdfdf6f60d842b898bbd22fc0a3342eab15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91e19bded6b52a5a0ab1baa0061648dbdc8a16317c7d0a2b781612e8344c79eece075981aa05305282129225058267480b150dd1195e84ae4e9ecfbdeb306d04d298;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8e54123625467a66633bbb8fe07e1ace8376e4cb2e1a3f5b60b722eabbb39311804a96e7b5ae93c972f429188c7e41201c3a3863c6c48c0df27f324daf1058329ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf3dd51d51c82829402c0dc13b3b8eafaae6d90330d0206636d324da46658735f4b527dc6c64abc044a997927b40ea01fbb20c3ec19516a297c4860c8d66656c3e15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32c99bef5b7cabebbd5dc2b5766b6d88f5ab51e54e374c8e75c8d74774e5ae3674224e7f0f905db9874520aed2b35e7d0d66cce614dcbd53e2674dd72119642eff91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f389c77446f459f59b114bc392279b93e5b8d4b364a9285ecca985009a7190de2553496ef34dbb11208fb946f03b3767bdf18378f3b637a622ea1d453fa201896c67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108b7c9735fdd65a0b2a6cd361e3e255524799d9ed53206619ea8a1146cc0dd808d5974dbf439c472562decb4d1f06cf20f805d0f9230585e771c85c2f7dd0b18c98f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1ef4a8ad52a0cb587666854b85f612cb5d41631c9544c45476750b342a85b019b4ca9c87e06cb52826d6cd03cf0625b901383a3e4c4cee82734b561701fa455c10e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ef8d49449a77487a63ea1cd52be65d3f46f8d4ca8dfd860a59cde25bfda3c44ffe91953874719910e33ccd319c67362dd041f449ff4c2c0294d3107e555cb157e6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca28aca8034c3a7b7e1b679d58f8565d408a87be9b018442bc61088adbb4e40ac7860a689b3606071c8a97763c6e742148aa69fd2290d7a2133a00163a8252f70a5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2cadf05a9801420c506e5d634b19380a6b43ba4e80bbd6ed3a8c873e97fd1c153c44e4305e5367c822a89cd1ad9596e2c52003b82b7de41797b8d41d7a94d7da36e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12503bc2158d22ce603a98dfdd87438bc8ae8695add97a8d3a2fc74cf049c91832e902dd5c6ec46dbba5cf72e69e55f2dd8101ed875facd62ee16fc02f0ec0a1c13c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34eb2ad7eab3f19014f006221d604cd9fbabb06d7ee888a30281e154aa875501ea4854d6c1107cf061aa5db62bd306c5064d010c01395b1f3d5eaa7a49d130130be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f938911bc418ce5e82993695860f10f0efbd038fa82a8fb9356d1e9c67c8b98bad9eb4599651ee67a1bcbac5e54e67a0bd6cff6e45685febbc97be4e471d067f270;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc44a539d5bf4f7478fd2664462d452eddd5790a63404ee2487b53ce60dde8d1504258fcb6ed0a9a5b75e07bab70c9ea0373dbd6ee532afc133597d088131fbe332e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184284b0f9aaeef5942ea78a039b2500c22f1818a118079ecc8f4ca3daec85a9a303bc10e0c88db40f45e599756b4b94b2170e54b2c5d3f25b12c216f44230e82e7bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a90d002e5d8eed202131848743cbfe5d4b435881e306ae393d1ee6a2afe397db4b79f980f1ff6dc80877e890476b1f0d4778926b3c85eada4b8a73e4c45ae99d2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af3123da393a0fc659b0b782e66a2123eb943a98174a4439a2ea9580201dc9f165b72c431e7181026cb80ba89187935dbd170a817ee23611b9cfd7370d67636bb264;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10879e79be3ebca7f1ef9365b96b6cc0bd1292f0eeccdbdac6f35aa4d977cb96d6be7303c0970a7b1c6c50d9cc88d4a54dc39dc483c5da1fb3718b560f24bcd54bee8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b42eab7b7e59d33e3f8a37d6fd51faf7df397615214c5cd548d351d7c04740bb4773fcca26ff642a1f20793f175ff5843e534503b6d24112ca67cb6b998ff98a6358;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fdde76a9991f38c3bb0cef8da70f3a94b80282f10f4ca0bc7fa0996887e0849ae799cdfa6c510a03dd282aba27d2db8a8b6dbf07713f0d7a8f1dc7f7b6316b101d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e99366779ddf0c03d723dac1eaab5315225f183348e172e79e9917b98b84e5552b4aeddf75c64e8130a0dcabaa1cfea5038e3530a96bafd29663c2b80fc16822370;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c0a149e80d5099dec1c2315a712c257f9e43f3297fbd885eb564c522342848da445c16859edf0140c3b04f703ca9e7d3471b9c0c40ba65f1218f835bbed4d3e916f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1929e84525e1eeb1009607c0c4d77b23b8872090ac39cb6a3885cfa8d6ae5c93007b18897ef9250324e6555eb67b6a320ff985b0cb75536eedea2ee9548a63ec10c02;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha593f5672f3c3e6cdde72ff1ec3d617d9d6d90b7d4fa0b6cc9a9a71482664905142e6fcf39bdd6e51eb0784edd7e7f1b0d47fb4bb9c5384d9c1b315ae560431cd415;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1229ca1f77d9f2ef4831d016eba918c92ff783216333777361139bd4b44f10d71e4e1f60b25805590468f04809e1a83e29ffb206ee159848487627b0419ab3db1bbbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb352c874323d5181e3470f8128e28ee57bf4d6190715cbede338586c77544498fa5d610cd7213c9c3513896ba6e02af657bf2b37ce5e6542940c160b122723cd3ac7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fe612dbfda605679c1042319ce7a7d6fbf71f88c718d633f38a0cd7f6a630cd4ab3a7fe7bb7faa28c82ac6dbbed808068fb429d690c0bd51b728253be77b8759c35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bdeb77dccd27de31785cac02572162be560e10d1f72c3b61f8a113ca6d2525233ac320ba4be11a8410d117ab3767089dcdf3b38ed08fc8e2e6604436c209ff436bd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10565f0289925aa37c180c6416a2c543243f8da792b3490001b51e2c37cee5c1e7ccedee44724adf6a71092fa403686f0d8e1001dfe599d8ebea7500c5eee3fa76d6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5ac00004b3f10e64b6c521fdf988b7e0771ff3a34b5a61e2632a479b6122974b685712de9cedbfe3555c975b4a69a598f0d8e7c8aa1b64d35323c69e4367a03b4f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6b5547076c58714e023b7e2eba275f7eb2f7f65fdd38f0c178089ff0a2263dddd088b85a7b4dcc1f47b5f76c70f6540aac4aff2e4995e7faa1fb3db1f9cf6cfa1e5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1090453fc88c5d8400b7805116ca0c8cb34cded90860478d93cf019ce26d516b06e62b01613d7ec720d392de8e9e69eddb474c1910fd1a7c60b2f05f8a1d09256116a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b269c95319c6b2703fcf35a8d42e9dd12600396409dcabb44b4543da857c3f1c13b63b3dd88e32c809167c86cc97784992b9d82d01f5632ebacc896f02a953afce6d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6c97989ad642b9188dc486136a719460a89de2e9a7a0ff0db43b3d5b640f44cf272b0becd26a763c984380d694d69ff960434fe60686f58e8e5605d20911ebf19b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4201e2ef7f33fb6eceadcfc9ccd8b4977ae22c833bb1e0aebde5d3fed07fc648405d223a4194ebffbb8e7dc6622ec9e732285665ddc3358cc6e99b05e648ce723d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139ae8f355fd5e0571c8fb4f977edd488e29c26a0673fdd681409e3b15cad98657483221fc9a8161b997a151c723f7e1aea35b82db0023a9f442bb09f838e95526d8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c830a27875e21c3c929f90ae61ff185f14471ebf4b859e280f8fbe9c5f07967744fd0f809114f918d11dd103c958d0bf9df718042079dadd379e937e12b60d27b458;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97ca983bdf4b78e796a6c9679a221ad765ce97015aae9ff4459924b7414907fa5f0051f4726a2f33f0744f6e552902b98b3cc97245e0ae34bfd136b3fd54b598295b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a16c9320c67e2a3f6faa060147123b6e894360d7e6bbf7c7785035facf2bdb7fca9e312bc2304596535ba258ac5c44b905739841ae1971503dc199df5931e6088a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b15c76e3b41e5be0db7d468f323c9b2029f6bbb54fd1bd4b711aed6a7bea50e0937da6ebbd2e6649165a104ee787e2e9823bea38e8a68edaa0d2bb47772e6cea53ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fbbba1aed72f3f19cc15bb82f025cca3ebeb029996120797542bf0fa84fcab231dc1410531f6ae29b6e0bc7cce3bc348a0e8f1fd6f7d55d370d937277cd816fbdb6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14524b3415c6d4289fbe2cd1364e5b4a19641f69994411f6ca9edac2f703f100939d40e4c7546e87022105de1efd917b5f8237fa57c9f8df9e65481473fa2f9f99a94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117b0608e8e28daa756385fbf53a68511047cf3df8e7608475bda7bc4f6775a3129e854e62e333706cdb0ca4f304b1ea58fd5ccc64c18895b6d3e991e73579d9efba3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h658caa96beec6a2b471f5e2d94b4331b264311a81aec513919ea70d41dbb8e2b581d1f3ec1a6a557dd47dda6638a05755071b152dade17d1be3af1e6cc92024dfed6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e046f0c80a2d58a0ad21f0e5b53cd5aa781e46dc2f1ba3743d31b05271b35cd5953a9554ec61cefc9b4c068ad537c1f8217f1c99e12ccd691baf92a814e4e1eeddd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14aa11aa725998f90b534f5de1394d73ce33ff9cd19c5543381c6faf68de034b5709767089d1c59e804367843e499f81a312f7ed6cdd22c272e466c6fc40801edab10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10382784b7e39d632ca8e3a657dfbfe8804022b5119fbe2e71c9ac6e02025515fabc6d24c8921a60e44cd7f16b077c346210625242ba3e694a587e3d6c0e5b93870db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152f0a3d97cbe6d479896c0144f771fb24946b8ee3a6599f5cd6d367b5d8e5fd26de534d6b834f4acb3cbe3348b2bcaeb8b7e2862d6bb81805ff2fc6a4fb5648963a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36234cf6c9b3f711d145c6aefcd93a91dd9ef607f1b2a5f2b487efa9f4de69a2e5995dd119791f1cbf324c1bb4badd9888999d1cd9975be8d06eb9afd0566e06063e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe7974a2813ff90e86e090bf8d5979e3f8cf8624721f67747bfa74dfb2b98f1d8e43609badc86caff63d1c18d0f68a8a17f317aa7bf484061c2a8c9c1b180a157948;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8415a6d011af2e326d78d1cf14c9ce51a79f3791ab64aa2119f20ed13153de599e57cea59bcdf4c690dd98e3f4fdffdf5b1dfc3989335ad9e1952f8f3c7cc6af819;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc95444e0c52422b4f9d1128bda904937c404afc03b44cbc40bd8fea08d3d59277ed59af89d7d0bfeb9252a58dbb6125446ed5e61bc2708b9aeb094d905db926f277;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a09a9943ef5912a0506f8b262443082a389312019234a09a6d9a313fc7df32bc95f758eb18f250ea1e512eb298e84e6c7c24cbbe5a00ba736380e547265fd28851f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18139245e1cdaa4a22631950fd85f47f3164c281e40a3f920264940d272f4007873fcd24cd76021b40134afad07552102b8695480f52566049efa2ca9b5312cb5ff3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9913204b8785f6708b9d1a32e9dbcd5235645dcb3650e7c994a1dbfdc2328c66da742ff35b1a232be154b60ad893962ea43492974b7b12d503340ed0f7bdfb7ad49d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10798063fd31d6f6d9122b3ea1478952f543c3d5932aa7ff06de8955a7c7fad34f2e103a844882c169aa35ffd5fe4a6e6f5216467fbeec0fa74ab83549486bac59862;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8d13c70550cf5eff101928adcd985f321ba107433eab0b9de8e184842c83c2a0d09c0c16cc7f19498f2c36050ab42818ade3c2411f033a1b5e5d0644c28526ea5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c78b48f875629304471289d6d28853d8091e093e9daa74452146f13df1fbc57a3d493c0bf4b59d3547e8ca845f08099355773324ca0d9536da47c0b8ed3d0b52a535;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f587c0852111a858729a1410c5971aa33c12f0a5e6f18debf3fe61404070192295754d5d245158058c928eb38d116809460c6ba4ea0f1a5399199b015a8968db0fa5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h790c8c34e159efb698da884f3c4ed5a6c637d83a2ec9d97c7a6f7b6d86b59c3e476a3681bdaf3ac33ee3cea30bcd01b71358aa7fd6fdeacd666e5c9d322c18f9996e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35a7423c44ae0060f649f68d8591bc0ce5e927b2967ca1e2431472841c3a2802bb4c0fda4e560ee43aecf4b9dea7f67b31ab74eaa5cb16098ce6a00540f6a4cc0bab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3af41715cec526640a3ff7ea88cc174dfba76d34e5797a1760847f432c3980f0a27637ef7ed4dcde7744a20ec8b44302f9d93ad4cc166ffaafb2904b180046ac31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha059ac79705b79f128c410717537122c1f0a8302b9711c8da39ccdf722889fd91be486aca627d26660d8b3a9cf8b9de95537a0943c0fd61a5cdbd5077b3288e3f5dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e9f1da445bacbfdd2d361109cafb3709f4073209b94a88534c57e3b10f9f1f33e28db5f8e32f11b3b2803183b1361e4f27618d7bd7d50f5e202f98cf0eb3ea351bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165e37fe5f593e59c4bcd33698187c884c0410d9de410e5324db44209b799b58ecbba7fdd58150dfae2ce8172829499211b8f0b1b54c6f2ad273d3954e8deaf05b922;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1575a178cd3cd9bbfa08f577c669cb8a7dcafa58c41bec1c6c5a6293e57609f5ba3361498130c63b37160a4495c96e3f1e84151df857227795d45d293c49e73803ffb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e973f126f13ac159ddf46cde1339c0a763406aa27a9b97e5da9622f5c0ea3e00902ecaf2fac6cdf5b2f6d8ca31c9b281ed19d18928ae8172defe514aac9fbfe724dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae846d993078e64eb3dfd34b02f57bb5373a8f8e5542beee78d0869bbe05ee76885fbc00a40bd3459b37268f761fad1e04c96edf74ceb041e7f10700394256c4e01b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178850dbc1363224b944bbf3e0c18079e49bc6b97ddc3cc645070a1f79d1024dc8c36f359e26121b8c9184c854251894799e73097951fd41401b29f2ec47c0a204231;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125c97950586b0beff68725c879c85689394efc2d1aa260b9e4cd34bee59545e63b808df0a30d95b1769f8c0dec7756d23dc45863408966596634b7b40caf2043173e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h844762982bd191391d22bf9040be469b601b70ed031bac20364ac42e93d841b4394fc2d4c92c441f4d3aced4fec5377979568eacbfd5f2fa7f731402b565ff3040c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b34cc62adafd3042a39e3520dc185f7d271d36d2883ffcc7c2d4a4c27f849955bf989d0289341f982171522f4b0ae302e90e7789895420613acf27d894e043c18a54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e2bdca6295efc2d604980ad6fdba1d459637bf1057a4830161f2c3510999c362b3633105d219135f145471b1504d59c6959a1369c6e0a4ce40bb0ad940f76d4fa5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115392149c4fcc92214e1735cac86a9bea833e9add5459cdc7a07cedbb20c6ca4f6a231b60652cbed6270330503f0511bb27aee7613b5d108edc7f909e526429eee1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9b0db6c45a745048ac50750ea1c151ec28a0b05fc936ad9eaae315223cd5c0c31e7bceb2f280271dc2eac13fd5b9a50895943f329777b147f8bac3eacfaad7d2c06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcd6bbec6b5f92345ca9f5f8778791ef67c49c772b1ebf115c83f88a8b290e3d2b361052eb5eb3b74b68c36dff6fc92fdacda3ca7135e3ffdd185688d3437f88b191;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3994bf9873ae5951b7f64132b9f0cdc1f37b3e6bf3456996a8313940390faa8010cdbdf0cfdd7566fa7fda4b1098b5fd4c8edcb65f0fec1d8ac8a8f9eff17449a3fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18769b855898f8e191e0f346c3ef764e56d0c369261c72b200ce650278e574560611e4f1d4574c856089a03c7d341520d7fae3fe9d07a652fca42688adc8c53dbc15f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a4720ab2da77f6a17efe4a0160cbd27716ce468f55a1d5141b0b1ad7e858ce4d8dcce2fe608bdbc7f7214cc318f867891e133a2673bc615c177c495dc19103f2acf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d37da14653bcd62c2efa94dee2832d23fb4564d64ff036d982e2db768578e588a66b91293b02198b27d4797a6c7492bec402bfc7fdf1d759339d7d55bce6fb5485a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105b5c144251b42c42876fbecbe48ecc1033bafcb2697ff632b6841af208bf3649806989ab24b25ced671a9f4ba13308bd8f932667456a44b8ba4db52200b8ee21b08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a63df8e5b15b3f23b462167ec5080501f609c6fe565d6cec2083db69ddc7bd2444b899e97f92395fba83ee1004904c06506733d53f2eb7949ee131ac9bb1ac2d3ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149f145f0171c2958e4fe0cb30523a8463946b6016888beb20d801f13c9ff8795025539d4d79498b0f8e454b4491e0d3e75a317cf93307068015652b5a24ca20a5088;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182be601cd3df6a3aab4b3144db32709886f33667fe9435d710c9889934408219b7e57311a63a313773f9b04c25d430922c46d9288c15335adbaec441b1e953e5b4d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f808b719b86e1a48b0b4b3460584170bf3dbd1efaa1525b952afca2524c4499f4cf9b8d51ffc1639ad3bb42b7620e531545dc241d75e5135adceb955c1fa9115d7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9fbc4ccce7f445a34043e724eb46c141d9183e3df5412f692d3c705e17737c7cf6260a4046ec0844022062ebb8fa747a0838ec84b60ceb08548017ad24c069e7a0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16202e752c271a693c60882db8809b9f5ec306264dfbdd3d107de06f27ef274d78fed6314c5c65506f2153e319fe0b2c09c3fd8e076f4e93f04ddb457836f70b5f19b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a879cfa47d49b5b1042494d84534b531bf3ce8b7c2e1d8217507d9e0ff85f0438e594853b2af441adc283c1a370dd0e691b766a26819aad259b71cd3f408669db4b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f860a8339b5fdc5ed9cccf643bd61e76c80cc9a8bc49a97e7216c73daf777e05e1c37419974f08c4d2da8ee5ab5805c9ac74e46789110b84410cee7d7b79ebd6fb8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bf3536daafd6a3ffcd35ebccafbd2061e480137eedea5f257ab44133cebbe3128e2ba3a041143f60f27d815d646d6279ab1d4d279a0fa2683a4654c8d731239b727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b0227180c5e98e17fec56fc972b5553cbc87958d8d7d75b39b066e982427ceab4130bd6088bc640cdae334138f655edb218245b06de1a9cf058e3dc56c3ff558904;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56c77dac84d9e76d7baac6a711f9ed8191b036619e5d6c7aae73e09df6056450de53283e07dd554c2572da61258bc8425dcdbceb5179c327e775563c28e464579516;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd89242d07a35b7ec85857a4f165f9ac2f93542809dae8b978ed6a4440b8b663b114af0a222845b6c286e7fc3edb97a26f3203815b4840f9487630c1d2e307b47e8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1138486b8eac205123a0d74a9f1a8f4b73821ebcb61c12d8b8e34bc1813f8cb9e7c8e696dedbf67e9691f0303a8d03323be2473a29d861662b3dda398c73281f4a978;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7708ccff3028f417aafc26e8194ae8191052944844c694d27f5717ef465aa1c2ec3d09da09c1b8b6c393150a9b4ca8a4da98efd3f4ca0b9d07763100cc4c5bbb331;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85bbce571da837307d60903652aec2697ecd46fff3a207c954dd72d92ed215a7f7ee342e91a333a2b314df257dd77b8a5b8e034d8778101408aa44a004a35cc32fa7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb3388b75a23d040a78659a8a9bdf5d806ce9e576bba3325d5e1f271f622e20a8098ee0b3bacdac2c51be211ea6f3415478d4962ad349c0afae34697988f2cd3e13c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0371b6aced238862342d2687e3fb49a87459f536ab07d86f7b36b75a265a39adc3aa01c53c900495f7d23fea27d573341ea0fa478c16e23bd0b0050d00d65cc7d92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f5548bac402050785f60a52d5a154cb7e292787be9eaa5fe38953df1af53163b7bee7bd4feb5751f55d108f236d93d7cc270a273fa0cbaf1bf2870cd0f6212d507c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93a639a2bfd3b19052a5ed05421ea07a8a8677afe6fea8e66d267fc8d99ea15d90c8a9429be772ef49f353d352afda207be41c9d6e9d9d25ce1c848a574675d14ec7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f42b2be55ccb0c64d99d50cf5b67ee67ad8c41f201f12546e12bb601e89ce0bc9ad176c22d3df55f3c405078ac8ebf1b5901b0086177303a4adc36e4b21e3d62554e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140d8aaea41a75c91230b546c02560fcc5ead21542dd4009a25e4c990f80994200838dd72cdc9c33f7e13b8e2dd9e2f442d22893fcd86404695f6fb9538b101eacfb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bea3352e2e4de6d20bbe347e18c66e902fbec426427d696270908af9ca23edd7ac5ca56500ee722df0119eda352e47994c7ba7fe27dcc1b59d7cd953fa91aeaca6b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf67221b3fc4bbe3adcf77ee0df2424575e546f5871ea31b941d86bd7288c0fea3b0e7da70b947591906b5bdd23a87ca4c22fac693fc739f1adbda3e88b4db3329bf6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172c315670bc041035737de0d42b0a744112d29f6f1f22c56d4870651d521a9bf34cb803d02fa583404c3549a07d5f9888d84895f7751e2ef907824b47f457e5f38ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c62ae9569e970075e22a10c3e6107eab2c978b9557361d07199280b2fa1392edc14deae92894756051ecb216ab0b24bc1cbadaa42d3aea5ac9a74f89e9a10b102052;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a39414a09262a6fe207a4c8cbd40a5662fc27ca63358e3ddf1249c69e49cdb007ce4e7adfbdbf6e54e3af47c3fdfc2ead46af336fd5b34447edcc93e3d50211cbc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h894a4ef872a098391c2ef5dc549faccacd380cf1970293d1922a2dd0b10e649c8067c51f02d6e19f9fc2d6434c73aafc87a57cf91f8affdb2cf79b66fc2fc50c2abc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6eaca5c362f32f1ab0cafeeefcff48e8fb721a3e836692eb17d981b2d47686dcd2a2087fe1c1dd579cce97d2caffa1f2442a942f1f2484be4ea3f5df9a702d7d2e00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a898aabc4ebfe0263733f5595a92cb4338e0a186ab90c3b7fb7243358950fc106ef8a235c8f79ad289b30b85304a9c09eb88945d3b63d22d267e6ca87cbb69362bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b42da1556607bae9062a1fc6167e2792f578a3b2cd689710c75d62c7b7d4cefbdaa92d60c3272c3ff9e7e5b269edb52501caf642027a400276115b4ee8b2de52b8ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143fd85ea3bf5a564782aad3d0f18da545d9d394c464ca5bf370d704ee533ee39b13ceae1f0abcfa9aff011a7aa8bab9fbfa7e33ade9fcd2520bdf61d84bbe389463b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a3d592a963ad855354cb233c0b4e16d1dc5beacbc3762613ca8e519c431cc75329f042b3c3eb33d73edecdd634bb380860fcfdae47df950d05e898583b52ac06fcf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29d28f4768968958df5be730f02abd1ab1440b8365e61a5450f244b6a66d841dfa4d4cc08ad1758deb1b50f9e4e2493740aff49816dd34dad399f7b1aab7c098f200;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9b412ee0dc75daa257e917a0b8441583232759c004fc498f81c2c4484ffb2a60713863b69a2bc19565926ca4d2966aeb4e7c1ea80a6ba7645e3ee437ff55cbb06dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cb084741e311d5f84ca3ab5397a9c5cc72e6d9334cece1706957be376f71fd40b748714497ec7ded59ce8f11497537d7c76b987db6b61b4774fbc9ac6d889e4ace2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9ac52980d4f64cb20af2eceeba3a49bc2cfcf0ab5589ede42b4ecfa02f6aaf44935c85f1643f880b9d940bc445bd8bb7982bc77ca295cc6f27134bf2d9c38c78ccb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b55a139d2c0289b6f15637707b7bc4aa003bec8c87c017e4757fd69d1c048099d4383986eb8549a1c636466064a9f2f51d4a9c0a38375d03e48f5dafbd06dc01a000;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8781070589172c704dc4ba6f489e21b29e51122cdec6391f9efc8989249da86c949c0aba1384f5a813be28da5ba7af77a0fa9c407617e7c71bfef3e807286c67462;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfeae149b25d989cd0acb0d549838e14ef316117d6b7d4901de8865f6035b798fc6e7459a45a068b418580adfa1475cc3d59df9b92effb912ecff56cd0873b93cef00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e4a59d245ab8b11702b165c4e6e1f7db9f7e3aca6598bec7e981db4adaf19dee3900da7de8332c16b5e7ea8b340465d10142cbed95cce8894a212d7c7d4ec3fac38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10163cf1ace3aa5fbd345ca782fc77121c7af9630f1913d2af3cf28cfc9a5983d326c0a406a2bf3612ceb958fd09f77544115ed2ec54776dce06f1eafacf1163c627d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58dde11985b961d626fd31032e523bff62624cb43de684fee88334af957ab2261dabce442439b53093778d7b7ef6fe278b8070b7b0aad2554b8d3f312f23270b81eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1953116f79c845dbcb7bf33cdbf64502b00e0aedacf7d217dae08eb53565f3f7e617cf03c2321a5af5917f85da25308fc5dae6391ac6c7e127fe7236fd5c618783c55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd45efcccda8bf47eef900d16d65f9803161677201f80921861139aa2c91bb48c3483835723c37f9f5f8d25fb4dd67da7ea49cdae97852f8c25e98e8fe4be3b15374;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62a638c7eb793e75763a5426dd3b846f8b149bc26b98000659bed798348e05e708e0eee679ba200c740afe16686c534ac14358d6c5e2e4448bf9ed1aa61fe69fed19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2efe108e3f487db7d9c58b7c09434d3b875b0b8c7d6dcb50a989846bf3f51a47fd434bf560718932510d844ec01ff984edda94be9508ca47c85029614a27e0119d85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h298a582f593d25e13a3c2de7fd5515e3b60cd6cd84dd10d427ade31bf5f77a656ee8f9f7074bbad8d64bb952d706c52d94cbfb3732648c048d61095a96e9f851861b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104bd5d70144a7ff769a9dcbb0c6a6d74bd769e0c2c563c35a1d8f2a72cab9d3569cca655f309c601955d21f06c8a5964d8ea54b0a399333841afa0a1e9e111774ee0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76e61e0f911f8b34bf96574fe84383dd0ec36c49b5c5edf15db4b797d31c24186ea7f76e02f61c065d47bb2dabcb40f2ee60ad7f0ee150b6b364f6c5a2fa13512a3c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cea5f1dad1184a629146e6660424567607f47067e12cd7aa99d6c2f5a77ccd0b66bed25b8a9e4a026b3d34e844f03cce79d809e47126c9e953f0118379d99bf458bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d25f48c0c9a9d762b6c64e56c63ca0aa0428e63f8e1b8c3b607fad5d6b61a0b1b47a678cc8004faaa6249361b74adf46167794b63f48d19af75e5be4c853f48c0d08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fdd1173cf3e424d0f5b6970c1b5e091136ef7530ff6de3a0dceeb96d297a10c7015330fa4d6d073660c895f897ac6585d192d8997315010666511bb7e6c622b4325b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105b6fe7a1058773ea0e347b4d496d339071ab5bdc659fdd25a116ef9e549d18ebf8389e92e6ebae7b10290859e54786fa311f8a47c7a03938df4ec8532f3b22106f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8f3205010e0a29dbb424a67e31916ce5e9916da1f19503780370d29d1b7765465f2f5c9bd58436f5eadf2e8c15af2dfd9724b88efec9d79a4c135cf05cbb061b51d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd52870ef72c07c7c5ec87feac72ef1b0465243fab27fb3b831c1224ee10aee1fdd4cbbbdd8b4ea234272c261a2d60e5b907b2159a40e5a507fec36ad91ff45efb90a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b67c2fed081c337c167d0cb3cdf33b636abc29e50ed65c6631d184067b3e5cb9e889a56d73cffc5bdb4507847c2bda01d36332128aa280bc0db379506795ec8b0e59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bbb62e59ebb91864519c5915cdb0ee7de58ae7886d321bf1f411274a2d41a45e5025520f99663501f7b42a418abfc8822554db1998580b587c51ed6e6a21381aa32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f56704b1d79545e0a58e71e9fe2a2e501eaf8b04a6352b1c6ae8bcc4740e32765ea383cf8284e40ab1bb5b26d87919bcdfd120aecfc16ccb5a6f2702b8c0c678afa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77cd6734e77aeb210d24537d5dde3617122e9714089351ead5593e806bac86ef91d9d8d111deee83e8eec9dcb49049615d881081d4217cdba14e819eb323153bf4ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c77a8b31248f556a8a22a51f5692c3d6771243d5a113678e5ac6af6055061bb1145425b4f8c3e4d048c6b893c63b95e44a5fed406ae8fc4f51553d382292c630d489;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e751acf9e0517dbc7d8c8ee026efacadbb9741532f500e1fcf5a26ee09019237498ca51cfe50fed4f640b86ac9200485ff46627b4113544bc5b44cae6800a5137cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h628aa1a8057e9d12cdb712838aa72a38ad59191791c26e75279ce9d81fd2fd34bf85a10a72bc0aedf04b76b18e6b1a57248d87065971bb6f408b5b4627d7cbe410e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6a00a3ce1e328167c12e84294b778c8c5c9ecc24c579dca6fcd440f3976abe84e850e6d038e718b0dfb2a72487cbf2cf23784bfc608d3c5c2c5e5ff73f8685e1d85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98b4db61c9e7f44b0bfbaad37461fabeca5cc373ea5e57c37399db5e1d33d1ce3b2a546571cee2ea92a5bfc15619120fd91164102355cc08bd07b403a0f38593f1b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14988e4970a681b68e4bd6c8b7bc29e14e634596e1a6088d470f9777dac492ceac106e315261d25280ca01d0f7a96f5b8e8dc31caa15a3d9c77b5d8ee55e3ff22388c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h612e5385dfe9c2e0a153a8145f74488c7db5afa2b5e655e4c109d898be3dfb4a1d28b8c338904b7ed4d3924b5b81cd1a2c57d98e1862ac95accd4abdc13e76b94e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1342d8c92ef92315b6d8566add68ac233a6e3e4816c0fc3cb4326f7c8636277f04273e5100c0fd782b0006968f6e42dbf3051e264226d09b078f2a910d80fa240de96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac6257b8a11f07d938ddab646339cb1d203a06da57c9e191fec8c9175cafa6295a2759e51cfa04fbb5c843fa4eb60a1d1d82b0bb73108535093716f402b604da6d8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113f2efea133443dc76feaaea6bfc83f8e7985cc8de192d30dc498f4d4488a82ed9d31718aa23272fff20e3f2725283aeb67eeb7a769ed5fef6b216b6c4862bfd6612;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf95d42a8b28fe569b4d5782d15d7f16a1ae9be8bfbec296feead444d2dc9f5b5f704f183d239e69b77284bb8d7126989aeb28072e1e716037157e67968d4ae42bd9a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c7cd4ff2d0bf23ee9f6652daaa35ddc99de4c0b593a27a89637fddcb41f741edfa988a93964bb30cce4a7878b97a79db908c1b0adab257ea8808871ad8ee847c9fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0d6c31cf7ba0bca2280b27b630046ee69440c93067af9f1fc2297933be6973f9fc279c7b69d1a143862381348540709b50f1260d0ca3e866c84af4d5c2a39c657ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a156c8cb217879db128297b72325185be0dfdcc4e1a49d10eb2231f756f56da9b41ba696c6d8d01cee5a34806bc5e1a64e8f1ad35cfba38d0143a7ca78e06a8cd382;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ae3ba686571f817bd476fc07346b689ee176e2396544bdd0a109f543a59f4e6453898a2bd29e2dddd8ce269afb65dbc989877317950a4e44b8f4b514ef7a709de51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6bae38be761bad9e2ef2cac7762f7c12ab26dd2f337c43ba7f97bef0708f0fd226be2392fa4e1afcaeb83e8161489b10cd5fc73208737a12ee8e4000ea260e4f3a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106b616aada1e4db63ac451cb465da297e17e33d35b5e14a2a2967c545404a58ff99e3aa2fe45e5ac5d72ae6b316078684229b3337bef3b04d4150a6ac558fcfb1282;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fa4a98b9b0d5b366872daa20f4461998aae365419bd9d7483e5d5ab0e34ab5043bde1d9715020b310bc572aaf4ee8587b5df7219ba7c985a4b510ace5efb0a0ecb5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c86986eec71209397f4121462a39dffd645c39465110803f3787f34c663af58dd4c12a0665fb16cac54902fd435de36826c8d42ef457627d588e910582829ead818;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f4806751e4d5a90b9559898ecfaa3e57f40be02e82a16cdeb182becf1b2f54152205a7b2ceb5fb44ab8cad4e020fc9ab1b4f9c28dc2245658361f2bd958193b9f00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafa5d426a6b383eb17c6870e50ab38ffb3cf89b4e9a90a315f928d5d4efa701b186d43256cefe686c4c75efa44744c35cd97b9e31af058950d7f5d3c6d30cdb5a5f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c43c773b6f9ecac4ee748da5ce28bba01a24374fee09be722efc5a5b6ef6f0755a455a364d775f5db105a1dfa6ef004b172c05e7de1036914626a7169b79b538567;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3440102c3a032ac286ea2d6e5ab299c4a24d36ec18f552d642f3f10e513dd0ca24a036ab3c055ff0a05d75fd1f97cdc4b7a662e7325906f3e00509119baa99a54aba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8be7b7677066b6fa6c88dcbcb57e19e369fccbc29bd398b2884c337adf28c3ab279a54039c8398b9df9ba6770b4d3ecb7237cd6393e6572142234ad63f51599aedf7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46382d669cfd5177d4e7bc59a80e3240518310ea5b3282dacff2b69aa78b7506f45cf81fd5d21041424cd00fe8fa2f58538f9461ecdc8d2c148a5f0f4b3d38e2002e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186b0df918c4e1906bffac7a5a199b68ffffdadebd9c48a09c588387a2b810657028771b4ed16e347cf43ffb86f6346480473037158611a18b805d9e71cb852d3a2f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbbff7c59106bac9a4b36f0989667ed0187d7f1d7b4a08c4429953a83d61be2cb628a1a066779e21915dbb23b7cc8b4fdf5ba72e3e5f0c586d46ce96f440d5b47e15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83a23fdfc25051cdaa9d7d076c53c9c08d287bd69f3eda408657cd1b5e302310cdd8cbf2ce0824f071d74790cfec5cdb8042ef79eef415bdc9e582a463f2afd488aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145d1bb000d8df066f46fc21ce4a338e0c298adc0658c72f1b1a6c71b845467b1c103e32d36092251d11b825e083ef71568c442438edf126a3a5feb29c992f403336f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11159b29da5c9fc63ce11cbee5aa00fd512ee06154365ddbcd2afa162ae19aadfe7fff9345a6069d3987810afd8ec3cc29c094f811c13c9a804776bfa1606b434d701;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fcfa03385051cb79d4289beb4584c30fa089a50e33f0a4d8862b3f37dd634424096cae44713eda3f3cf7a272d8be382cb56778043abf56c8c16ce5201a40c7fc5959;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfedac434e4912644edccc0d5a9acf4368985a955b04611d6e6742b21b3e83daa560c802d8ac38dacbe06c37ff7d2301c11ce9696798ab2e537f3ae86c46b64b9571;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17336eb7a19fd39c700603c22227c1017daf60cfcecbb015d55014e3fbb90c0566dbe56bc9a66968d2a66f8d55cb45a4cfecd52cf38a8e69e2d27b188b348cbcd7c61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119a31dc4fe27701e9ab8d90bd57851f92cfb4c75907786b46586bd6503e9b60e2bb5af97d474f193c0722d74255181073b5d04d46fe25b76ffe5df9c4baa781693c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b34ab0444926a9d560c030cbf0c78a0b2114bdf71ed81df792c863cce212394781ed15c7e10fd505bb0bf8396c24b5b465422b22cef1e7ef5505aece7f19bc48939;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29622df7ac4a9a81784e78568c9db4bf84faf7f59d7f616eb57000bee70921159047e84a924c0c4bbd3cf975adf1b21be4dd52dd48409846070ba028859cf98db39a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152bbc1aa7aa8f9014317f41d1b6b9bb8130b0cb14567b04f14cdc6224a455153c59fb210458a2777dffc0cff2fd0343f48c81e08369db222f91a637bdb2659b94fa2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cee73cabc15f5ae31cd83378fb1d06c48b239cfcf72c19c9961466bbaad0358a43646a47309d453031841a59325fa7fa453582f84e313b386cdc9761c268940341b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f00a963498a971fc228a92fa9e62954056f4a43bf9ce5ccc653512319e9189d8f9a41f6ff73b4f5467d98e9f7d620cdbf269ac474a37a74630321a10da3a28faa71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b4c3af2c0fee64f7dd4ae2655279b20d5472aa4d30714bb97d3628c86609d91cd8bee8b275bfe60c5ebf014bad7e0a2254d4252e113f3607e105349a8fbf1db2188;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d715248c14547c3ef3995dcc96c6128adfb6071e96eeb7893a8618ca5c62827ebd2824480367baf3a8014e57b924b52bc068c0dd0a28abf135033d539aaebd23211;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e80938e4127ac43cb2b2c30ca87b490267dcd46d71dbd95fa1001a539a749f46ca874c5092333b96e3558f9872193b2a7320bf28100a84c70a48da08ce6c2c20573;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc74d8f03020c24518d79f58982522f75a4debe58015ef004d1d824f6be76ae78797bec88b9b9b268e58c4d60d4279bef30022fb8f48f57caed1e877d3f19e40c4d00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16fba6c655f8823e976483ef1a407be5783114b27ecf7cae10857efa8b3a9bf0f9d6df2ae37d27912889d71b9d8511e77f05e5f135196877ce35399d81bddc665caeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ea227ef302b8837344cc2f2550ece4011c9b8d9917c01314bddf235e922f9741688e247b9f28b4b9fb11f351f21f15a0d30459d6b1ec7b7058bcc33b46ef8b12ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd2b8b1d612604931fffdede57f915ddd52e9f774f305d19ad1ec4d336093fb9d879ee32ab4488cb2760d65e1376721090a3c0bca8f5b2b01507ffd2c44e5bbaecad6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1313d5e91c1b0fd9e75d4e71ca292deef25cd16bf95c913d98c795e905307cabd0d80ee5b664d7e0ae5bf983e6f6974387ec61ff23e761ef9a8f798616e15a935a616;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h338c8dde68db7a06b00cad8d0163c4ef4bd5d5612f4c5a1052af2d3fe2600e8dbc6930383a9f6bb62959938d3e8e16a252cc831afc2a3dfba8066f8f00d38bba8210;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4491c7f9d812b121f962eacecec33d2b4bcffaaeac141588674d5cd5d2a488ecc5d0a157a95102f1e4eaaadc795482bb7614368f0e2989044495c04a7e048eefd971;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d4412a6ad427d71b280b1e7fd51c5a94b7dcbd0c8c0a56421cdee4e12ad26850b0c114a2b97ff02053b88d96ce6cdc4d2e5c3418b2303e3cbe0064df7c75d3d40d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde06725a08f69e95774b2e31e9f0a58996a689104bd771a5ba559f29c314698e2c84470549c424cea0ff684ac7f05a99d5c817298885592372e73576f60f85aad5df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6af089d697b0a5438e7ee84c53b74dbd4cb8371d733b17c58e0582e13deb3cafa91f7d93931881847c60a1df70795a2d90e1fdd552083694a48eb6ef158c47a20a84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6adb7adba9cb0b595cad328d20296f2a1475d524d842455ae809a4bcfc9b2b17f3767d1d1e9058d04b6478ff5f638a6a9d3a72d31a2e165d68bc6d1e69c7d03584d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa8cf280feb299651e534ac3f8a06ff4c56b18fdcfdf9af67a22041b44d2ec03b023b7de6fc4a6ed808affb308045360b47ba811c8cabc2d767fc70dca0657ebe2a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9c095002e2882d97a5db0e50eab81bc95b8d26735fd4170114e48257bee9290c366309da286af9143ac6c1da85caaccf2afa1eaeb3710c448e50e1ba416d6a4cd55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f797ed7eb25e04b7643b040e4f5ed22a5e31419fe2a4094e6b4a5212174c4580f5dc37476a5c82fd064b49121ce9cd4c139d0da3fb30367c122830f574696ef945a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e470e6a65db2355280a09e07463f8664c30a03c966e57a169e7055f15cd58d36f2c781f7afa072da803aec95d18c5ac7c0c7851c44e8d9cb4227bcccc15f426f39c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166a7e8a5d721b135564c3428de40bcc3156c8221b80f075f8471ec8c5940c94f5e2e62a410e73792024ae6a1dda771fd4b5203daadc03ec89ed09d708a2d1cf03d6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25a82d2e9d7971626965027f2fadc83de9d031349a426c0cf38c8af01e107eae61826be6183b9553024206a14cb63ff48d1b13de1877b8bdb442510bf0b6f1496976;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h943be95812f6a34c163c20af29c3709f00db015a134bd59276259a38fae88e4d52318864e99285f2192daab28c556724c38b48c3bf7f1b88aa458ab55404b9748dcf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19dc71a0f8d6ade32f617d272f226f2dcad06f670c20929123a7f7ef58d786752f023b2464152753176a8c872c9a8ce003aeb5765995affcfa8747f2067f106c2a242;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f376d0a0065a345db53938fc98e0eeb01080a5f515d11b27b166659ed680dd8cea0dc335ae9045e5bc10cc26139dc36b37e1b039f54605ab8ef03ff4dd1ef4f703f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6122fe496f2af60fa613dc2d94d368c65a77c7256a1225b6663d77480a894565613f9827c4297072854cf05b93dc2892c64085bd97ab2815886b27f3daea1e299177;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b3963e87beaf2e67c21af4f390158c96755323b6f6e2f5691770ae292d30f473d9161317bd171afc56beaffb5e99908df3503a9aa189b62dcb8aee5a6f274fbaea07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab65b938605071a03537fc20673f38853de66a36ef25b3663b1f5cba6c41edcc01fba1b0994353067a2e3be408198dec3918623c9583cc32f6c53ceba5697d35f813;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195458f542893e8a55c7822a2a56d730f472cdba55869b214cde329fb8fac96aa1362dd873f711d99f88e054e66f167bc73270bfe34df94f249f7cab78659bb9965a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac58669c392213981c220c9107ce1094a9fa0b09fc6d3638107a3e00bc0d854a5e0f6fcb26479c73a3ffb42d29eec5bd645c6c92551e3528de1764dc1a121d12cc29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc61a4db0a9994cdd05091abd88235a160643f6008b9a1c284869c690f45227828f311d8a285b92c0eb228a1554b1a2de600d1279c1649b1bffc9f431c5e5385bd1bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2971d4fd5136e2c7b36e21beaee8eec68bae22096ad36e9e41cfc01ca721a920858fa4ad68936f8abd7ff3854170267f9e6507fe4ab4ea084ca80e758bf9d8288b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119aceeaf393a838bd1bdbf686c760efea18c38f94e789ea6ede10cbca3c235268262cd2b0eb8b889d6cdd383158baceeb72a7aab2bd8050fe7de8ae65723c08f4e21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf999ce8c11fde3506e6e7586a1c0c9c2bab2633a93b4916db88a0ccd541264838a837b32c5cb33c4285b7697c0f4d05b90ad3ee7cd369d460c9fc3c8361654d59a1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbcf099d9beffdd14444074f1b4f269ea0549419da7906e5240860650cbd3f35752363ea0d06ee3133fbc30b3c1923767230dff8d03033bfdda99c66fbf8ffa96fbc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde6cceaab2f1354083acf9d399fbabc932c00e7b12f1c10ea9ff3bc95d15dfedbd6c4a713054cf0bfbfe5fda81364010d0975eade6321bf41e8f337d152d3b77d96a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15446b6bf052444540e519bc161df5234499b8dfd66ad1368651a52229fd062edc8969e06757b3defb313634188087e88127fa2fc54c4440ca439f7dd1a3715dd2775;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f9e6b4b290cb05b3b80ca9f9fef4c88423e5f5a3a7aedfcf20c2a8ac91a9529eeb5cd69c0a3e3b7ace3bb4d2920a5b6895e8b3cdf12d84b4a6efefaee7066767fc3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b386367268cea945056335d15916179e556f83db4857c549915045a62ae6972c0c787f33769abdf1eabe1d4580c01aaf08a086a30ac6024fbaeb2f02871f52db0b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5276224fec820b72b968a2d345960ead6513c1b919dcf38d396e886c6f1c04056dbbe73f74ef0fc0d370abff43bffb282ded89ea0401c1ea54a4de5cab8743af1101;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h436bcb3556b7c6a5a5c1fff2b16c9bc8e11bc65ac0d4506fceac4b7a3194042b7b31edcdaabf1402f5d0e50c670bbdc1a00a76ee9192bcdf20536590c0cb61410c7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fd530dfcc896594c9f4c66f03ce210fec5c2bfd1eecd91357e4898f4dae78c969297f2c90f190235d0a9a1ada97894ea0c39484918491538fa1f1c985516dc9934a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4237d85fb00f557db82e6e6517066755a39a91860b47ea5c911388cdbdaad30f99d981f95ae1b6670cab3105463303451979e63911b39228dc67d358960724f2b82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad838474638a93d1c30dee7e6683deedc4527e7138fda312ad2fd830cf81e03fb8ba6c8abd0433ea0e0e229e9d534b15d82ca6d4d790a9adca8203cc19334ef841fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he62f491b13d31fe1326750999e5d9afeefd49beaf6a860ac907b0126b569908e7c5202079e92448ba6add33ebc009775ecc28eb8318119bf687bfbed05cc504e9d33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c52c5477d17168cb73853d87e0bb06c0c9648c23707d67aa9cbbdb28873ba5e35ae0acfbe34e3e549d44364a6469352a7862c9d3e723d11d9923efc916c883eabc5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc595ba3ea7bcf596a65eb8fa073d0dd4419ad8d594ca2538d8d26763e92a5611f681e5488be16e1019b4d10bf23aded156b206923bf284ef5ed6eff2f8b8a84d2ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fb5b909c93ee95569c47d548ac2425bb9547de6a00748a117455cb3cab27ee6da4c8252f9b67951f1381a7e5713bb8c5097a57ac24a05a3646b987cdc02b1d39e57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2943d9d0ffebd16f7315448bc848e148cdf0d99f700c5ec7dbed48f324f382768dce67065e6df366c05364e6a161f8956cd54f8ad73bbfa73631990eb9eb442e2011;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1856c00cf6149759d590b576c821e490c11c25ed4b800500708bf6da6352f9a700801eba3bab5cd52e6c706bda2f1f24aa381d70fb55cb3e8ee25cb8c61ee608f3a61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d963ca9995bf62a1f56a01a463e765e628a2e35b121c2f279d6e0d6e78947051928d1f23d3188925d501aeaae85e9c3c39f3852e0e832a4a5f5e69556250e2cfa89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1178acc70e381cdd827fe829cb5abd33f70ef959f89a3e4cbe3becf974e98704be34e2e0379db3c4348a73834485c9e92d7406fbb305e9512f8e512c4c3de66e428f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1313047d711305d5ea14edb4849d7a2811ef185bbc6910587443aa2d72b984d4840249c42739b91d47b33c301b74d7d5b9b81691c146d200a9a15863b5e20fe9a8dff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76aed796b90cd2b44a7bc9d67df919c794c32922227909969c915c8df02da7d5dd97bf214951ee4c19efb93509f1c30b844b432def41fe799f705f89e248e3c921a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9b3074da94c6ef9b527bdea00cdbb0293bea7974f65d85028c60d5638b93ce2c55182c1e65688bd9ff0a2ad0d3eb96132c6898592ef2fe940a036f8d3b8aaa24e58;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162835f2cd24fe573247292fc8a5ade3c947456c83c7009408c43ffe1f201c53c59040bda9f3f86f8b1534776385dbe3b4faa2a764ba68094edcbcf27a10ca9ed81b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb25bee27ef642c550aae82b1f1c9faff606ff34d8964ccbcfee0d5915f18c933b14fb8652321413e9f415a4fc3e54e1f24b4218f026108bbb9a9c3047edcf99cfa8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f518158148948693520f192f014843169d7fc976780352d77e8e9f827b2b4787e785c002664d917bd032da88adaea7f975416d32460f80e7cf5867ef822bebff75fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b34b9d5b6cb1aacab7250b2da025a86ee2581240cfb147ab1995c96d7bd244ab29aca77b02716dde4e54644b1b7247deee28d2809bf88f8f32f81c3fa32ae798c10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16275fa0342b3b787629e59c5ae5a8640f3b2e64a49f2354c85e76fbe7a6ccaaca539fb8b51f94e7cdb2bb5d15473b221e07b95bc2bdbc6e8709d7268080e8b3a188a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c7af6d40d4c3569d6de231615b61337b969b4b35866db34263f3feb8880068ffd79d02623772ee3d217d573e6617f07773c937527e27b449ce37901839d104485e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dee13537ec358667b7897e744773ce2ad178cb7ec592785ddd2ba65f1b29ad5b3ab1b71cea975506f2f31f3ac43fe3e7e0a893afbc57b3ffa0ba00585c07b27ad951;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8f3b42a5cab078cc542511627ad488998e22016d25821be838b872f5c9a5c37305fc25a42fa9c5f4161d96c4001f7d856c9beea33e294cf2e48a817a313da8dface;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b12119079a9622387184f651f994ca9d0545719b3a375b7e096c5183a82f5ca2e543e0847d7bb623804a618ec3af808c9aa99aa3be8da76e7b440d8d2f8963e861b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69753e23c1cdf448dad6bee7304add254ddc3e146ee33b9661a355a61cfe80c2d20c5c32da2478afb054d1084d5e28c05bbc016e13705278d5833f02bad928c12580;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc901772c21ffa981450df7db6a40116b67a3b34194f8b8cd5bd372f7ef7cf7525a75eea0f074d0fd861400e87a9ebdafe978ab639c435341b200be7a37185033fbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c242749b23f88148d2c6471a8af57cdb117dbcfacf8ee1d72ac1bb07405a34052c24babd496e9c7d1bf10b5e49c4bf14d4fdab7923326f0c5e91c5d946d0905ec498;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a7c0c2336f44a2a39c7be4d9a66c46ad9ae2ecc9cac4680989a60c0c96125f0ee5766235bbf313dfbc9ebd10217480ba403d03a1298acc30fed7e5dc302dbb7b4e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59fc5bfa897d35e65f6405bdcf92e1246d724256e833df28ebeb0f0b2c79fa1958cf504861fa41de386207fb188b1aebddb35ad7edb38464578f5d9abad1de6241ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8fd9c67da7d1429cf6f93b6ee8b3fd5b9a5a112854c48f756e42672da5235da6811fb10da7b0a9ef2379ff049ff01ffdf93bb00b2559ed28d91c6b3c3a94ea09888;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53a3be5251d4e10c04079bbf6edc43b3b6870e072518a19f9c9ebf820eee6b7369c9c90541c9be7321e3eaada03ba8edb889ed3a55dbaef2ce723fdb2a9bc5a174bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60ddf670d4f6505cca9d17de84427f5463d46680f315776792a9a4d3da458cd403b461d3b84a67bd9a965a2e2370239f0d801d43c8315043d87a53f79673adc3d8f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17874f28ab2c428f0fd888440c37135dd3287c79acd298cff8701d31914a400b278f7ace20c54dbefe5a2ae6832f0685b72b853c013afcf84aaa7f4dbef52705dfd18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1691a16d0dc0e29597d8032282b49859b79ba339c81ca27b172a9cc380068be507d53072159b39f1e325245ffdb3f056a3b973e567755ec7f967bf633873bc5c11735;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfe06084c3d3f5476ee059cabb7f33e65e5f366570802fc3f3bdeda22f73e7f5556bacf390a6917682741b44b35f96574ca720b81038390cd9a29cf9bc420fd5cf9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efbc0702b55f3cd9b156c4d0bf02666e62693a7368ab10128ac294fc24463a0237ae5a012bab1c9bc9bd125f521101ccb6093e53cf89b7a6f286c7bff269d96ba6ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ffd09fb14e7530522301467aacf87486a005b67dcb3b28a32cb67a25eb875c9c94966769b9e0260b24c75d1ac9771e9b2af7bd40728a3072c5177aeceb00ed3f53b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebe390c50cabbcbeed57f6d48121425feceafc9b2f910374d594e0ec04f257bfa293cac18b08d0034a9b498f3af1fef778cce647a2496a79deacc0e4d801e789b5d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfddbfda0c71e96fdff0e2a21bde72f227da8ed63e45a3d9ef005ca337a60ebcfd9563927b10907f7f5e352ab315cce2a61612fd9885405ad5e78484b6d2420fabd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h292bcf071f7649477173676a2b804c19bb36dd1a661fdbf45ba2d4f94fccc27c1c5db23ffa9423c1f9178c3c4ffe06359d0614801ee988b6449086806d49620cbc91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c9a3e2d210226eb1ace193c7237e79ad83728de85dae05aa0818d935eaa955e904c2866318dacf02ab8eff90ab88f7823a4fe88d2fcbae2800ceff42b97c164f2f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had2418850a4ba1067687e7616d85df9194a26bb215c740c23fcbfbe0e521671f7d8f5b073a33017f437a4e7689e74582e6494d836fe5d4ee500045960c88bccd404e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2afd286a014a0f51bc8f110ce8a05520644227d741caf4aecac546e7a100925bd22b266d347d23c204daedfe8650bac9e98cf209dc928b5443baabfcc4bb164a4528;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca2f49aa8673a9147c34e409c91a4192c63d037bcd3f547bd76f2fc8b5454938c75af8a9e52ed1e880fbf6cbebcd760a491c137dab0851bff2e9f6f21a12a949cfef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he09d0688c5f9cdace5ee2d401e8d8cfaaa2c994b3cc373d72e761f037d922a69e79051463fdf32ee147f00341c8ff80080d65009ec3a18064637d7324de600f7a0ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb07a3ade097b178360203ad28c6c55755bd197401f1b8d3db5c1fc328e2a56172f72c0fb5d8efc2cf9b5ef0611c18c8ca4fec58db20cad2624a44c94cbe37904710f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a576c46eaf980dcfbf7704b6c27e8ae8ce574197348a112e35a990f1b2f6165dbddc20e6630a02f47c965fa4164385c01b8b0fbaf5ec4c697c5c2ca8f414a0c180f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfbda8a82bbbccab686fa87ff713c1561ba871e92858e1464983a617dd62508f0861fed8d32372529758210337cecd8cafe3bb4a676088b2c599fc883908f62f93707;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1767618172894e0a0cd3faa4f74d1057ce2c12fd4940d4aae1d80d5050040996cfd711063778fa1f40082d68bfc3f7506e9386a13d284210633ada3619737124b8d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c45115def381185657ea72c4626a7d4cba1e730431fd615d16e29c9c3ca816bc409d34edcec31a61dccc1dec36b47092c128d2f07b08de0e768c152a9488849c895;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac663116e4e3b6e505fd737e21260c674ed7ee15cb4f36e886300e0deac26b866a06bbf3b459c8ed9279ba28d7db267f85a9648eb4d6f30b8a5841a2aa351578b3eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdeaf4361fbe571cf57449e2559d5047fbf8b1c4e60307136ba88dbc9ea122068c0c77f938db9804adb6c2ddbc65bd752876cfdce950a26159c068da05c2f2d4f2706;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c8eeea87818c3649526fbcb73bb87c196762ca9fb159473c971c218f102a8c32b7c36821ead6fffb5cfee08eec27c2fc51e823be1fb635886310c74afb44b3bd893;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc54a43cf9caefed6ec40d3509a30c9371b9096cac353728fa585f3c22d0321cc77d0eb92ad71a85ca6b346eb7781ece8338078fbfae1ab11dec92b4812b8baed3ff7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba9528bd117fdbabf29242a030977cd12c954dc9592f9ece3b5df639ae08c88a20582542586d3edeb144a03bf86c9db822c80e1db1306af026d7e83f6c372550d982;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155be3877db009fea7765cd15d52c2ac653d118fb5abe93e29a95ffe176d9f600406f9563e1b9ce38f31a6551308585af0875c140b555f3b167a7a5ae34c1f9216c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h232220578d1b158e0a4cf520e58003116972d016dcfcd42c97899cfcef834e66cff4de71a983a04bfd17dd79bd83c85b1b6e27f8b794f2af69a3e8adb2eeab48cbbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd69fb0db3b808a6cd6da462aef90c2d4518bd548bbb3da41562608c4c1650d0955ce6309e0a470a571d308ff45d217f7516d00001af7ef783f8d6b0cd7c3c1e01ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heff576e05d41380a6fb20248c46c95086b48605f88317b23d2f00711fd18cce707e2fa0e90f2a10e00b92d57b39ff5a0d248d367064ba896176abd81c959d379f0b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbad0fb9a2ac391cb6f43aa8e67bde4bfae1bd7df273b26dfb04782eac8a64fbcc0700547616567b59e87fb78fbe6aa8a73972a543017935e598dde3fcbe25fd511d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126979b828a4f074a3cb124d44b9c2f832e566549b35c9bc04ecd01dac54f5724ec0c7c49bd69a31173201fac46f73c6716a7e2dd71221d340659c3ba955d741bcffa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb865a18e30ff1915be935af64a0e960c36fc14df7e959657cf82b329e826e70f38fa9544460dd075a8e36abfbc7a5dd942e72c79102ed21406c69dda1e87296fdf25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h932f1a39e3fc0c3c90883af936f6d972fbce819b19a6d04291aba062bee83beb7d6c59d45ae2cb26064b9796d06471e89ee975dd2454a787772f15c100a0bec3c7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133bbea46044ba68a64f883094759c64139b77e761942cfb95590a7de6ebe6f01902cc04dbdaffd1862e021681e652f5ee62d5d6e6af658db95e5270ffc8a3b7830dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd830212890336e073e58f20d6184e2623dba124182ea1e4d74998585477ec5b3aab56b0ce3c70b84801935e7a3e6337d16244e13e252f638e2211ad40275f49833c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ab4ee412a0745d1308e86561fba48c6cba8ef31530ef05b17a46d236f3615972961ec1483c90d35588c9fdaf0a4916e8ba346ddb1a63d7e59c61667b0bd21c44;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159cf15825154fdfd836af15f23cfdc91b45740fe8abfd146637869dd0708c67043d35a1b7346465dfad8a1242baf17782a992adf6d417b9b0538636533e3d00897ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74b8bf2596c64b96a2579a89aba6fba96e4b0da5ca516646f2156181114fdb759cedb8272c8dd59625ed410cb59d9f5d7860fc8af9fcb6dc05cf0fd522a0b7f70997;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a68e39316e0b774a259ef17ebd8c07ba56eb5c07f26ce6286b2a01c4b4a5e875e0aca8316a31e7dcef47f695c731416eddb1f6bba2a86d37a35ae60dcbbbae9ebef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3dda7833474e938c65ce5e44dd1bd08be8a2372bebd49053fbc847d28c63d64c58adbd019d816105afda6660990dccdcc11e8560c41b1aaf9cf18adbbd5f79ad245b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e4247b79cca2e1ab281def464d1cadf398bfb6c7fedc2fae011a70e07dfc117dbaa24c78335ba0a2c7e4d91828bf6126fdf75ef60a3379d9fd0b5edddb025989712;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1756666402afc8933e08abfa56cefd8f6b8a872045450a0cd61be31b7ef8f8aed01efdaf706b72dd198fa56d4db3c99f091ab3bf6e915acac5ef07d889f4bce420e13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13af2d8db5dec5598e0a1bb838bf9f9a344c98a5e6b903f5acd63d9e77f4cf94126fcc9971848d6117e2cab7f2bdd0cc9ec11145bac746caf293f016f11674ecd285b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ae33d3e43982f55470c28f3a713b505bb368487bd9b0d26bed053eeaf129c73fa7dafa9df9d206288f4e2c9c7a70fc01b82c7827bb4e8e1c98fa7151bbb9296cb0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18df3cc78b524872d1fe2665e817dcf5bcc25d7526f1c087b997a79568f2c36838c256fbc121fb2990ab3214d1c09ac493ec56b2289d42a2f0b796df98d5dc2b94deb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0bffced00210fd23871076db7633356ef35684cf5cdbbb3011135ccf46ef0ed6b4f46ff3fb5c9145162138ddf9d21bb7ce94c50802af3933b93a15513df5953c6e5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab54fa4929582394785bacf398ab9f19645caf0867e05f677672b3e49972ec00ea379d4275893219cdad2c29d23f75516f51b05646028e2a2f2fc92968c6d1949b16;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130ee9113fea7dc2b1402b40dc84a30341718b692df769964e150fea93afb9e65c5547a68e8240cf0441b0bc6dc9187a6b68c459f517a857af1435e884ce3a553a415;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1085379b948a285b46ed7a02f5071cb13c30bcdbdcbdcef4c4aa647cb61565848fcf75a6ffcccf56e12501ddc4f739cde9761a9a12259a2a2a843cb995a2c1f23e964;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1f5c13a1cecd69dd127f8e573d08474f3b90a7878a6a93ed98e9275c27d8256b28eea7e0b4474df8af207ec4b56c8b5679fec458c0d00a5b551b9eb584df8909057;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4a28e8e94b8bd312514cc4d35f7974a5585f780f871f971179af9c61dcd624f99bfffaad28bdb6627235d4c3b1fd98484b1c090177fc77bdd8615f9d13b35d1bf19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd686730ff39f0cb1d0e2c5060ab750b8180b1f6df537493b5b6c542432442cfde4e89ad9d25033b9ed6b8e2b7b4f6a1d48c242592cd63cfcd3ba64e16bb7402804fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h264a63a856a7e78fcff015824cf0ab295372db3cc81d83678bf089ac0f3855cf6b38ccf0eb3ad62944a4ffbf5fbb6c7f6102e1d20c44d5b2a4eedba8767bf9a708cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7912c3972054a0e9033101e99c0527c7ee3df04d70dac95c81602126d1ea69789b68da5efee93b78cc6e83512c138f126b93e42625d6bc53eed36fd8cdb8ebd3e34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13949638bb883de555cd5892e775d75a19f371c6a62aa81fa061ac6c3aae5af1d44717bd17daa7f507d748a754d9be775fa55e2bfb8e399b4f16f8bac2a6d8e59534f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3de7927e5990789ddb6dc00d78c01e37f38cef3b16593e2edbdd75a5e79cb01922c6597fcd32238efbd81c3bd913ebe7a108f776ca0b8c9c2865aa7fedb9f767126e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c324b80e1f7c2dbfafd8f6d1bfb49800f0d1fa53c581a30cf43e7fce184c74a6e1e569aa6cd79fcfc7a6767750b2bd7e38ed60f17fb5f1aea58fa6a2c4763103c88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb11bf31c45f8451c3730534e68793fd7d3dd181cc04e666a64319dd1a82c849a4ae9f3a569ad09236cb20d6b7a02bdce1acf06e57fd9b41e700973deec419c6cabf4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1730abf7445c40cd5987e4f1d76908dbb4b2b6d86c1bba78519f70a8c61a3fff7fc3156ac725ccaf9fc5ec905737ec582896e113e9bcc5f28b8f1b0291b97dbf265b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14cd70617c0226f50195e33cae9afab99def62ae079080c81a3df58cc16721925c412f077d6dd8d72f901a1daa6126f4c93b4cfa8ed5e1c5dd7c66fc34c27bebddb1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ad87091c987379fade55c84241f2f7ffae5e19224739c85dac6cc5dff9fb01d37be7b13ef2c046980855f9b7bcc1530a69abb1fab7d77299510b83a7d028a1d23ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6bc8d7799d07d0bf36c70397b3a418c453c4bd3b06be3c078b2a4fab25d2f4ca7126654fcfb6b4fe4e94dda1237d83829443b91411b75b5e97283b065f5a6ddfb98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10573c3ff90c2917f1a23ef673f3b78826e411cd7d195ac1a0a900fc861db7a5b107ec0f41718599b7bdb47f99b8484d664d2dfd1008c47ca5507f88df1b0addbe681;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c8a7410c13f29cc48ef14b3aee78c3df6c085bb3a41caf7d32f42af1deccc2de3d7776d7cabd55743fbd0cdf6df50ddad419604d31830204f42593c69a42ec81c32b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf32c60f38a6cba4f954c507146d6988a576ee49db496a1cf258024f16378be8b598f3f3c9cfcd390d85297322038004e5ca89eec0f739d816fcb13b7a275afdcf2e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f0c6db9dc0b5e9426e109bd6b86f03ea410b1d0149bd736e1a47cfb2fd73ed804726d3ecf13f13503fe9233cebc133cb00a6b9ed68b26d112fefb296b58c68c429e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136fff9b53e903d66e8903de5f45a4ea40a0559b52cdf399ef9ba2ba640529cb4db4cd5b3ee83ce68c36cc7e4f3edc61317da8054871b022347b35f81d0e8bec4cd8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f01162a84c8f6872274ecbe429725e66990376b794ba1f2b5924558534749fbe5c3da52522d41d8deae4d0d020f07fce3540c3ada448d375acd11be0aa62baa757d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fed93cfc5bf51866d822d7321e7fa0de25ee932f63982be020657a2f403c9f63f380b79089b4a03620d613f95a2bb54b520c530357ba10cecd308def1f65627b3315;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa44700760d9a391d4222344a0f1f9019d9a9c5e45ff7d5d8a376bcdae69d08d00aa079b0dbdb6a2ef83b6fff97fdb45ce2efab251e22276ebb102f519e2f7617cd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h538f5bdf8d029056169e68822b68f9744c4ab4e1533e1ae9da0be6be3006d91b75ba7fc52ed67ae0931d32a07cd4a1e641ee5a5cb9a59a2c4635577f53066fcf651f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129a0841815b1ff737eed336dc2c84014c191df2671640eb2f960a5c1d4a4521394209c8d9d955e570f54f5fab70ad8e4a311f68b403cdc45ef405dc50bc230bbd47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3e90a16e591421815e588078e1e5eb8732045815effd2297c1f2c53aeb4ef9a34162bfc2694e601cdaade61d8e756bee825415669267d128a90d35daf7bc11f8619;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb89eddfde428113ed570406761a1c33b435b23fe1b556a67ab16917c102e03fcd85ad8be9a77e6626dab938b6ca771c011dbe02eff2aa05e7fbaa0ee4a8fc4c702dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1036c900bf31122699881cf221536d910b467c7a23fe087640426e7edf6d79f8354e0fcd1713592108bcf80ded2dec6c42c450d7642b4789e0733a7a1f0bc0b06119a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6af6a5bd63644dac596342ec3c3f62865a1778349cfd2f7c67c84abf572e13b3e49275167f2d41cef7b69e7c16af74e51e4ae5c3f0c5a07a375e048ae3474beab006;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118c2b9657fa9d02a484f2f727c71cbff0e62b1b238ee7b9cba3796f0101e10b31dc6db4cf8d7a4c7be6dd042a6a96f59fc9f2b6dc20d504b4a2b0dc2d622dfde5330;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1baec98e9b12987e3d3ba0822e2fe72d4a7b733e81933aa86ab125ba9f46c12889295090e9014b9527dc53c5a71c8d218d9666498b801b6a3ad8e3bb78758b096d9de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ccd202e1a0dc7c8c8ba630918e7f568a8dabf2a5770b0b25375c14abc7a2a3718ccd4a300b1df7675c2dcc90769b7122eab683941fece0c2b60abd8d3cd19d2cf30;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1469e765de19a0b3516b4367091bbdedc215aa615b05b3142ff51d61e0bc4f1ab3a6a4248031db3ba053ad698453209cdb284b4b667055e8df3fdf1c321b693d310c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adcf73afaa6c1a5404e148d6c0384a0696ee234573842c4e1fbe1e8933497d4a822cb8c176a45db460a8fe04a3ffa4d7ac15101727b3de00d18e2798ce45994e065f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2da87368869c06b0c52a42c667958355e9c9d86d82873e90ce632d2a5f24c431b190ce713698942be0dc0155bc96eedbff5491852a8d0ddf841dabf1ec1d5524144;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6dbaac53025edc8c724e62c271097720c62088029cead5536d755c31b581c0736a497591f09e4fb3aa2b2380e83d54d257d80a1871786e260e5daf6f2910b8b117b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h839011c4336d570f129cbbadec0217933ef44fe2a36f68b6dda9ad2d33083dc910cc0e19743d278b8f75cbf7a78a281463811d6616baa695d8c6df71b255bf7508de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191fd502ce380893d9cc947993256d648be7b783d85366ac26b5c18e9ffcaea9ede404145481ded226da129344372be8478637334a247ca0b15299c521ca8ed5760a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c232b88c1b58a4bd90dadeab4c076c5c474fdd24da0ad4e94143155b9d037c328395b49327c19b10fee7f464b0c278445216e9137931fb1e324c55c5dfd08e76f2bd;
        #1
        $finish();
    end
endmodule
