module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    compressor_CLA128_32 compressor_CLA128_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
        src16 <= 128'h0;
        src17 <= 128'h0;
        src18 <= 128'h0;
        src19 <= 128'h0;
        src20 <= 128'h0;
        src21 <= 128'h0;
        src22 <= 128'h0;
        src23 <= 128'h0;
        src24 <= 128'h0;
        src25 <= 128'h0;
        src26 <= 128'h0;
        src27 <= 128'h0;
        src28 <= 128'h0;
        src29 <= 128'h0;
        src30 <= 128'h0;
        src31 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA128_32(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    input [127:0]src16,
    input [127:0]src17,
    input [127:0]src18,
    input [127:0]src19,
    input [127:0]src20,
    input [127:0]src21,
    input [127:0]src22,
    input [127:0]src23,
    input [127:0]src24,
    input [127:0]src25,
    input [127:0]src26,
    input [127:0]src27,
    input [127:0]src28,
    input [127:0]src29,
    input [127:0]src30,
    input [127:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [0:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], 1'h0, comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      input wire [127:0] src16,
      input wire [127:0] src17,
      input wire [127:0] src18,
      input wire [127:0] src19,
      input wire [127:0] src20,
      input wire [127:0] src21,
      input wire [127:0] src22,
      input wire [127:0] src23,
      input wire [127:0] src24,
      input wire [127:0] src25,
      input wire [127:0] src26,
      input wire [127:0] src27,
      input wire [127:0] src28,
      input wire [127:0] src29,
      input wire [127:0] src30,
      input wire [127:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [0:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [127:0] stage0_16;
   wire [127:0] stage0_17;
   wire [127:0] stage0_18;
   wire [127:0] stage0_19;
   wire [127:0] stage0_20;
   wire [127:0] stage0_21;
   wire [127:0] stage0_22;
   wire [127:0] stage0_23;
   wire [127:0] stage0_24;
   wire [127:0] stage0_25;
   wire [127:0] stage0_26;
   wire [127:0] stage0_27;
   wire [127:0] stage0_28;
   wire [127:0] stage0_29;
   wire [127:0] stage0_30;
   wire [127:0] stage0_31;
   wire [35:0] stage1_0;
   wire [39:0] stage1_1;
   wire [57:0] stage1_2;
   wire [58:0] stage1_3;
   wire [66:0] stage1_4;
   wire [62:0] stage1_5;
   wire [49:0] stage1_6;
   wire [69:0] stage1_7;
   wire [55:0] stage1_8;
   wire [60:0] stage1_9;
   wire [53:0] stage1_10;
   wire [57:0] stage1_11;
   wire [57:0] stage1_12;
   wire [60:0] stage1_13;
   wire [45:0] stage1_14;
   wire [46:0] stage1_15;
   wire [86:0] stage1_16;
   wire [62:0] stage1_17;
   wire [65:0] stage1_18;
   wire [42:0] stage1_19;
   wire [65:0] stage1_20;
   wire [64:0] stage1_21;
   wire [60:0] stage1_22;
   wire [43:0] stage1_23;
   wire [89:0] stage1_24;
   wire [69:0] stage1_25;
   wire [68:0] stage1_26;
   wire [55:0] stage1_27;
   wire [55:0] stage1_28;
   wire [56:0] stage1_29;
   wire [60:0] stage1_30;
   wire [70:0] stage1_31;
   wire [33:0] stage1_32;
   wire [15:0] stage1_33;
   wire [35:0] stage2_0;
   wire [19:0] stage2_1;
   wire [26:0] stage2_2;
   wire [33:0] stage2_3;
   wire [25:0] stage2_4;
   wire [30:0] stage2_5;
   wire [47:0] stage2_6;
   wire [19:0] stage2_7;
   wire [38:0] stage2_8;
   wire [22:0] stage2_9;
   wire [21:0] stage2_10;
   wire [26:0] stage2_11;
   wire [20:0] stage2_12;
   wire [34:0] stage2_13;
   wire [26:0] stage2_14;
   wire [22:0] stage2_15;
   wire [22:0] stage2_16;
   wire [48:0] stage2_17;
   wire [37:0] stage2_18;
   wire [20:0] stage2_19;
   wire [55:0] stage2_20;
   wire [20:0] stage2_21;
   wire [26:0] stage2_22;
   wire [33:0] stage2_23;
   wire [32:0] stage2_24;
   wire [46:0] stage2_25;
   wire [36:0] stage2_26;
   wire [30:0] stage2_27;
   wire [35:0] stage2_28;
   wire [31:0] stage2_29;
   wire [18:0] stage2_30;
   wire [33:0] stage2_31;
   wire [28:0] stage2_32;
   wire [17:0] stage2_33;
   wire [5:0] stage2_34;
   wire [1:0] stage2_35;
   wire [6:0] stage3_0;
   wire [12:0] stage3_1;
   wire [7:0] stage3_2;
   wire [12:0] stage3_3;
   wire [17:0] stage3_4;
   wire [8:0] stage3_5;
   wire [33:0] stage3_6;
   wire [12:0] stage3_7;
   wire [16:0] stage3_8;
   wire [8:0] stage3_9;
   wire [12:0] stage3_10;
   wire [13:0] stage3_11;
   wire [18:0] stage3_12;
   wire [10:0] stage3_13;
   wire [21:0] stage3_14;
   wire [11:0] stage3_15;
   wire [12:0] stage3_16;
   wire [24:0] stage3_17;
   wire [13:0] stage3_18;
   wire [25:0] stage3_19;
   wire [15:0] stage3_20;
   wire [13:0] stage3_21;
   wire [15:0] stage3_22;
   wire [10:0] stage3_23;
   wire [18:0] stage3_24;
   wire [13:0] stage3_25;
   wire [18:0] stage3_26;
   wire [13:0] stage3_27;
   wire [10:0] stage3_28;
   wire [17:0] stage3_29;
   wire [14:0] stage3_30;
   wire [8:0] stage3_31;
   wire [14:0] stage3_32;
   wire [20:0] stage3_33;
   wire [8:0] stage3_34;
   wire [1:0] stage3_35;
   wire [0:0] stage3_36;
   wire [1:0] stage4_0;
   wire [7:0] stage4_1;
   wire [3:0] stage4_2;
   wire [6:0] stage4_3;
   wire [7:0] stage4_4;
   wire [8:0] stage4_5;
   wire [10:0] stage4_6;
   wire [10:0] stage4_7;
   wire [10:0] stage4_8;
   wire [5:0] stage4_9;
   wire [6:0] stage4_10;
   wire [3:0] stage4_11;
   wire [8:0] stage4_12;
   wire [6:0] stage4_13;
   wire [5:0] stage4_14;
   wire [8:0] stage4_15;
   wire [6:0] stage4_16;
   wire [6:0] stage4_17;
   wire [11:0] stage4_18;
   wire [7:0] stage4_19;
   wire [6:0] stage4_20;
   wire [9:0] stage4_21;
   wire [6:0] stage4_22;
   wire [7:0] stage4_23;
   wire [10:0] stage4_24;
   wire [5:0] stage4_25;
   wire [12:0] stage4_26;
   wire [5:0] stage4_27;
   wire [6:0] stage4_28;
   wire [5:0] stage4_29;
   wire [4:0] stage4_30;
   wire [5:0] stage4_31;
   wire [6:0] stage4_32;
   wire [12:0] stage4_33;
   wire [11:0] stage4_34;
   wire [2:0] stage4_35;
   wire [1:0] stage4_36;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [4:0] stage5_3;
   wire [2:0] stage5_4;
   wire [3:0] stage5_5;
   wire [3:0] stage5_6;
   wire [3:0] stage5_7;
   wire [7:0] stage5_8;
   wire [2:0] stage5_9;
   wire [2:0] stage5_10;
   wire [5:0] stage5_11;
   wire [2:0] stage5_12;
   wire [2:0] stage5_13;
   wire [1:0] stage5_14;
   wire [6:0] stage5_15;
   wire [2:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [5:0] stage5_19;
   wire [2:0] stage5_20;
   wire [5:0] stage5_21;
   wire [2:0] stage5_22;
   wire [5:0] stage5_23;
   wire [4:0] stage5_24;
   wire [2:0] stage5_25;
   wire [3:0] stage5_26;
   wire [3:0] stage5_27;
   wire [3:0] stage5_28;
   wire [1:0] stage5_29;
   wire [6:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [3:0] stage5_33;
   wire [3:0] stage5_34;
   wire [3:0] stage5_35;
   wire [2:0] stage5_36;
   wire [1:0] stage5_37;
   wire [0:0] stage5_38;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [0:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [0:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[3]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[4]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[5]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[6]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[7]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc615_5 gpc20 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[48]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[49]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_1[50]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_1[51]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc1343_5 gpc36 (
      {stage0_2[104], stage0_2[105], stage0_2[106]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83]},
      {stage0_4[0], stage0_4[1], stage0_4[2]},
      {stage0_5[0]},
      {stage1_6[0],stage1_5[12],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_5[1]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[1],stage1_5[13],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage0_4[9]},
      {stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7]},
      {stage1_7[1],stage1_6[2],stage1_5[14],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[10]},
      {stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13]},
      {stage1_7[2],stage1_6[3],stage1_5[15],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[11]},
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage1_7[3],stage1_6[4],stage1_5[16],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[12]},
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage1_7[4],stage1_6[5],stage1_5[17],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[13]},
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage1_7[5],stage1_6[6],stage1_5[18],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage1_8[0],stage1_7[6],stage1_6[7],stage1_5[19],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12]},
      {stage1_8[1],stage1_7[7],stage1_6[8],stage1_5[20],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18]},
      {stage1_8[2],stage1_7[8],stage1_6[9],stage1_5[21],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37]},
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24]},
      {stage1_8[3],stage1_7[9],stage1_6[10],stage1_5[22],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30]},
      {stage1_8[4],stage1_7[10],stage1_6[11],stage1_5[23],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35], stage0_6[36]},
      {stage1_8[5],stage1_7[11],stage1_6[12],stage1_5[24],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage1_8[6],stage1_7[12],stage1_6[13],stage1_5[25],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage1_8[7],stage1_7[13],stage1_6[14],stage1_5[26],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53], stage0_6[54]},
      {stage1_8[8],stage1_7[14],stage1_6[15],stage1_5[27],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59], stage0_6[60]},
      {stage1_8[9],stage1_7[15],stage1_6[16],stage1_5[28],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65], stage0_6[66]},
      {stage1_8[10],stage1_7[16],stage1_6[17],stage1_5[29],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72]},
      {stage1_8[11],stage1_7[17],stage1_6[18],stage1_5[30],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage1_8[12],stage1_7[18],stage1_6[19],stage1_5[31],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83], stage0_6[84]},
      {stage1_8[13],stage1_7[19],stage1_6[20],stage1_5[32],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89], stage0_6[90]},
      {stage1_8[14],stage1_7[20],stage1_6[21],stage1_5[33],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95], stage0_6[96]},
      {stage1_8[15],stage1_7[21],stage1_6[22],stage1_5[34],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102]},
      {stage1_8[16],stage1_7[22],stage1_6[23],stage1_5[35],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage1_8[17],stage1_7[23],stage1_6[24],stage1_5[36],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[18],stage1_7[24],stage1_6[25],stage1_5[37]}
   );
   gpc606_5 gpc62 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[19],stage1_7[25],stage1_6[26],stage1_5[38]}
   );
   gpc606_5 gpc63 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[20],stage1_7[26],stage1_6[27],stage1_5[39]}
   );
   gpc606_5 gpc64 (
      {stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[21],stage1_7[27],stage1_6[28],stage1_5[40]}
   );
   gpc606_5 gpc65 (
      {stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[22],stage1_7[28],stage1_6[29],stage1_5[41]}
   );
   gpc606_5 gpc66 (
      {stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[23],stage1_7[29],stage1_6[30],stage1_5[42]}
   );
   gpc606_5 gpc67 (
      {stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[24],stage1_7[30],stage1_6[31],stage1_5[43]}
   );
   gpc606_5 gpc68 (
      {stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[25],stage1_7[31],stage1_6[32],stage1_5[44]}
   );
   gpc606_5 gpc69 (
      {stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[26],stage1_7[32],stage1_6[33],stage1_5[45]}
   );
   gpc606_5 gpc70 (
      {stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[27],stage1_7[33],stage1_6[34],stage1_5[46]}
   );
   gpc606_5 gpc71 (
      {stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[28],stage1_7[34],stage1_6[35],stage1_5[47]}
   );
   gpc606_5 gpc72 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[29],stage1_7[35],stage1_6[36],stage1_5[48]}
   );
   gpc606_5 gpc73 (
      {stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[30],stage1_7[36],stage1_6[37],stage1_5[49]}
   );
   gpc606_5 gpc74 (
      {stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[31],stage1_7[37],stage1_6[38],stage1_5[50]}
   );
   gpc615_5 gpc75 (
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage0_7[84]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[14],stage1_8[32],stage1_7[38],stage1_6[39]}
   );
   gpc615_5 gpc76 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[85]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[15],stage1_8[33],stage1_7[39],stage1_6[40]}
   );
   gpc615_5 gpc77 (
      {stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89], stage0_7[90]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[16],stage1_8[34],stage1_7[40]}
   );
   gpc615_5 gpc78 (
      {stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage0_8[13]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[3],stage1_9[17],stage1_8[35],stage1_7[41]}
   );
   gpc615_5 gpc79 (
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100]},
      {stage0_8[14]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[4],stage1_9[18],stage1_8[36],stage1_7[42]}
   );
   gpc207_4 gpc80 (
      {stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[3],stage1_10[5],stage1_9[19],stage1_8[37]}
   );
   gpc606_5 gpc81 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage1_12[0],stage1_11[4],stage1_10[6],stage1_9[20],stage1_8[38]}
   );
   gpc606_5 gpc82 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13]},
      {stage1_12[1],stage1_11[5],stage1_10[7],stage1_9[21],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19]},
      {stage1_12[2],stage1_11[6],stage1_10[8],stage1_9[22],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25]},
      {stage1_12[3],stage1_11[7],stage1_10[9],stage1_9[23],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31]},
      {stage1_12[4],stage1_11[8],stage1_10[10],stage1_9[24],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37]},
      {stage1_12[5],stage1_11[9],stage1_10[11],stage1_9[25],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage1_12[6],stage1_11[10],stage1_10[12],stage1_9[26],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69]},
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49]},
      {stage1_12[7],stage1_11[11],stage1_10[13],stage1_9[27],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54], stage0_10[55]},
      {stage1_12[8],stage1_11[12],stage1_10[14],stage1_9[28],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage1_12[9],stage1_11[13],stage1_10[15],stage1_9[29],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65], stage0_10[66], stage0_10[67]},
      {stage1_12[10],stage1_11[14],stage1_10[16],stage1_9[30],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93]},
      {stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71], stage0_10[72], stage0_10[73]},
      {stage1_12[11],stage1_11[15],stage1_10[17],stage1_9[31],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99]},
      {stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77], stage0_10[78], stage0_10[79]},
      {stage1_12[12],stage1_11[16],stage1_10[18],stage1_9[32],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105]},
      {stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83], stage0_10[84], stage0_10[85]},
      {stage1_12[13],stage1_11[17],stage1_10[19],stage1_9[33],stage1_8[51]}
   );
   gpc606_5 gpc95 (
      {stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89], stage0_10[90], stage0_10[91]},
      {stage1_12[14],stage1_11[18],stage1_10[20],stage1_9[34],stage1_8[52]}
   );
   gpc606_5 gpc96 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95], stage0_10[96], stage0_10[97]},
      {stage1_12[15],stage1_11[19],stage1_10[21],stage1_9[35],stage1_8[53]}
   );
   gpc615_5 gpc97 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[18]},
      {stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101], stage0_10[102], stage0_10[103]},
      {stage1_12[16],stage1_11[20],stage1_10[22],stage1_9[36],stage1_8[54]}
   );
   gpc615_5 gpc98 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[19]},
      {stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107], stage0_10[108], stage0_10[109]},
      {stage1_12[17],stage1_11[21],stage1_10[23],stage1_9[37],stage1_8[55]}
   );
   gpc606_5 gpc99 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[18],stage1_11[22],stage1_10[24],stage1_9[38]}
   );
   gpc606_5 gpc100 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[19],stage1_11[23],stage1_10[25],stage1_9[39]}
   );
   gpc606_5 gpc101 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[20],stage1_11[24],stage1_10[26],stage1_9[40]}
   );
   gpc606_5 gpc102 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[21],stage1_11[25],stage1_10[27],stage1_9[41]}
   );
   gpc606_5 gpc103 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[22],stage1_11[26],stage1_10[28],stage1_9[42]}
   );
   gpc606_5 gpc104 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[23],stage1_11[27],stage1_10[29],stage1_9[43]}
   );
   gpc606_5 gpc105 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[24],stage1_11[28],stage1_10[30],stage1_9[44]}
   );
   gpc606_5 gpc106 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[25],stage1_11[29],stage1_10[31],stage1_9[45]}
   );
   gpc606_5 gpc107 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[26],stage1_11[30],stage1_10[32],stage1_9[46]}
   );
   gpc606_5 gpc108 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[27],stage1_11[31],stage1_10[33],stage1_9[47]}
   );
   gpc606_5 gpc109 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[28],stage1_11[32],stage1_10[34],stage1_9[48]}
   );
   gpc606_5 gpc110 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[29],stage1_11[33],stage1_10[35],stage1_9[49]}
   );
   gpc606_5 gpc111 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[30],stage1_11[34],stage1_10[36],stage1_9[50]}
   );
   gpc606_5 gpc112 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[31],stage1_11[35],stage1_10[37],stage1_9[51]}
   );
   gpc606_5 gpc113 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[32],stage1_11[36],stage1_10[38],stage1_9[52]}
   );
   gpc606_5 gpc114 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[33],stage1_11[37],stage1_10[39],stage1_9[53]}
   );
   gpc606_5 gpc115 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[34],stage1_11[38],stage1_10[40],stage1_9[54]}
   );
   gpc606_5 gpc116 (
      {stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[17],stage1_12[35],stage1_11[39],stage1_10[41]}
   );
   gpc615_5 gpc117 (
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106]},
      {stage0_12[6]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[18],stage1_12[36],stage1_11[40]}
   );
   gpc615_5 gpc118 (
      {stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111]},
      {stage0_12[7]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[2],stage1_13[19],stage1_12[37],stage1_11[41]}
   );
   gpc606_5 gpc119 (
      {stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[2],stage1_14[3],stage1_13[20],stage1_12[38]}
   );
   gpc606_5 gpc120 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[3],stage1_14[4],stage1_13[21],stage1_12[39]}
   );
   gpc606_5 gpc121 (
      {stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[4],stage1_14[5],stage1_13[22],stage1_12[40]}
   );
   gpc606_5 gpc122 (
      {stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[5],stage1_14[6],stage1_13[23],stage1_12[41]}
   );
   gpc606_5 gpc123 (
      {stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[6],stage1_14[7],stage1_13[24],stage1_12[42]}
   );
   gpc606_5 gpc124 (
      {stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[7],stage1_14[8],stage1_13[25],stage1_12[43]}
   );
   gpc606_5 gpc125 (
      {stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[8],stage1_14[9],stage1_13[26],stage1_12[44]}
   );
   gpc606_5 gpc126 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[9],stage1_14[10],stage1_13[27],stage1_12[45]}
   );
   gpc606_5 gpc127 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[10],stage1_14[11],stage1_13[28],stage1_12[46]}
   );
   gpc606_5 gpc128 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[11],stage1_14[12],stage1_13[29],stage1_12[47]}
   );
   gpc606_5 gpc129 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[12],stage1_14[13],stage1_13[30],stage1_12[48]}
   );
   gpc606_5 gpc130 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[13],stage1_14[14],stage1_13[31],stage1_12[49]}
   );
   gpc606_5 gpc131 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[14],stage1_14[15],stage1_13[32],stage1_12[50]}
   );
   gpc606_5 gpc132 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[15],stage1_14[16],stage1_13[33],stage1_12[51]}
   );
   gpc606_5 gpc133 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[16],stage1_14[17],stage1_13[34],stage1_12[52]}
   );
   gpc606_5 gpc134 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[17],stage1_14[18],stage1_13[35],stage1_12[53]}
   );
   gpc606_5 gpc135 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[18],stage1_14[19],stage1_13[36],stage1_12[54]}
   );
   gpc606_5 gpc136 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[19],stage1_14[20],stage1_13[37],stage1_12[55]}
   );
   gpc606_5 gpc137 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[20],stage1_14[21],stage1_13[38],stage1_12[56]}
   );
   gpc606_5 gpc138 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[21],stage1_14[22],stage1_13[39],stage1_12[57]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[20],stage1_15[22],stage1_14[23],stage1_13[40]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[21],stage1_15[23],stage1_14[24],stage1_13[41]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[22],stage1_15[24],stage1_14[25],stage1_13[42]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[23],stage1_15[25],stage1_14[26],stage1_13[43]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[24],stage1_15[26],stage1_14[27],stage1_13[44]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[25],stage1_15[27],stage1_14[28],stage1_13[45]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[26],stage1_15[28],stage1_14[29],stage1_13[46]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[27],stage1_15[29],stage1_14[30],stage1_13[47]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[28],stage1_15[30],stage1_14[31],stage1_13[48]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[29],stage1_15[31],stage1_14[32],stage1_13[49]}
   );
   gpc606_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[30],stage1_15[32],stage1_14[33],stage1_13[50]}
   );
   gpc606_5 gpc150 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[31],stage1_15[33],stage1_14[34],stage1_13[51]}
   );
   gpc606_5 gpc151 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[32],stage1_15[34],stage1_14[35],stage1_13[52]}
   );
   gpc606_5 gpc152 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[33],stage1_15[35],stage1_14[36],stage1_13[53]}
   );
   gpc606_5 gpc153 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[34],stage1_15[36],stage1_14[37],stage1_13[54]}
   );
   gpc606_5 gpc154 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[35],stage1_15[37],stage1_14[38],stage1_13[55]}
   );
   gpc606_5 gpc155 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[36],stage1_15[38],stage1_14[39],stage1_13[56]}
   );
   gpc606_5 gpc156 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[37],stage1_15[39],stage1_14[40],stage1_13[57]}
   );
   gpc606_5 gpc157 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[38],stage1_15[40],stage1_14[41],stage1_13[58]}
   );
   gpc615_5 gpc158 (
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124]},
      {stage0_15[114]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[19],stage1_16[39],stage1_15[41],stage1_14[42]}
   );
   gpc615_5 gpc159 (
      {stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage0_16[6]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[1],stage1_17[20],stage1_16[40],stage1_15[42]}
   );
   gpc615_5 gpc160 (
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124]},
      {stage0_16[7]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[2],stage1_17[21],stage1_16[41],stage1_15[43]}
   );
   gpc606_5 gpc161 (
      {stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[2],stage1_18[3],stage1_17[22],stage1_16[42]}
   );
   gpc606_5 gpc162 (
      {stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[3],stage1_18[4],stage1_17[23],stage1_16[43]}
   );
   gpc606_5 gpc163 (
      {stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[4],stage1_18[5],stage1_17[24],stage1_16[44]}
   );
   gpc606_5 gpc164 (
      {stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[5],stage1_18[6],stage1_17[25],stage1_16[45]}
   );
   gpc606_5 gpc165 (
      {stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[6],stage1_18[7],stage1_17[26],stage1_16[46]}
   );
   gpc606_5 gpc166 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[7],stage1_18[8],stage1_17[27],stage1_16[47]}
   );
   gpc606_5 gpc167 (
      {stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[8],stage1_18[9],stage1_17[28],stage1_16[48]}
   );
   gpc606_5 gpc168 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[9],stage1_18[10],stage1_17[29],stage1_16[49]}
   );
   gpc606_5 gpc169 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[10],stage1_18[11],stage1_17[30],stage1_16[50]}
   );
   gpc606_5 gpc170 (
      {stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[11],stage1_18[12],stage1_17[31],stage1_16[51]}
   );
   gpc606_5 gpc171 (
      {stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[12],stage1_18[13],stage1_17[32],stage1_16[52]}
   );
   gpc606_5 gpc172 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[13],stage1_18[14],stage1_17[33],stage1_16[53]}
   );
   gpc606_5 gpc173 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[14],stage1_18[15],stage1_17[34],stage1_16[54]}
   );
   gpc606_5 gpc174 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[15],stage1_18[16],stage1_17[35],stage1_16[55]}
   );
   gpc606_5 gpc175 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[16],stage1_18[17],stage1_17[36],stage1_16[56]}
   );
   gpc606_5 gpc176 (
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[15],stage1_19[17],stage1_18[18],stage1_17[37]}
   );
   gpc606_5 gpc177 (
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[16],stage1_19[18],stage1_18[19],stage1_17[38]}
   );
   gpc606_5 gpc178 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[17],stage1_19[19],stage1_18[20],stage1_17[39]}
   );
   gpc606_5 gpc179 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[18],stage1_19[20],stage1_18[21],stage1_17[40]}
   );
   gpc606_5 gpc180 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[19],stage1_19[21],stage1_18[22],stage1_17[41]}
   );
   gpc606_5 gpc181 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[20],stage1_19[22],stage1_18[23],stage1_17[42]}
   );
   gpc606_5 gpc182 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[21],stage1_19[23],stage1_18[24],stage1_17[43]}
   );
   gpc606_5 gpc183 (
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[22],stage1_19[24],stage1_18[25],stage1_17[44]}
   );
   gpc606_5 gpc184 (
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[23],stage1_19[25],stage1_18[26],stage1_17[45]}
   );
   gpc606_5 gpc185 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[24],stage1_19[26],stage1_18[27],stage1_17[46]}
   );
   gpc606_5 gpc186 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[25],stage1_19[27],stage1_18[28],stage1_17[47]}
   );
   gpc606_5 gpc187 (
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[26],stage1_19[28],stage1_18[29],stage1_17[48]}
   );
   gpc606_5 gpc188 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[27],stage1_19[29],stage1_18[30],stage1_17[49]}
   );
   gpc606_5 gpc189 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[28],stage1_19[30],stage1_18[31],stage1_17[50]}
   );
   gpc606_5 gpc190 (
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[29],stage1_19[31],stage1_18[32],stage1_17[51]}
   );
   gpc606_5 gpc191 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[30],stage1_19[32],stage1_18[33],stage1_17[52]}
   );
   gpc606_5 gpc192 (
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[31],stage1_19[33],stage1_18[34],stage1_17[53]}
   );
   gpc606_5 gpc193 (
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[32],stage1_19[34],stage1_18[35],stage1_17[54]}
   );
   gpc615_5 gpc194 (
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94]},
      {stage0_19[108]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[18],stage1_20[33],stage1_19[35],stage1_18[36]}
   );
   gpc615_5 gpc195 (
      {stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99]},
      {stage0_19[109]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[19],stage1_20[34],stage1_19[36],stage1_18[37]}
   );
   gpc615_5 gpc196 (
      {stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113], stage0_19[114]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[20],stage1_20[35],stage1_19[37]}
   );
   gpc615_5 gpc197 (
      {stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage0_20[13]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[3],stage1_21[21],stage1_20[36],stage1_19[38]}
   );
   gpc615_5 gpc198 (
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124]},
      {stage0_20[14]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[4],stage1_21[22],stage1_20[37],stage1_19[39]}
   );
   gpc606_5 gpc199 (
      {stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[3],stage1_22[5],stage1_21[23],stage1_20[38]}
   );
   gpc606_5 gpc200 (
      {stage0_20[21], stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[4],stage1_22[6],stage1_21[24],stage1_20[39]}
   );
   gpc606_5 gpc201 (
      {stage0_20[27], stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[5],stage1_22[7],stage1_21[25],stage1_20[40]}
   );
   gpc606_5 gpc202 (
      {stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[6],stage1_22[8],stage1_21[26],stage1_20[41]}
   );
   gpc606_5 gpc203 (
      {stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43], stage0_20[44]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[7],stage1_22[9],stage1_21[27],stage1_20[42]}
   );
   gpc606_5 gpc204 (
      {stage0_20[45], stage0_20[46], stage0_20[47], stage0_20[48], stage0_20[49], stage0_20[50]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[8],stage1_22[10],stage1_21[28],stage1_20[43]}
   );
   gpc606_5 gpc205 (
      {stage0_20[51], stage0_20[52], stage0_20[53], stage0_20[54], stage0_20[55], stage0_20[56]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[9],stage1_22[11],stage1_21[29],stage1_20[44]}
   );
   gpc606_5 gpc206 (
      {stage0_20[57], stage0_20[58], stage0_20[59], stage0_20[60], stage0_20[61], stage0_20[62]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[10],stage1_22[12],stage1_21[30],stage1_20[45]}
   );
   gpc606_5 gpc207 (
      {stage0_20[63], stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[11],stage1_22[13],stage1_21[31],stage1_20[46]}
   );
   gpc606_5 gpc208 (
      {stage0_20[69], stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[12],stage1_22[14],stage1_21[32],stage1_20[47]}
   );
   gpc606_5 gpc209 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[13],stage1_22[15],stage1_21[33],stage1_20[48]}
   );
   gpc606_5 gpc210 (
      {stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[14],stage1_22[16],stage1_21[34],stage1_20[49]}
   );
   gpc606_5 gpc211 (
      {stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[15],stage1_22[17],stage1_21[35],stage1_20[50]}
   );
   gpc606_5 gpc212 (
      {stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[16],stage1_22[18],stage1_21[36],stage1_20[51]}
   );
   gpc606_5 gpc213 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[17],stage1_22[19],stage1_21[37],stage1_20[52]}
   );
   gpc606_5 gpc214 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[18],stage1_22[20],stage1_21[38],stage1_20[53]}
   );
   gpc606_5 gpc215 (
      {stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[19],stage1_22[21],stage1_21[39],stage1_20[54]}
   );
   gpc606_5 gpc216 (
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[17],stage1_23[20],stage1_22[22],stage1_21[40]}
   );
   gpc606_5 gpc217 (
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[18],stage1_23[21],stage1_22[23],stage1_21[41]}
   );
   gpc606_5 gpc218 (
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[19],stage1_23[22],stage1_22[24],stage1_21[42]}
   );
   gpc606_5 gpc219 (
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[20],stage1_23[23],stage1_22[25],stage1_21[43]}
   );
   gpc606_5 gpc220 (
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[21],stage1_23[24],stage1_22[26],stage1_21[44]}
   );
   gpc606_5 gpc221 (
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[22],stage1_23[25],stage1_22[27],stage1_21[45]}
   );
   gpc606_5 gpc222 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[23],stage1_23[26],stage1_22[28],stage1_21[46]}
   );
   gpc606_5 gpc223 (
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[24],stage1_23[27],stage1_22[29],stage1_21[47]}
   );
   gpc606_5 gpc224 (
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[25],stage1_23[28],stage1_22[30],stage1_21[48]}
   );
   gpc606_5 gpc225 (
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[26],stage1_23[29],stage1_22[31],stage1_21[49]}
   );
   gpc606_5 gpc226 (
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[27],stage1_23[30],stage1_22[32],stage1_21[50]}
   );
   gpc606_5 gpc227 (
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[28],stage1_23[31],stage1_22[33],stage1_21[51]}
   );
   gpc606_5 gpc228 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[29],stage1_23[32],stage1_22[34],stage1_21[52]}
   );
   gpc606_5 gpc229 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[30],stage1_23[33],stage1_22[35],stage1_21[53]}
   );
   gpc606_5 gpc230 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[31],stage1_23[34],stage1_22[36],stage1_21[54]}
   );
   gpc606_5 gpc231 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[32],stage1_23[35],stage1_22[37],stage1_21[55]}
   );
   gpc606_5 gpc232 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[33],stage1_23[36],stage1_22[38],stage1_21[56]}
   );
   gpc615_5 gpc233 (
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106]},
      {stage0_23[102]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[17],stage1_24[34],stage1_23[37],stage1_22[39]}
   );
   gpc606_5 gpc234 (
      {stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[18],stage1_24[35],stage1_23[38]}
   );
   gpc606_5 gpc235 (
      {stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[2],stage1_25[19],stage1_24[36],stage1_23[39]}
   );
   gpc606_5 gpc236 (
      {stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[3],stage1_25[20],stage1_24[37],stage1_23[40]}
   );
   gpc615_5 gpc237 (
      {stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage0_24[6]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[4],stage1_25[21],stage1_24[38],stage1_23[41]}
   );
   gpc606_5 gpc238 (
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[4],stage1_26[5],stage1_25[22],stage1_24[39]}
   );
   gpc606_5 gpc239 (
      {stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[5],stage1_26[6],stage1_25[23],stage1_24[40]}
   );
   gpc606_5 gpc240 (
      {stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[6],stage1_26[7],stage1_25[24],stage1_24[41]}
   );
   gpc606_5 gpc241 (
      {stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[7],stage1_26[8],stage1_25[25],stage1_24[42]}
   );
   gpc606_5 gpc242 (
      {stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[8],stage1_26[9],stage1_25[26],stage1_24[43]}
   );
   gpc606_5 gpc243 (
      {stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[9],stage1_26[10],stage1_25[27],stage1_24[44]}
   );
   gpc606_5 gpc244 (
      {stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47], stage0_24[48]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[10],stage1_26[11],stage1_25[28],stage1_24[45]}
   );
   gpc606_5 gpc245 (
      {stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53], stage0_24[54]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[11],stage1_26[12],stage1_25[29],stage1_24[46]}
   );
   gpc606_5 gpc246 (
      {stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59], stage0_24[60]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[12],stage1_26[13],stage1_25[30],stage1_24[47]}
   );
   gpc606_5 gpc247 (
      {stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65], stage0_24[66]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[13],stage1_26[14],stage1_25[31],stage1_24[48]}
   );
   gpc606_5 gpc248 (
      {stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71], stage0_24[72]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[14],stage1_26[15],stage1_25[32],stage1_24[49]}
   );
   gpc606_5 gpc249 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[15],stage1_26[16],stage1_25[33],stage1_24[50]}
   );
   gpc606_5 gpc250 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[16],stage1_26[17],stage1_25[34],stage1_24[51]}
   );
   gpc606_5 gpc251 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[17],stage1_26[18],stage1_25[35],stage1_24[52]}
   );
   gpc606_5 gpc252 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[14],stage1_27[18],stage1_26[19],stage1_25[36]}
   );
   gpc606_5 gpc253 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[15],stage1_27[19],stage1_26[20],stage1_25[37]}
   );
   gpc606_5 gpc254 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[16],stage1_27[20],stage1_26[21],stage1_25[38]}
   );
   gpc606_5 gpc255 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[17],stage1_27[21],stage1_26[22],stage1_25[39]}
   );
   gpc606_5 gpc256 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[18],stage1_27[22],stage1_26[23],stage1_25[40]}
   );
   gpc606_5 gpc257 (
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[19],stage1_27[23],stage1_26[24],stage1_25[41]}
   );
   gpc606_5 gpc258 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[20],stage1_27[24],stage1_26[25],stage1_25[42]}
   );
   gpc606_5 gpc259 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[21],stage1_27[25],stage1_26[26],stage1_25[43]}
   );
   gpc606_5 gpc260 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[22],stage1_27[26],stage1_26[27],stage1_25[44]}
   );
   gpc606_5 gpc261 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[23],stage1_27[27],stage1_26[28],stage1_25[45]}
   );
   gpc606_5 gpc262 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[24],stage1_27[28],stage1_26[29],stage1_25[46]}
   );
   gpc606_5 gpc263 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[25],stage1_27[29],stage1_26[30],stage1_25[47]}
   );
   gpc606_5 gpc264 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[26],stage1_27[30],stage1_26[31],stage1_25[48]}
   );
   gpc606_5 gpc265 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[27],stage1_27[31],stage1_26[32],stage1_25[49]}
   );
   gpc615_5 gpc266 (
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88]},
      {stage0_27[84]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[14],stage1_28[28],stage1_27[32],stage1_26[33]}
   );
   gpc615_5 gpc267 (
      {stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93]},
      {stage0_27[85]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[15],stage1_28[29],stage1_27[33],stage1_26[34]}
   );
   gpc615_5 gpc268 (
      {stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89], stage0_27[90]},
      {stage0_28[12]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[2],stage1_29[16],stage1_28[30],stage1_27[34]}
   );
   gpc615_5 gpc269 (
      {stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage0_28[13]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[3],stage1_29[17],stage1_28[31],stage1_27[35]}
   );
   gpc615_5 gpc270 (
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100]},
      {stage0_28[14]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[4],stage1_29[18],stage1_28[32],stage1_27[36]}
   );
   gpc615_5 gpc271 (
      {stage0_27[101], stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105]},
      {stage0_28[15]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[5],stage1_29[19],stage1_28[33],stage1_27[37]}
   );
   gpc615_5 gpc272 (
      {stage0_27[106], stage0_27[107], stage0_27[108], stage0_27[109], stage0_27[110]},
      {stage0_28[16]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[6],stage1_29[20],stage1_28[34],stage1_27[38]}
   );
   gpc606_5 gpc273 (
      {stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[5],stage1_30[7],stage1_29[21],stage1_28[35]}
   );
   gpc606_5 gpc274 (
      {stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[6],stage1_30[8],stage1_29[22],stage1_28[36]}
   );
   gpc606_5 gpc275 (
      {stage0_28[29], stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[7],stage1_30[9],stage1_29[23],stage1_28[37]}
   );
   gpc606_5 gpc276 (
      {stage0_28[35], stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[8],stage1_30[10],stage1_29[24],stage1_28[38]}
   );
   gpc606_5 gpc277 (
      {stage0_28[41], stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[9],stage1_30[11],stage1_29[25],stage1_28[39]}
   );
   gpc606_5 gpc278 (
      {stage0_28[47], stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[10],stage1_30[12],stage1_29[26],stage1_28[40]}
   );
   gpc606_5 gpc279 (
      {stage0_28[53], stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[11],stage1_30[13],stage1_29[27],stage1_28[41]}
   );
   gpc606_5 gpc280 (
      {stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[12],stage1_30[14],stage1_29[28],stage1_28[42]}
   );
   gpc606_5 gpc281 (
      {stage0_28[65], stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[13],stage1_30[15],stage1_29[29],stage1_28[43]}
   );
   gpc606_5 gpc282 (
      {stage0_28[71], stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[14],stage1_30[16],stage1_29[30],stage1_28[44]}
   );
   gpc606_5 gpc283 (
      {stage0_28[77], stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[15],stage1_30[17],stage1_29[31],stage1_28[45]}
   );
   gpc606_5 gpc284 (
      {stage0_28[83], stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[16],stage1_30[18],stage1_29[32],stage1_28[46]}
   );
   gpc606_5 gpc285 (
      {stage0_28[89], stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[17],stage1_30[19],stage1_29[33],stage1_28[47]}
   );
   gpc606_5 gpc286 (
      {stage0_28[95], stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[18],stage1_30[20],stage1_29[34],stage1_28[48]}
   );
   gpc606_5 gpc287 (
      {stage0_28[101], stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[19],stage1_30[21],stage1_29[35],stage1_28[49]}
   );
   gpc606_5 gpc288 (
      {stage0_28[107], stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[20],stage1_30[22],stage1_29[36],stage1_28[50]}
   );
   gpc606_5 gpc289 (
      {stage0_28[113], stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[21],stage1_30[23],stage1_29[37],stage1_28[51]}
   );
   gpc606_5 gpc290 (
      {stage0_28[119], stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[22],stage1_30[24],stage1_29[38],stage1_28[52]}
   );
   gpc606_5 gpc291 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[18],stage1_31[23],stage1_30[25],stage1_29[39]}
   );
   gpc606_5 gpc292 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[19],stage1_31[24],stage1_30[26],stage1_29[40]}
   );
   gpc606_5 gpc293 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[20],stage1_31[25],stage1_30[27],stage1_29[41]}
   );
   gpc606_5 gpc294 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[21],stage1_31[26],stage1_30[28],stage1_29[42]}
   );
   gpc606_5 gpc295 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[22],stage1_31[27],stage1_30[29],stage1_29[43]}
   );
   gpc606_5 gpc296 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[23],stage1_31[28],stage1_30[30],stage1_29[44]}
   );
   gpc606_5 gpc297 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[24],stage1_31[29],stage1_30[31],stage1_29[45]}
   );
   gpc606_5 gpc298 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[25],stage1_31[30],stage1_30[32],stage1_29[46]}
   );
   gpc606_5 gpc299 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[26],stage1_31[31],stage1_30[33],stage1_29[47]}
   );
   gpc606_5 gpc300 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[27],stage1_31[32],stage1_30[34],stage1_29[48]}
   );
   gpc606_5 gpc301 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[28],stage1_31[33],stage1_30[35],stage1_29[49]}
   );
   gpc606_5 gpc302 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[29],stage1_31[34],stage1_30[36],stage1_29[50]}
   );
   gpc606_5 gpc303 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[30],stage1_31[35],stage1_30[37],stage1_29[51]}
   );
   gpc606_5 gpc304 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[31],stage1_31[36],stage1_30[38],stage1_29[52]}
   );
   gpc606_5 gpc305 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[32],stage1_31[37],stage1_30[39],stage1_29[53]}
   );
   gpc606_5 gpc306 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[33],stage1_31[38],stage1_30[40],stage1_29[54]}
   );
   gpc1_1 gpc307 (
      {stage0_0[116]},
      {stage1_0[24]}
   );
   gpc1_1 gpc308 (
      {stage0_0[117]},
      {stage1_0[25]}
   );
   gpc1_1 gpc309 (
      {stage0_0[118]},
      {stage1_0[26]}
   );
   gpc1_1 gpc310 (
      {stage0_0[119]},
      {stage1_0[27]}
   );
   gpc1_1 gpc311 (
      {stage0_0[120]},
      {stage1_0[28]}
   );
   gpc1_1 gpc312 (
      {stage0_0[121]},
      {stage1_0[29]}
   );
   gpc1_1 gpc313 (
      {stage0_0[122]},
      {stage1_0[30]}
   );
   gpc1_1 gpc314 (
      {stage0_0[123]},
      {stage1_0[31]}
   );
   gpc1_1 gpc315 (
      {stage0_0[124]},
      {stage1_0[32]}
   );
   gpc1_1 gpc316 (
      {stage0_0[125]},
      {stage1_0[33]}
   );
   gpc1_1 gpc317 (
      {stage0_0[126]},
      {stage1_0[34]}
   );
   gpc1_1 gpc318 (
      {stage0_0[127]},
      {stage1_0[35]}
   );
   gpc1_1 gpc319 (
      {stage0_1[124]},
      {stage1_1[36]}
   );
   gpc1_1 gpc320 (
      {stage0_1[125]},
      {stage1_1[37]}
   );
   gpc1_1 gpc321 (
      {stage0_1[126]},
      {stage1_1[38]}
   );
   gpc1_1 gpc322 (
      {stage0_1[127]},
      {stage1_1[39]}
   );
   gpc1_1 gpc323 (
      {stage0_2[107]},
      {stage1_2[37]}
   );
   gpc1_1 gpc324 (
      {stage0_2[108]},
      {stage1_2[38]}
   );
   gpc1_1 gpc325 (
      {stage0_2[109]},
      {stage1_2[39]}
   );
   gpc1_1 gpc326 (
      {stage0_2[110]},
      {stage1_2[40]}
   );
   gpc1_1 gpc327 (
      {stage0_2[111]},
      {stage1_2[41]}
   );
   gpc1_1 gpc328 (
      {stage0_2[112]},
      {stage1_2[42]}
   );
   gpc1_1 gpc329 (
      {stage0_2[113]},
      {stage1_2[43]}
   );
   gpc1_1 gpc330 (
      {stage0_2[114]},
      {stage1_2[44]}
   );
   gpc1_1 gpc331 (
      {stage0_2[115]},
      {stage1_2[45]}
   );
   gpc1_1 gpc332 (
      {stage0_2[116]},
      {stage1_2[46]}
   );
   gpc1_1 gpc333 (
      {stage0_2[117]},
      {stage1_2[47]}
   );
   gpc1_1 gpc334 (
      {stage0_2[118]},
      {stage1_2[48]}
   );
   gpc1_1 gpc335 (
      {stage0_2[119]},
      {stage1_2[49]}
   );
   gpc1_1 gpc336 (
      {stage0_2[120]},
      {stage1_2[50]}
   );
   gpc1_1 gpc337 (
      {stage0_2[121]},
      {stage1_2[51]}
   );
   gpc1_1 gpc338 (
      {stage0_2[122]},
      {stage1_2[52]}
   );
   gpc1_1 gpc339 (
      {stage0_2[123]},
      {stage1_2[53]}
   );
   gpc1_1 gpc340 (
      {stage0_2[124]},
      {stage1_2[54]}
   );
   gpc1_1 gpc341 (
      {stage0_2[125]},
      {stage1_2[55]}
   );
   gpc1_1 gpc342 (
      {stage0_2[126]},
      {stage1_2[56]}
   );
   gpc1_1 gpc343 (
      {stage0_2[127]},
      {stage1_2[57]}
   );
   gpc1_1 gpc344 (
      {stage0_3[112]},
      {stage1_3[43]}
   );
   gpc1_1 gpc345 (
      {stage0_3[113]},
      {stage1_3[44]}
   );
   gpc1_1 gpc346 (
      {stage0_3[114]},
      {stage1_3[45]}
   );
   gpc1_1 gpc347 (
      {stage0_3[115]},
      {stage1_3[46]}
   );
   gpc1_1 gpc348 (
      {stage0_3[116]},
      {stage1_3[47]}
   );
   gpc1_1 gpc349 (
      {stage0_3[117]},
      {stage1_3[48]}
   );
   gpc1_1 gpc350 (
      {stage0_3[118]},
      {stage1_3[49]}
   );
   gpc1_1 gpc351 (
      {stage0_3[119]},
      {stage1_3[50]}
   );
   gpc1_1 gpc352 (
      {stage0_3[120]},
      {stage1_3[51]}
   );
   gpc1_1 gpc353 (
      {stage0_3[121]},
      {stage1_3[52]}
   );
   gpc1_1 gpc354 (
      {stage0_3[122]},
      {stage1_3[53]}
   );
   gpc1_1 gpc355 (
      {stage0_3[123]},
      {stage1_3[54]}
   );
   gpc1_1 gpc356 (
      {stage0_3[124]},
      {stage1_3[55]}
   );
   gpc1_1 gpc357 (
      {stage0_3[125]},
      {stage1_3[56]}
   );
   gpc1_1 gpc358 (
      {stage0_3[126]},
      {stage1_3[57]}
   );
   gpc1_1 gpc359 (
      {stage0_3[127]},
      {stage1_3[58]}
   );
   gpc1_1 gpc360 (
      {stage0_4[122]},
      {stage1_4[61]}
   );
   gpc1_1 gpc361 (
      {stage0_4[123]},
      {stage1_4[62]}
   );
   gpc1_1 gpc362 (
      {stage0_4[124]},
      {stage1_4[63]}
   );
   gpc1_1 gpc363 (
      {stage0_4[125]},
      {stage1_4[64]}
   );
   gpc1_1 gpc364 (
      {stage0_4[126]},
      {stage1_4[65]}
   );
   gpc1_1 gpc365 (
      {stage0_4[127]},
      {stage1_4[66]}
   );
   gpc1_1 gpc366 (
      {stage0_5[116]},
      {stage1_5[51]}
   );
   gpc1_1 gpc367 (
      {stage0_5[117]},
      {stage1_5[52]}
   );
   gpc1_1 gpc368 (
      {stage0_5[118]},
      {stage1_5[53]}
   );
   gpc1_1 gpc369 (
      {stage0_5[119]},
      {stage1_5[54]}
   );
   gpc1_1 gpc370 (
      {stage0_5[120]},
      {stage1_5[55]}
   );
   gpc1_1 gpc371 (
      {stage0_5[121]},
      {stage1_5[56]}
   );
   gpc1_1 gpc372 (
      {stage0_5[122]},
      {stage1_5[57]}
   );
   gpc1_1 gpc373 (
      {stage0_5[123]},
      {stage1_5[58]}
   );
   gpc1_1 gpc374 (
      {stage0_5[124]},
      {stage1_5[59]}
   );
   gpc1_1 gpc375 (
      {stage0_5[125]},
      {stage1_5[60]}
   );
   gpc1_1 gpc376 (
      {stage0_5[126]},
      {stage1_5[61]}
   );
   gpc1_1 gpc377 (
      {stage0_5[127]},
      {stage1_5[62]}
   );
   gpc1_1 gpc378 (
      {stage0_6[119]},
      {stage1_6[41]}
   );
   gpc1_1 gpc379 (
      {stage0_6[120]},
      {stage1_6[42]}
   );
   gpc1_1 gpc380 (
      {stage0_6[121]},
      {stage1_6[43]}
   );
   gpc1_1 gpc381 (
      {stage0_6[122]},
      {stage1_6[44]}
   );
   gpc1_1 gpc382 (
      {stage0_6[123]},
      {stage1_6[45]}
   );
   gpc1_1 gpc383 (
      {stage0_6[124]},
      {stage1_6[46]}
   );
   gpc1_1 gpc384 (
      {stage0_6[125]},
      {stage1_6[47]}
   );
   gpc1_1 gpc385 (
      {stage0_6[126]},
      {stage1_6[48]}
   );
   gpc1_1 gpc386 (
      {stage0_6[127]},
      {stage1_6[49]}
   );
   gpc1_1 gpc387 (
      {stage0_7[101]},
      {stage1_7[43]}
   );
   gpc1_1 gpc388 (
      {stage0_7[102]},
      {stage1_7[44]}
   );
   gpc1_1 gpc389 (
      {stage0_7[103]},
      {stage1_7[45]}
   );
   gpc1_1 gpc390 (
      {stage0_7[104]},
      {stage1_7[46]}
   );
   gpc1_1 gpc391 (
      {stage0_7[105]},
      {stage1_7[47]}
   );
   gpc1_1 gpc392 (
      {stage0_7[106]},
      {stage1_7[48]}
   );
   gpc1_1 gpc393 (
      {stage0_7[107]},
      {stage1_7[49]}
   );
   gpc1_1 gpc394 (
      {stage0_7[108]},
      {stage1_7[50]}
   );
   gpc1_1 gpc395 (
      {stage0_7[109]},
      {stage1_7[51]}
   );
   gpc1_1 gpc396 (
      {stage0_7[110]},
      {stage1_7[52]}
   );
   gpc1_1 gpc397 (
      {stage0_7[111]},
      {stage1_7[53]}
   );
   gpc1_1 gpc398 (
      {stage0_7[112]},
      {stage1_7[54]}
   );
   gpc1_1 gpc399 (
      {stage0_7[113]},
      {stage1_7[55]}
   );
   gpc1_1 gpc400 (
      {stage0_7[114]},
      {stage1_7[56]}
   );
   gpc1_1 gpc401 (
      {stage0_7[115]},
      {stage1_7[57]}
   );
   gpc1_1 gpc402 (
      {stage0_7[116]},
      {stage1_7[58]}
   );
   gpc1_1 gpc403 (
      {stage0_7[117]},
      {stage1_7[59]}
   );
   gpc1_1 gpc404 (
      {stage0_7[118]},
      {stage1_7[60]}
   );
   gpc1_1 gpc405 (
      {stage0_7[119]},
      {stage1_7[61]}
   );
   gpc1_1 gpc406 (
      {stage0_7[120]},
      {stage1_7[62]}
   );
   gpc1_1 gpc407 (
      {stage0_7[121]},
      {stage1_7[63]}
   );
   gpc1_1 gpc408 (
      {stage0_7[122]},
      {stage1_7[64]}
   );
   gpc1_1 gpc409 (
      {stage0_7[123]},
      {stage1_7[65]}
   );
   gpc1_1 gpc410 (
      {stage0_7[124]},
      {stage1_7[66]}
   );
   gpc1_1 gpc411 (
      {stage0_7[125]},
      {stage1_7[67]}
   );
   gpc1_1 gpc412 (
      {stage0_7[126]},
      {stage1_7[68]}
   );
   gpc1_1 gpc413 (
      {stage0_7[127]},
      {stage1_7[69]}
   );
   gpc1_1 gpc414 (
      {stage0_9[122]},
      {stage1_9[55]}
   );
   gpc1_1 gpc415 (
      {stage0_9[123]},
      {stage1_9[56]}
   );
   gpc1_1 gpc416 (
      {stage0_9[124]},
      {stage1_9[57]}
   );
   gpc1_1 gpc417 (
      {stage0_9[125]},
      {stage1_9[58]}
   );
   gpc1_1 gpc418 (
      {stage0_9[126]},
      {stage1_9[59]}
   );
   gpc1_1 gpc419 (
      {stage0_9[127]},
      {stage1_9[60]}
   );
   gpc1_1 gpc420 (
      {stage0_10[116]},
      {stage1_10[42]}
   );
   gpc1_1 gpc421 (
      {stage0_10[117]},
      {stage1_10[43]}
   );
   gpc1_1 gpc422 (
      {stage0_10[118]},
      {stage1_10[44]}
   );
   gpc1_1 gpc423 (
      {stage0_10[119]},
      {stage1_10[45]}
   );
   gpc1_1 gpc424 (
      {stage0_10[120]},
      {stage1_10[46]}
   );
   gpc1_1 gpc425 (
      {stage0_10[121]},
      {stage1_10[47]}
   );
   gpc1_1 gpc426 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc427 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc428 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc429 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc430 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc431 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc432 (
      {stage0_11[112]},
      {stage1_11[42]}
   );
   gpc1_1 gpc433 (
      {stage0_11[113]},
      {stage1_11[43]}
   );
   gpc1_1 gpc434 (
      {stage0_11[114]},
      {stage1_11[44]}
   );
   gpc1_1 gpc435 (
      {stage0_11[115]},
      {stage1_11[45]}
   );
   gpc1_1 gpc436 (
      {stage0_11[116]},
      {stage1_11[46]}
   );
   gpc1_1 gpc437 (
      {stage0_11[117]},
      {stage1_11[47]}
   );
   gpc1_1 gpc438 (
      {stage0_11[118]},
      {stage1_11[48]}
   );
   gpc1_1 gpc439 (
      {stage0_11[119]},
      {stage1_11[49]}
   );
   gpc1_1 gpc440 (
      {stage0_11[120]},
      {stage1_11[50]}
   );
   gpc1_1 gpc441 (
      {stage0_11[121]},
      {stage1_11[51]}
   );
   gpc1_1 gpc442 (
      {stage0_11[122]},
      {stage1_11[52]}
   );
   gpc1_1 gpc443 (
      {stage0_11[123]},
      {stage1_11[53]}
   );
   gpc1_1 gpc444 (
      {stage0_11[124]},
      {stage1_11[54]}
   );
   gpc1_1 gpc445 (
      {stage0_11[125]},
      {stage1_11[55]}
   );
   gpc1_1 gpc446 (
      {stage0_11[126]},
      {stage1_11[56]}
   );
   gpc1_1 gpc447 (
      {stage0_11[127]},
      {stage1_11[57]}
   );
   gpc1_1 gpc448 (
      {stage0_13[126]},
      {stage1_13[59]}
   );
   gpc1_1 gpc449 (
      {stage0_13[127]},
      {stage1_13[60]}
   );
   gpc1_1 gpc450 (
      {stage0_14[125]},
      {stage1_14[43]}
   );
   gpc1_1 gpc451 (
      {stage0_14[126]},
      {stage1_14[44]}
   );
   gpc1_1 gpc452 (
      {stage0_14[127]},
      {stage1_14[45]}
   );
   gpc1_1 gpc453 (
      {stage0_15[125]},
      {stage1_15[44]}
   );
   gpc1_1 gpc454 (
      {stage0_15[126]},
      {stage1_15[45]}
   );
   gpc1_1 gpc455 (
      {stage0_15[127]},
      {stage1_15[46]}
   );
   gpc1_1 gpc456 (
      {stage0_16[98]},
      {stage1_16[57]}
   );
   gpc1_1 gpc457 (
      {stage0_16[99]},
      {stage1_16[58]}
   );
   gpc1_1 gpc458 (
      {stage0_16[100]},
      {stage1_16[59]}
   );
   gpc1_1 gpc459 (
      {stage0_16[101]},
      {stage1_16[60]}
   );
   gpc1_1 gpc460 (
      {stage0_16[102]},
      {stage1_16[61]}
   );
   gpc1_1 gpc461 (
      {stage0_16[103]},
      {stage1_16[62]}
   );
   gpc1_1 gpc462 (
      {stage0_16[104]},
      {stage1_16[63]}
   );
   gpc1_1 gpc463 (
      {stage0_16[105]},
      {stage1_16[64]}
   );
   gpc1_1 gpc464 (
      {stage0_16[106]},
      {stage1_16[65]}
   );
   gpc1_1 gpc465 (
      {stage0_16[107]},
      {stage1_16[66]}
   );
   gpc1_1 gpc466 (
      {stage0_16[108]},
      {stage1_16[67]}
   );
   gpc1_1 gpc467 (
      {stage0_16[109]},
      {stage1_16[68]}
   );
   gpc1_1 gpc468 (
      {stage0_16[110]},
      {stage1_16[69]}
   );
   gpc1_1 gpc469 (
      {stage0_16[111]},
      {stage1_16[70]}
   );
   gpc1_1 gpc470 (
      {stage0_16[112]},
      {stage1_16[71]}
   );
   gpc1_1 gpc471 (
      {stage0_16[113]},
      {stage1_16[72]}
   );
   gpc1_1 gpc472 (
      {stage0_16[114]},
      {stage1_16[73]}
   );
   gpc1_1 gpc473 (
      {stage0_16[115]},
      {stage1_16[74]}
   );
   gpc1_1 gpc474 (
      {stage0_16[116]},
      {stage1_16[75]}
   );
   gpc1_1 gpc475 (
      {stage0_16[117]},
      {stage1_16[76]}
   );
   gpc1_1 gpc476 (
      {stage0_16[118]},
      {stage1_16[77]}
   );
   gpc1_1 gpc477 (
      {stage0_16[119]},
      {stage1_16[78]}
   );
   gpc1_1 gpc478 (
      {stage0_16[120]},
      {stage1_16[79]}
   );
   gpc1_1 gpc479 (
      {stage0_16[121]},
      {stage1_16[80]}
   );
   gpc1_1 gpc480 (
      {stage0_16[122]},
      {stage1_16[81]}
   );
   gpc1_1 gpc481 (
      {stage0_16[123]},
      {stage1_16[82]}
   );
   gpc1_1 gpc482 (
      {stage0_16[124]},
      {stage1_16[83]}
   );
   gpc1_1 gpc483 (
      {stage0_16[125]},
      {stage1_16[84]}
   );
   gpc1_1 gpc484 (
      {stage0_16[126]},
      {stage1_16[85]}
   );
   gpc1_1 gpc485 (
      {stage0_16[127]},
      {stage1_16[86]}
   );
   gpc1_1 gpc486 (
      {stage0_17[120]},
      {stage1_17[55]}
   );
   gpc1_1 gpc487 (
      {stage0_17[121]},
      {stage1_17[56]}
   );
   gpc1_1 gpc488 (
      {stage0_17[122]},
      {stage1_17[57]}
   );
   gpc1_1 gpc489 (
      {stage0_17[123]},
      {stage1_17[58]}
   );
   gpc1_1 gpc490 (
      {stage0_17[124]},
      {stage1_17[59]}
   );
   gpc1_1 gpc491 (
      {stage0_17[125]},
      {stage1_17[60]}
   );
   gpc1_1 gpc492 (
      {stage0_17[126]},
      {stage1_17[61]}
   );
   gpc1_1 gpc493 (
      {stage0_17[127]},
      {stage1_17[62]}
   );
   gpc1_1 gpc494 (
      {stage0_18[100]},
      {stage1_18[38]}
   );
   gpc1_1 gpc495 (
      {stage0_18[101]},
      {stage1_18[39]}
   );
   gpc1_1 gpc496 (
      {stage0_18[102]},
      {stage1_18[40]}
   );
   gpc1_1 gpc497 (
      {stage0_18[103]},
      {stage1_18[41]}
   );
   gpc1_1 gpc498 (
      {stage0_18[104]},
      {stage1_18[42]}
   );
   gpc1_1 gpc499 (
      {stage0_18[105]},
      {stage1_18[43]}
   );
   gpc1_1 gpc500 (
      {stage0_18[106]},
      {stage1_18[44]}
   );
   gpc1_1 gpc501 (
      {stage0_18[107]},
      {stage1_18[45]}
   );
   gpc1_1 gpc502 (
      {stage0_18[108]},
      {stage1_18[46]}
   );
   gpc1_1 gpc503 (
      {stage0_18[109]},
      {stage1_18[47]}
   );
   gpc1_1 gpc504 (
      {stage0_18[110]},
      {stage1_18[48]}
   );
   gpc1_1 gpc505 (
      {stage0_18[111]},
      {stage1_18[49]}
   );
   gpc1_1 gpc506 (
      {stage0_18[112]},
      {stage1_18[50]}
   );
   gpc1_1 gpc507 (
      {stage0_18[113]},
      {stage1_18[51]}
   );
   gpc1_1 gpc508 (
      {stage0_18[114]},
      {stage1_18[52]}
   );
   gpc1_1 gpc509 (
      {stage0_18[115]},
      {stage1_18[53]}
   );
   gpc1_1 gpc510 (
      {stage0_18[116]},
      {stage1_18[54]}
   );
   gpc1_1 gpc511 (
      {stage0_18[117]},
      {stage1_18[55]}
   );
   gpc1_1 gpc512 (
      {stage0_18[118]},
      {stage1_18[56]}
   );
   gpc1_1 gpc513 (
      {stage0_18[119]},
      {stage1_18[57]}
   );
   gpc1_1 gpc514 (
      {stage0_18[120]},
      {stage1_18[58]}
   );
   gpc1_1 gpc515 (
      {stage0_18[121]},
      {stage1_18[59]}
   );
   gpc1_1 gpc516 (
      {stage0_18[122]},
      {stage1_18[60]}
   );
   gpc1_1 gpc517 (
      {stage0_18[123]},
      {stage1_18[61]}
   );
   gpc1_1 gpc518 (
      {stage0_18[124]},
      {stage1_18[62]}
   );
   gpc1_1 gpc519 (
      {stage0_18[125]},
      {stage1_18[63]}
   );
   gpc1_1 gpc520 (
      {stage0_18[126]},
      {stage1_18[64]}
   );
   gpc1_1 gpc521 (
      {stage0_18[127]},
      {stage1_18[65]}
   );
   gpc1_1 gpc522 (
      {stage0_19[125]},
      {stage1_19[40]}
   );
   gpc1_1 gpc523 (
      {stage0_19[126]},
      {stage1_19[41]}
   );
   gpc1_1 gpc524 (
      {stage0_19[127]},
      {stage1_19[42]}
   );
   gpc1_1 gpc525 (
      {stage0_20[117]},
      {stage1_20[55]}
   );
   gpc1_1 gpc526 (
      {stage0_20[118]},
      {stage1_20[56]}
   );
   gpc1_1 gpc527 (
      {stage0_20[119]},
      {stage1_20[57]}
   );
   gpc1_1 gpc528 (
      {stage0_20[120]},
      {stage1_20[58]}
   );
   gpc1_1 gpc529 (
      {stage0_20[121]},
      {stage1_20[59]}
   );
   gpc1_1 gpc530 (
      {stage0_20[122]},
      {stage1_20[60]}
   );
   gpc1_1 gpc531 (
      {stage0_20[123]},
      {stage1_20[61]}
   );
   gpc1_1 gpc532 (
      {stage0_20[124]},
      {stage1_20[62]}
   );
   gpc1_1 gpc533 (
      {stage0_20[125]},
      {stage1_20[63]}
   );
   gpc1_1 gpc534 (
      {stage0_20[126]},
      {stage1_20[64]}
   );
   gpc1_1 gpc535 (
      {stage0_20[127]},
      {stage1_20[65]}
   );
   gpc1_1 gpc536 (
      {stage0_21[120]},
      {stage1_21[57]}
   );
   gpc1_1 gpc537 (
      {stage0_21[121]},
      {stage1_21[58]}
   );
   gpc1_1 gpc538 (
      {stage0_21[122]},
      {stage1_21[59]}
   );
   gpc1_1 gpc539 (
      {stage0_21[123]},
      {stage1_21[60]}
   );
   gpc1_1 gpc540 (
      {stage0_21[124]},
      {stage1_21[61]}
   );
   gpc1_1 gpc541 (
      {stage0_21[125]},
      {stage1_21[62]}
   );
   gpc1_1 gpc542 (
      {stage0_21[126]},
      {stage1_21[63]}
   );
   gpc1_1 gpc543 (
      {stage0_21[127]},
      {stage1_21[64]}
   );
   gpc1_1 gpc544 (
      {stage0_22[107]},
      {stage1_22[40]}
   );
   gpc1_1 gpc545 (
      {stage0_22[108]},
      {stage1_22[41]}
   );
   gpc1_1 gpc546 (
      {stage0_22[109]},
      {stage1_22[42]}
   );
   gpc1_1 gpc547 (
      {stage0_22[110]},
      {stage1_22[43]}
   );
   gpc1_1 gpc548 (
      {stage0_22[111]},
      {stage1_22[44]}
   );
   gpc1_1 gpc549 (
      {stage0_22[112]},
      {stage1_22[45]}
   );
   gpc1_1 gpc550 (
      {stage0_22[113]},
      {stage1_22[46]}
   );
   gpc1_1 gpc551 (
      {stage0_22[114]},
      {stage1_22[47]}
   );
   gpc1_1 gpc552 (
      {stage0_22[115]},
      {stage1_22[48]}
   );
   gpc1_1 gpc553 (
      {stage0_22[116]},
      {stage1_22[49]}
   );
   gpc1_1 gpc554 (
      {stage0_22[117]},
      {stage1_22[50]}
   );
   gpc1_1 gpc555 (
      {stage0_22[118]},
      {stage1_22[51]}
   );
   gpc1_1 gpc556 (
      {stage0_22[119]},
      {stage1_22[52]}
   );
   gpc1_1 gpc557 (
      {stage0_22[120]},
      {stage1_22[53]}
   );
   gpc1_1 gpc558 (
      {stage0_22[121]},
      {stage1_22[54]}
   );
   gpc1_1 gpc559 (
      {stage0_22[122]},
      {stage1_22[55]}
   );
   gpc1_1 gpc560 (
      {stage0_22[123]},
      {stage1_22[56]}
   );
   gpc1_1 gpc561 (
      {stage0_22[124]},
      {stage1_22[57]}
   );
   gpc1_1 gpc562 (
      {stage0_22[125]},
      {stage1_22[58]}
   );
   gpc1_1 gpc563 (
      {stage0_22[126]},
      {stage1_22[59]}
   );
   gpc1_1 gpc564 (
      {stage0_22[127]},
      {stage1_22[60]}
   );
   gpc1_1 gpc565 (
      {stage0_23[126]},
      {stage1_23[42]}
   );
   gpc1_1 gpc566 (
      {stage0_23[127]},
      {stage1_23[43]}
   );
   gpc1_1 gpc567 (
      {stage0_24[91]},
      {stage1_24[53]}
   );
   gpc1_1 gpc568 (
      {stage0_24[92]},
      {stage1_24[54]}
   );
   gpc1_1 gpc569 (
      {stage0_24[93]},
      {stage1_24[55]}
   );
   gpc1_1 gpc570 (
      {stage0_24[94]},
      {stage1_24[56]}
   );
   gpc1_1 gpc571 (
      {stage0_24[95]},
      {stage1_24[57]}
   );
   gpc1_1 gpc572 (
      {stage0_24[96]},
      {stage1_24[58]}
   );
   gpc1_1 gpc573 (
      {stage0_24[97]},
      {stage1_24[59]}
   );
   gpc1_1 gpc574 (
      {stage0_24[98]},
      {stage1_24[60]}
   );
   gpc1_1 gpc575 (
      {stage0_24[99]},
      {stage1_24[61]}
   );
   gpc1_1 gpc576 (
      {stage0_24[100]},
      {stage1_24[62]}
   );
   gpc1_1 gpc577 (
      {stage0_24[101]},
      {stage1_24[63]}
   );
   gpc1_1 gpc578 (
      {stage0_24[102]},
      {stage1_24[64]}
   );
   gpc1_1 gpc579 (
      {stage0_24[103]},
      {stage1_24[65]}
   );
   gpc1_1 gpc580 (
      {stage0_24[104]},
      {stage1_24[66]}
   );
   gpc1_1 gpc581 (
      {stage0_24[105]},
      {stage1_24[67]}
   );
   gpc1_1 gpc582 (
      {stage0_24[106]},
      {stage1_24[68]}
   );
   gpc1_1 gpc583 (
      {stage0_24[107]},
      {stage1_24[69]}
   );
   gpc1_1 gpc584 (
      {stage0_24[108]},
      {stage1_24[70]}
   );
   gpc1_1 gpc585 (
      {stage0_24[109]},
      {stage1_24[71]}
   );
   gpc1_1 gpc586 (
      {stage0_24[110]},
      {stage1_24[72]}
   );
   gpc1_1 gpc587 (
      {stage0_24[111]},
      {stage1_24[73]}
   );
   gpc1_1 gpc588 (
      {stage0_24[112]},
      {stage1_24[74]}
   );
   gpc1_1 gpc589 (
      {stage0_24[113]},
      {stage1_24[75]}
   );
   gpc1_1 gpc590 (
      {stage0_24[114]},
      {stage1_24[76]}
   );
   gpc1_1 gpc591 (
      {stage0_24[115]},
      {stage1_24[77]}
   );
   gpc1_1 gpc592 (
      {stage0_24[116]},
      {stage1_24[78]}
   );
   gpc1_1 gpc593 (
      {stage0_24[117]},
      {stage1_24[79]}
   );
   gpc1_1 gpc594 (
      {stage0_24[118]},
      {stage1_24[80]}
   );
   gpc1_1 gpc595 (
      {stage0_24[119]},
      {stage1_24[81]}
   );
   gpc1_1 gpc596 (
      {stage0_24[120]},
      {stage1_24[82]}
   );
   gpc1_1 gpc597 (
      {stage0_24[121]},
      {stage1_24[83]}
   );
   gpc1_1 gpc598 (
      {stage0_24[122]},
      {stage1_24[84]}
   );
   gpc1_1 gpc599 (
      {stage0_24[123]},
      {stage1_24[85]}
   );
   gpc1_1 gpc600 (
      {stage0_24[124]},
      {stage1_24[86]}
   );
   gpc1_1 gpc601 (
      {stage0_24[125]},
      {stage1_24[87]}
   );
   gpc1_1 gpc602 (
      {stage0_24[126]},
      {stage1_24[88]}
   );
   gpc1_1 gpc603 (
      {stage0_24[127]},
      {stage1_24[89]}
   );
   gpc1_1 gpc604 (
      {stage0_25[108]},
      {stage1_25[50]}
   );
   gpc1_1 gpc605 (
      {stage0_25[109]},
      {stage1_25[51]}
   );
   gpc1_1 gpc606 (
      {stage0_25[110]},
      {stage1_25[52]}
   );
   gpc1_1 gpc607 (
      {stage0_25[111]},
      {stage1_25[53]}
   );
   gpc1_1 gpc608 (
      {stage0_25[112]},
      {stage1_25[54]}
   );
   gpc1_1 gpc609 (
      {stage0_25[113]},
      {stage1_25[55]}
   );
   gpc1_1 gpc610 (
      {stage0_25[114]},
      {stage1_25[56]}
   );
   gpc1_1 gpc611 (
      {stage0_25[115]},
      {stage1_25[57]}
   );
   gpc1_1 gpc612 (
      {stage0_25[116]},
      {stage1_25[58]}
   );
   gpc1_1 gpc613 (
      {stage0_25[117]},
      {stage1_25[59]}
   );
   gpc1_1 gpc614 (
      {stage0_25[118]},
      {stage1_25[60]}
   );
   gpc1_1 gpc615 (
      {stage0_25[119]},
      {stage1_25[61]}
   );
   gpc1_1 gpc616 (
      {stage0_25[120]},
      {stage1_25[62]}
   );
   gpc1_1 gpc617 (
      {stage0_25[121]},
      {stage1_25[63]}
   );
   gpc1_1 gpc618 (
      {stage0_25[122]},
      {stage1_25[64]}
   );
   gpc1_1 gpc619 (
      {stage0_25[123]},
      {stage1_25[65]}
   );
   gpc1_1 gpc620 (
      {stage0_25[124]},
      {stage1_25[66]}
   );
   gpc1_1 gpc621 (
      {stage0_25[125]},
      {stage1_25[67]}
   );
   gpc1_1 gpc622 (
      {stage0_25[126]},
      {stage1_25[68]}
   );
   gpc1_1 gpc623 (
      {stage0_25[127]},
      {stage1_25[69]}
   );
   gpc1_1 gpc624 (
      {stage0_26[94]},
      {stage1_26[35]}
   );
   gpc1_1 gpc625 (
      {stage0_26[95]},
      {stage1_26[36]}
   );
   gpc1_1 gpc626 (
      {stage0_26[96]},
      {stage1_26[37]}
   );
   gpc1_1 gpc627 (
      {stage0_26[97]},
      {stage1_26[38]}
   );
   gpc1_1 gpc628 (
      {stage0_26[98]},
      {stage1_26[39]}
   );
   gpc1_1 gpc629 (
      {stage0_26[99]},
      {stage1_26[40]}
   );
   gpc1_1 gpc630 (
      {stage0_26[100]},
      {stage1_26[41]}
   );
   gpc1_1 gpc631 (
      {stage0_26[101]},
      {stage1_26[42]}
   );
   gpc1_1 gpc632 (
      {stage0_26[102]},
      {stage1_26[43]}
   );
   gpc1_1 gpc633 (
      {stage0_26[103]},
      {stage1_26[44]}
   );
   gpc1_1 gpc634 (
      {stage0_26[104]},
      {stage1_26[45]}
   );
   gpc1_1 gpc635 (
      {stage0_26[105]},
      {stage1_26[46]}
   );
   gpc1_1 gpc636 (
      {stage0_26[106]},
      {stage1_26[47]}
   );
   gpc1_1 gpc637 (
      {stage0_26[107]},
      {stage1_26[48]}
   );
   gpc1_1 gpc638 (
      {stage0_26[108]},
      {stage1_26[49]}
   );
   gpc1_1 gpc639 (
      {stage0_26[109]},
      {stage1_26[50]}
   );
   gpc1_1 gpc640 (
      {stage0_26[110]},
      {stage1_26[51]}
   );
   gpc1_1 gpc641 (
      {stage0_26[111]},
      {stage1_26[52]}
   );
   gpc1_1 gpc642 (
      {stage0_26[112]},
      {stage1_26[53]}
   );
   gpc1_1 gpc643 (
      {stage0_26[113]},
      {stage1_26[54]}
   );
   gpc1_1 gpc644 (
      {stage0_26[114]},
      {stage1_26[55]}
   );
   gpc1_1 gpc645 (
      {stage0_26[115]},
      {stage1_26[56]}
   );
   gpc1_1 gpc646 (
      {stage0_26[116]},
      {stage1_26[57]}
   );
   gpc1_1 gpc647 (
      {stage0_26[117]},
      {stage1_26[58]}
   );
   gpc1_1 gpc648 (
      {stage0_26[118]},
      {stage1_26[59]}
   );
   gpc1_1 gpc649 (
      {stage0_26[119]},
      {stage1_26[60]}
   );
   gpc1_1 gpc650 (
      {stage0_26[120]},
      {stage1_26[61]}
   );
   gpc1_1 gpc651 (
      {stage0_26[121]},
      {stage1_26[62]}
   );
   gpc1_1 gpc652 (
      {stage0_26[122]},
      {stage1_26[63]}
   );
   gpc1_1 gpc653 (
      {stage0_26[123]},
      {stage1_26[64]}
   );
   gpc1_1 gpc654 (
      {stage0_26[124]},
      {stage1_26[65]}
   );
   gpc1_1 gpc655 (
      {stage0_26[125]},
      {stage1_26[66]}
   );
   gpc1_1 gpc656 (
      {stage0_26[126]},
      {stage1_26[67]}
   );
   gpc1_1 gpc657 (
      {stage0_26[127]},
      {stage1_26[68]}
   );
   gpc1_1 gpc658 (
      {stage0_27[111]},
      {stage1_27[39]}
   );
   gpc1_1 gpc659 (
      {stage0_27[112]},
      {stage1_27[40]}
   );
   gpc1_1 gpc660 (
      {stage0_27[113]},
      {stage1_27[41]}
   );
   gpc1_1 gpc661 (
      {stage0_27[114]},
      {stage1_27[42]}
   );
   gpc1_1 gpc662 (
      {stage0_27[115]},
      {stage1_27[43]}
   );
   gpc1_1 gpc663 (
      {stage0_27[116]},
      {stage1_27[44]}
   );
   gpc1_1 gpc664 (
      {stage0_27[117]},
      {stage1_27[45]}
   );
   gpc1_1 gpc665 (
      {stage0_27[118]},
      {stage1_27[46]}
   );
   gpc1_1 gpc666 (
      {stage0_27[119]},
      {stage1_27[47]}
   );
   gpc1_1 gpc667 (
      {stage0_27[120]},
      {stage1_27[48]}
   );
   gpc1_1 gpc668 (
      {stage0_27[121]},
      {stage1_27[49]}
   );
   gpc1_1 gpc669 (
      {stage0_27[122]},
      {stage1_27[50]}
   );
   gpc1_1 gpc670 (
      {stage0_27[123]},
      {stage1_27[51]}
   );
   gpc1_1 gpc671 (
      {stage0_27[124]},
      {stage1_27[52]}
   );
   gpc1_1 gpc672 (
      {stage0_27[125]},
      {stage1_27[53]}
   );
   gpc1_1 gpc673 (
      {stage0_27[126]},
      {stage1_27[54]}
   );
   gpc1_1 gpc674 (
      {stage0_27[127]},
      {stage1_27[55]}
   );
   gpc1_1 gpc675 (
      {stage0_28[125]},
      {stage1_28[53]}
   );
   gpc1_1 gpc676 (
      {stage0_28[126]},
      {stage1_28[54]}
   );
   gpc1_1 gpc677 (
      {stage0_28[127]},
      {stage1_28[55]}
   );
   gpc1_1 gpc678 (
      {stage0_29[126]},
      {stage1_29[55]}
   );
   gpc1_1 gpc679 (
      {stage0_29[127]},
      {stage1_29[56]}
   );
   gpc1_1 gpc680 (
      {stage0_30[108]},
      {stage1_30[41]}
   );
   gpc1_1 gpc681 (
      {stage0_30[109]},
      {stage1_30[42]}
   );
   gpc1_1 gpc682 (
      {stage0_30[110]},
      {stage1_30[43]}
   );
   gpc1_1 gpc683 (
      {stage0_30[111]},
      {stage1_30[44]}
   );
   gpc1_1 gpc684 (
      {stage0_30[112]},
      {stage1_30[45]}
   );
   gpc1_1 gpc685 (
      {stage0_30[113]},
      {stage1_30[46]}
   );
   gpc1_1 gpc686 (
      {stage0_30[114]},
      {stage1_30[47]}
   );
   gpc1_1 gpc687 (
      {stage0_30[115]},
      {stage1_30[48]}
   );
   gpc1_1 gpc688 (
      {stage0_30[116]},
      {stage1_30[49]}
   );
   gpc1_1 gpc689 (
      {stage0_30[117]},
      {stage1_30[50]}
   );
   gpc1_1 gpc690 (
      {stage0_30[118]},
      {stage1_30[51]}
   );
   gpc1_1 gpc691 (
      {stage0_30[119]},
      {stage1_30[52]}
   );
   gpc1_1 gpc692 (
      {stage0_30[120]},
      {stage1_30[53]}
   );
   gpc1_1 gpc693 (
      {stage0_30[121]},
      {stage1_30[54]}
   );
   gpc1_1 gpc694 (
      {stage0_30[122]},
      {stage1_30[55]}
   );
   gpc1_1 gpc695 (
      {stage0_30[123]},
      {stage1_30[56]}
   );
   gpc1_1 gpc696 (
      {stage0_30[124]},
      {stage1_30[57]}
   );
   gpc1_1 gpc697 (
      {stage0_30[125]},
      {stage1_30[58]}
   );
   gpc1_1 gpc698 (
      {stage0_30[126]},
      {stage1_30[59]}
   );
   gpc1_1 gpc699 (
      {stage0_30[127]},
      {stage1_30[60]}
   );
   gpc1_1 gpc700 (
      {stage0_31[96]},
      {stage1_31[39]}
   );
   gpc1_1 gpc701 (
      {stage0_31[97]},
      {stage1_31[40]}
   );
   gpc1_1 gpc702 (
      {stage0_31[98]},
      {stage1_31[41]}
   );
   gpc1_1 gpc703 (
      {stage0_31[99]},
      {stage1_31[42]}
   );
   gpc1_1 gpc704 (
      {stage0_31[100]},
      {stage1_31[43]}
   );
   gpc1_1 gpc705 (
      {stage0_31[101]},
      {stage1_31[44]}
   );
   gpc1_1 gpc706 (
      {stage0_31[102]},
      {stage1_31[45]}
   );
   gpc1_1 gpc707 (
      {stage0_31[103]},
      {stage1_31[46]}
   );
   gpc1_1 gpc708 (
      {stage0_31[104]},
      {stage1_31[47]}
   );
   gpc1_1 gpc709 (
      {stage0_31[105]},
      {stage1_31[48]}
   );
   gpc1_1 gpc710 (
      {stage0_31[106]},
      {stage1_31[49]}
   );
   gpc1_1 gpc711 (
      {stage0_31[107]},
      {stage1_31[50]}
   );
   gpc1_1 gpc712 (
      {stage0_31[108]},
      {stage1_31[51]}
   );
   gpc1_1 gpc713 (
      {stage0_31[109]},
      {stage1_31[52]}
   );
   gpc1_1 gpc714 (
      {stage0_31[110]},
      {stage1_31[53]}
   );
   gpc1_1 gpc715 (
      {stage0_31[111]},
      {stage1_31[54]}
   );
   gpc1_1 gpc716 (
      {stage0_31[112]},
      {stage1_31[55]}
   );
   gpc1_1 gpc717 (
      {stage0_31[113]},
      {stage1_31[56]}
   );
   gpc1_1 gpc718 (
      {stage0_31[114]},
      {stage1_31[57]}
   );
   gpc1_1 gpc719 (
      {stage0_31[115]},
      {stage1_31[58]}
   );
   gpc1_1 gpc720 (
      {stage0_31[116]},
      {stage1_31[59]}
   );
   gpc1_1 gpc721 (
      {stage0_31[117]},
      {stage1_31[60]}
   );
   gpc1_1 gpc722 (
      {stage0_31[118]},
      {stage1_31[61]}
   );
   gpc1_1 gpc723 (
      {stage0_31[119]},
      {stage1_31[62]}
   );
   gpc1_1 gpc724 (
      {stage0_31[120]},
      {stage1_31[63]}
   );
   gpc1_1 gpc725 (
      {stage0_31[121]},
      {stage1_31[64]}
   );
   gpc1_1 gpc726 (
      {stage0_31[122]},
      {stage1_31[65]}
   );
   gpc1_1 gpc727 (
      {stage0_31[123]},
      {stage1_31[66]}
   );
   gpc1_1 gpc728 (
      {stage0_31[124]},
      {stage1_31[67]}
   );
   gpc1_1 gpc729 (
      {stage0_31[125]},
      {stage1_31[68]}
   );
   gpc1_1 gpc730 (
      {stage0_31[126]},
      {stage1_31[69]}
   );
   gpc1_1 gpc731 (
      {stage0_31[127]},
      {stage1_31[70]}
   );
   gpc606_5 gpc732 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0]}
   );
   gpc606_5 gpc733 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc734 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc735 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc736 (
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc737 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc606_5 gpc738 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc739 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[24]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc740 (
      {stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage1_3[25]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc741 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32]},
      {stage1_3[26]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc742 (
      {stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37]},
      {stage1_3[27]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc743 (
      {stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage1_3[28]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[11],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc744 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[12],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc745 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[13],stage2_4[13],stage2_3[13]}
   );
   gpc606_5 gpc746 (
      {stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[2],stage2_6[10],stage2_5[14],stage2_4[14]}
   );
   gpc606_5 gpc747 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[11],stage2_5[15]}
   );
   gpc606_5 gpc748 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[12],stage2_5[16]}
   );
   gpc606_5 gpc749 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[13],stage2_5[17]}
   );
   gpc606_5 gpc750 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[14],stage2_5[18]}
   );
   gpc606_5 gpc751 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[15],stage2_5[19]}
   );
   gpc606_5 gpc752 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[6],stage2_7[8],stage2_6[16],stage2_5[20]}
   );
   gpc606_5 gpc753 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[7],stage2_7[9],stage2_6[17],stage2_5[21]}
   );
   gpc606_5 gpc754 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[7],stage2_8[8],stage2_7[10],stage2_6[18]}
   );
   gpc606_5 gpc755 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[8],stage2_8[9],stage2_7[11],stage2_6[19]}
   );
   gpc615_5 gpc756 (
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22]},
      {stage1_7[42]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[9],stage2_8[10],stage2_7[12],stage2_6[20]}
   );
   gpc615_5 gpc757 (
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[10],stage2_8[11],stage2_7[13]}
   );
   gpc615_5 gpc758 (
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[11],stage2_8[12],stage2_7[14]}
   );
   gpc615_5 gpc759 (
      {stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[12],stage2_8[13],stage2_7[15]}
   );
   gpc615_5 gpc760 (
      {stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[13],stage2_8[14],stage2_7[16]}
   );
   gpc615_5 gpc761 (
      {stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66], stage1_7[67]},
      {stage1_8[22]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[7],stage2_9[14],stage2_8[15],stage2_7[17]}
   );
   gpc606_5 gpc762 (
      {stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[5],stage2_10[8],stage2_9[15],stage2_8[16]}
   );
   gpc606_5 gpc763 (
      {stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[6],stage2_10[9],stage2_9[16],stage2_8[17]}
   );
   gpc606_5 gpc764 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[7],stage2_10[10],stage2_9[17]}
   );
   gpc606_5 gpc765 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[8],stage2_10[11],stage2_9[18]}
   );
   gpc606_5 gpc766 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[4],stage2_11[9],stage2_10[12],stage2_9[19]}
   );
   gpc606_5 gpc767 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[5],stage2_11[10],stage2_10[13],stage2_9[20]}
   );
   gpc606_5 gpc768 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[6],stage2_11[11],stage2_10[14],stage2_9[21]}
   );
   gpc606_5 gpc769 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[5],stage2_12[7],stage2_11[12],stage2_10[15]}
   );
   gpc606_5 gpc770 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[6],stage2_12[8],stage2_11[13],stage2_10[16]}
   );
   gpc606_5 gpc771 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[7],stage2_12[9],stage2_11[14],stage2_10[17]}
   );
   gpc606_5 gpc772 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[8],stage2_12[10],stage2_11[15],stage2_10[18]}
   );
   gpc606_5 gpc773 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[9],stage2_12[11],stage2_11[16],stage2_10[19]}
   );
   gpc606_5 gpc774 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[10],stage2_12[12],stage2_11[17],stage2_10[20]}
   );
   gpc606_5 gpc775 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[11],stage2_12[13],stage2_11[18],stage2_10[21]}
   );
   gpc615_5 gpc776 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[42]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[12],stage2_12[14],stage2_11[19]}
   );
   gpc615_5 gpc777 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[43]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[13],stage2_12[15],stage2_11[20]}
   );
   gpc615_5 gpc778 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], stage1_11[44]},
      {stage1_12[44]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[14],stage2_12[16],stage2_11[21]}
   );
   gpc615_5 gpc779 (
      {stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48], stage1_11[49]},
      {stage1_12[45]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[15],stage2_12[17],stage2_11[22]}
   );
   gpc615_5 gpc780 (
      {stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage1_12[46]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[16],stage2_12[18],stage2_11[23]}
   );
   gpc606_5 gpc781 (
      {stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[5],stage2_14[12],stage2_13[17],stage2_12[19]}
   );
   gpc606_5 gpc782 (
      {stage1_12[53], stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], 1'b0},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[6],stage2_14[13],stage2_13[18],stage2_12[20]}
   );
   gpc606_5 gpc783 (
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[2],stage2_15[7],stage2_14[14],stage2_13[19]}
   );
   gpc606_5 gpc784 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[3],stage2_15[8],stage2_14[15],stage2_13[20]}
   );
   gpc606_5 gpc785 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[4],stage2_15[9],stage2_14[16],stage2_13[21]}
   );
   gpc615_5 gpc786 (
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16]},
      {stage1_15[18]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[3],stage2_16[5],stage2_15[10],stage2_14[17]}
   );
   gpc615_5 gpc787 (
      {stage1_14[17], stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21]},
      {stage1_15[19]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[4],stage2_16[6],stage2_15[11],stage2_14[18]}
   );
   gpc615_5 gpc788 (
      {stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26]},
      {stage1_15[20]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[5],stage2_16[7],stage2_15[12],stage2_14[19]}
   );
   gpc615_5 gpc789 (
      {stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage1_15[21]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[6],stage2_16[8],stage2_15[13],stage2_14[20]}
   );
   gpc615_5 gpc790 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_15[22]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[7],stage2_16[9],stage2_15[14],stage2_14[21]}
   );
   gpc615_5 gpc791 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_15[23]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[8],stage2_16[10],stage2_15[15],stage2_14[22]}
   );
   gpc615_5 gpc792 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28]},
      {stage1_16[36]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[6],stage2_17[9],stage2_16[11],stage2_15[16]}
   );
   gpc615_5 gpc793 (
      {stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage1_16[37]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[7],stage2_17[10],stage2_16[12],stage2_15[17]}
   );
   gpc615_5 gpc794 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38]},
      {stage1_16[38]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[8],stage2_17[11],stage2_16[13],stage2_15[18]}
   );
   gpc615_5 gpc795 (
      {stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_16[39]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[9],stage2_17[12],stage2_16[14],stage2_15[19]}
   );
   gpc606_5 gpc796 (
      {stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[4],stage2_18[10],stage2_17[13],stage2_16[15]}
   );
   gpc606_5 gpc797 (
      {stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[5],stage2_18[11],stage2_17[14],stage2_16[16]}
   );
   gpc606_5 gpc798 (
      {stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[6],stage2_18[12],stage2_17[15],stage2_16[17]}
   );
   gpc606_5 gpc799 (
      {stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[7],stage2_18[13],stage2_17[16],stage2_16[18]}
   );
   gpc606_5 gpc800 (
      {stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[8],stage2_18[14],stage2_17[17],stage2_16[19]}
   );
   gpc606_5 gpc801 (
      {stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[9],stage2_18[15],stage2_17[18],stage2_16[20]}
   );
   gpc606_5 gpc802 (
      {stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[10],stage2_18[16],stage2_17[19],stage2_16[21]}
   );
   gpc615_5 gpc803 (
      {stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86]},
      {stage1_17[24]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[11],stage2_18[17],stage2_17[20],stage2_16[22]}
   );
   gpc606_5 gpc804 (
      {stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[8],stage2_19[12],stage2_18[18],stage2_17[21]}
   );
   gpc606_5 gpc805 (
      {stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[9],stage2_19[13],stage2_18[19],stage2_17[22]}
   );
   gpc615_5 gpc806 (
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[2],stage2_20[10],stage2_19[14]}
   );
   gpc615_5 gpc807 (
      {stage1_19[17], stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[3],stage2_20[11],stage2_19[15]}
   );
   gpc615_5 gpc808 (
      {stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25], stage1_19[26]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[4],stage2_20[12],stage2_19[16]}
   );
   gpc615_5 gpc809 (
      {stage1_19[27], stage1_19[28], stage1_19[29], stage1_19[30], stage1_19[31]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[5],stage2_20[13],stage2_19[17]}
   );
   gpc615_5 gpc810 (
      {stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35], stage1_19[36]},
      {stage1_20[4]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[6],stage2_20[14],stage2_19[18]}
   );
   gpc615_5 gpc811 (
      {stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage1_20[5]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[7],stage2_20[15],stage2_19[19]}
   );
   gpc606_5 gpc812 (
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[6],stage2_22[6],stage2_21[8],stage2_20[16]}
   );
   gpc606_5 gpc813 (
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[7],stage2_22[7],stage2_21[9],stage2_20[17]}
   );
   gpc606_5 gpc814 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[8],stage2_22[8],stage2_21[10],stage2_20[18]}
   );
   gpc606_5 gpc815 (
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[9],stage2_22[9],stage2_21[11],stage2_20[19]}
   );
   gpc606_5 gpc816 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[4],stage2_23[10],stage2_22[10],stage2_21[12]}
   );
   gpc606_5 gpc817 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[5],stage2_23[11],stage2_22[11],stage2_21[13]}
   );
   gpc606_5 gpc818 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[6],stage2_23[12],stage2_22[12],stage2_21[14]}
   );
   gpc606_5 gpc819 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[7],stage2_23[13],stage2_22[13],stage2_21[15]}
   );
   gpc606_5 gpc820 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[8],stage2_23[14],stage2_22[14]}
   );
   gpc606_5 gpc821 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[9],stage2_23[15],stage2_22[15]}
   );
   gpc606_5 gpc822 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[10],stage2_23[16],stage2_22[16]}
   );
   gpc606_5 gpc823 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[11],stage2_23[17],stage2_22[17]}
   );
   gpc615_5 gpc824 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52]},
      {stage1_23[24]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[12],stage2_23[18],stage2_22[18]}
   );
   gpc615_5 gpc825 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage1_24[30]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[5],stage2_25[9],stage2_24[13],stage2_23[19]}
   );
   gpc606_5 gpc826 (
      {stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[6],stage2_25[10],stage2_24[14]}
   );
   gpc606_5 gpc827 (
      {stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[7],stage2_25[11],stage2_24[15]}
   );
   gpc606_5 gpc828 (
      {stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[3],stage2_26[8],stage2_25[12],stage2_24[16]}
   );
   gpc606_5 gpc829 (
      {stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[4],stage2_26[9],stage2_25[13],stage2_24[17]}
   );
   gpc606_5 gpc830 (
      {stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59], stage1_24[60]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[5],stage2_26[10],stage2_25[14],stage2_24[18]}
   );
   gpc606_5 gpc831 (
      {stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65], stage1_24[66]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[6],stage2_26[11],stage2_25[15],stage2_24[19]}
   );
   gpc606_5 gpc832 (
      {stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71], stage1_24[72]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[7],stage2_26[12],stage2_25[16],stage2_24[20]}
   );
   gpc606_5 gpc833 (
      {stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77], stage1_24[78]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[8],stage2_26[13],stage2_25[17],stage2_24[21]}
   );
   gpc606_5 gpc834 (
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[8],stage2_27[9],stage2_26[14],stage2_25[18]}
   );
   gpc606_5 gpc835 (
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[9],stage2_27[10],stage2_26[15],stage2_25[19]}
   );
   gpc606_5 gpc836 (
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[10],stage2_27[11],stage2_26[16],stage2_25[20]}
   );
   gpc606_5 gpc837 (
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[11],stage2_27[12],stage2_26[17],stage2_25[21]}
   );
   gpc606_5 gpc838 (
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[12],stage2_27[13],stage2_26[18],stage2_25[22]}
   );
   gpc606_5 gpc839 (
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[13],stage2_27[14],stage2_26[19],stage2_25[23]}
   );
   gpc606_5 gpc840 (
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[14],stage2_27[15],stage2_26[20],stage2_25[24]}
   );
   gpc606_5 gpc841 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[7],stage2_28[15],stage2_27[16],stage2_26[21]}
   );
   gpc606_5 gpc842 (
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[0],stage2_30[1],stage2_29[8],stage2_28[16]}
   );
   gpc606_5 gpc843 (
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[1],stage2_30[2],stage2_29[9],stage2_28[17]}
   );
   gpc606_5 gpc844 (
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[2],stage2_30[3],stage2_29[10],stage2_28[18]}
   );
   gpc606_5 gpc845 (
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[3],stage2_30[4],stage2_29[11],stage2_28[19]}
   );
   gpc606_5 gpc846 (
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[4],stage2_30[5],stage2_29[12],stage2_28[20]}
   );
   gpc606_5 gpc847 (
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[5],stage2_30[6],stage2_29[13],stage2_28[21]}
   );
   gpc606_5 gpc848 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[6],stage2_31[6],stage2_30[7],stage2_29[14]}
   );
   gpc606_5 gpc849 (
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[7],stage2_31[7],stage2_30[8],stage2_29[15]}
   );
   gpc606_5 gpc850 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[8],stage2_31[8],stage2_30[9],stage2_29[16]}
   );
   gpc606_5 gpc851 (
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[9],stage2_31[9],stage2_30[10],stage2_29[17]}
   );
   gpc606_5 gpc852 (
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[10],stage2_31[10],stage2_30[11],stage2_29[18]}
   );
   gpc606_5 gpc853 (
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[11],stage2_31[11],stage2_30[12],stage2_29[19]}
   );
   gpc606_5 gpc854 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[12],stage2_31[12],stage2_30[13],stage2_29[20]}
   );
   gpc1325_5 gpc855 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46]},
      {stage1_30[36], stage1_30[37]},
      {stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_32[0]},
      {stage2_33[7],stage2_32[13],stage2_31[13],stage2_30[14],stage2_29[21]}
   );
   gpc606_5 gpc856 (
      {stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41], stage1_30[42], stage1_30[43]},
      {stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6]},
      {stage2_34[0],stage2_33[8],stage2_32[14],stage2_31[14],stage2_30[15]}
   );
   gpc606_5 gpc857 (
      {stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47], stage1_30[48], stage1_30[49]},
      {stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12]},
      {stage2_34[1],stage2_33[9],stage2_32[15],stage2_31[15],stage2_30[16]}
   );
   gpc606_5 gpc858 (
      {stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54], stage1_30[55]},
      {stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17], stage1_32[18]},
      {stage2_34[2],stage2_33[10],stage2_32[16],stage2_31[16],stage2_30[17]}
   );
   gpc606_5 gpc859 (
      {stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], 1'b0},
      {stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23], stage1_32[24]},
      {stage2_34[3],stage2_33[11],stage2_32[17],stage2_31[17],stage2_30[18]}
   );
   gpc606_5 gpc860 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[4],stage2_33[12],stage2_32[18],stage2_31[18]}
   );
   gpc606_5 gpc861 (
      {stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54], stage1_31[55], stage1_31[56]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[5],stage2_33[13],stage2_32[19],stage2_31[19]}
   );
   gpc1_1 gpc862 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc863 (
      {stage1_0[1]},
      {stage2_0[1]}
   );
   gpc1_1 gpc864 (
      {stage1_0[2]},
      {stage2_0[2]}
   );
   gpc1_1 gpc865 (
      {stage1_0[3]},
      {stage2_0[3]}
   );
   gpc1_1 gpc866 (
      {stage1_0[4]},
      {stage2_0[4]}
   );
   gpc1_1 gpc867 (
      {stage1_0[5]},
      {stage2_0[5]}
   );
   gpc1_1 gpc868 (
      {stage1_0[6]},
      {stage2_0[6]}
   );
   gpc1_1 gpc869 (
      {stage1_0[7]},
      {stage2_0[7]}
   );
   gpc1_1 gpc870 (
      {stage1_0[8]},
      {stage2_0[8]}
   );
   gpc1_1 gpc871 (
      {stage1_0[9]},
      {stage2_0[9]}
   );
   gpc1_1 gpc872 (
      {stage1_0[10]},
      {stage2_0[10]}
   );
   gpc1_1 gpc873 (
      {stage1_0[11]},
      {stage2_0[11]}
   );
   gpc1_1 gpc874 (
      {stage1_0[12]},
      {stage2_0[12]}
   );
   gpc1_1 gpc875 (
      {stage1_0[13]},
      {stage2_0[13]}
   );
   gpc1_1 gpc876 (
      {stage1_0[14]},
      {stage2_0[14]}
   );
   gpc1_1 gpc877 (
      {stage1_0[15]},
      {stage2_0[15]}
   );
   gpc1_1 gpc878 (
      {stage1_0[16]},
      {stage2_0[16]}
   );
   gpc1_1 gpc879 (
      {stage1_0[17]},
      {stage2_0[17]}
   );
   gpc1_1 gpc880 (
      {stage1_0[18]},
      {stage2_0[18]}
   );
   gpc1_1 gpc881 (
      {stage1_0[19]},
      {stage2_0[19]}
   );
   gpc1_1 gpc882 (
      {stage1_0[20]},
      {stage2_0[20]}
   );
   gpc1_1 gpc883 (
      {stage1_0[21]},
      {stage2_0[21]}
   );
   gpc1_1 gpc884 (
      {stage1_0[22]},
      {stage2_0[22]}
   );
   gpc1_1 gpc885 (
      {stage1_0[23]},
      {stage2_0[23]}
   );
   gpc1_1 gpc886 (
      {stage1_0[24]},
      {stage2_0[24]}
   );
   gpc1_1 gpc887 (
      {stage1_0[25]},
      {stage2_0[25]}
   );
   gpc1_1 gpc888 (
      {stage1_0[26]},
      {stage2_0[26]}
   );
   gpc1_1 gpc889 (
      {stage1_0[27]},
      {stage2_0[27]}
   );
   gpc1_1 gpc890 (
      {stage1_0[28]},
      {stage2_0[28]}
   );
   gpc1_1 gpc891 (
      {stage1_0[29]},
      {stage2_0[29]}
   );
   gpc1_1 gpc892 (
      {stage1_0[30]},
      {stage2_0[30]}
   );
   gpc1_1 gpc893 (
      {stage1_0[31]},
      {stage2_0[31]}
   );
   gpc1_1 gpc894 (
      {stage1_0[32]},
      {stage2_0[32]}
   );
   gpc1_1 gpc895 (
      {stage1_0[33]},
      {stage2_0[33]}
   );
   gpc1_1 gpc896 (
      {stage1_0[34]},
      {stage2_0[34]}
   );
   gpc1_1 gpc897 (
      {stage1_0[35]},
      {stage2_0[35]}
   );
   gpc1_1 gpc898 (
      {stage1_1[24]},
      {stage2_1[4]}
   );
   gpc1_1 gpc899 (
      {stage1_1[25]},
      {stage2_1[5]}
   );
   gpc1_1 gpc900 (
      {stage1_1[26]},
      {stage2_1[6]}
   );
   gpc1_1 gpc901 (
      {stage1_1[27]},
      {stage2_1[7]}
   );
   gpc1_1 gpc902 (
      {stage1_1[28]},
      {stage2_1[8]}
   );
   gpc1_1 gpc903 (
      {stage1_1[29]},
      {stage2_1[9]}
   );
   gpc1_1 gpc904 (
      {stage1_1[30]},
      {stage2_1[10]}
   );
   gpc1_1 gpc905 (
      {stage1_1[31]},
      {stage2_1[11]}
   );
   gpc1_1 gpc906 (
      {stage1_1[32]},
      {stage2_1[12]}
   );
   gpc1_1 gpc907 (
      {stage1_1[33]},
      {stage2_1[13]}
   );
   gpc1_1 gpc908 (
      {stage1_1[34]},
      {stage2_1[14]}
   );
   gpc1_1 gpc909 (
      {stage1_1[35]},
      {stage2_1[15]}
   );
   gpc1_1 gpc910 (
      {stage1_1[36]},
      {stage2_1[16]}
   );
   gpc1_1 gpc911 (
      {stage1_1[37]},
      {stage2_1[17]}
   );
   gpc1_1 gpc912 (
      {stage1_1[38]},
      {stage2_1[18]}
   );
   gpc1_1 gpc913 (
      {stage1_1[39]},
      {stage2_1[19]}
   );
   gpc1_1 gpc914 (
      {stage1_2[43]},
      {stage2_2[12]}
   );
   gpc1_1 gpc915 (
      {stage1_2[44]},
      {stage2_2[13]}
   );
   gpc1_1 gpc916 (
      {stage1_2[45]},
      {stage2_2[14]}
   );
   gpc1_1 gpc917 (
      {stage1_2[46]},
      {stage2_2[15]}
   );
   gpc1_1 gpc918 (
      {stage1_2[47]},
      {stage2_2[16]}
   );
   gpc1_1 gpc919 (
      {stage1_2[48]},
      {stage2_2[17]}
   );
   gpc1_1 gpc920 (
      {stage1_2[49]},
      {stage2_2[18]}
   );
   gpc1_1 gpc921 (
      {stage1_2[50]},
      {stage2_2[19]}
   );
   gpc1_1 gpc922 (
      {stage1_2[51]},
      {stage2_2[20]}
   );
   gpc1_1 gpc923 (
      {stage1_2[52]},
      {stage2_2[21]}
   );
   gpc1_1 gpc924 (
      {stage1_2[53]},
      {stage2_2[22]}
   );
   gpc1_1 gpc925 (
      {stage1_2[54]},
      {stage2_2[23]}
   );
   gpc1_1 gpc926 (
      {stage1_2[55]},
      {stage2_2[24]}
   );
   gpc1_1 gpc927 (
      {stage1_2[56]},
      {stage2_2[25]}
   );
   gpc1_1 gpc928 (
      {stage1_2[57]},
      {stage2_2[26]}
   );
   gpc1_1 gpc929 (
      {stage1_3[39]},
      {stage2_3[14]}
   );
   gpc1_1 gpc930 (
      {stage1_3[40]},
      {stage2_3[15]}
   );
   gpc1_1 gpc931 (
      {stage1_3[41]},
      {stage2_3[16]}
   );
   gpc1_1 gpc932 (
      {stage1_3[42]},
      {stage2_3[17]}
   );
   gpc1_1 gpc933 (
      {stage1_3[43]},
      {stage2_3[18]}
   );
   gpc1_1 gpc934 (
      {stage1_3[44]},
      {stage2_3[19]}
   );
   gpc1_1 gpc935 (
      {stage1_3[45]},
      {stage2_3[20]}
   );
   gpc1_1 gpc936 (
      {stage1_3[46]},
      {stage2_3[21]}
   );
   gpc1_1 gpc937 (
      {stage1_3[47]},
      {stage2_3[22]}
   );
   gpc1_1 gpc938 (
      {stage1_3[48]},
      {stage2_3[23]}
   );
   gpc1_1 gpc939 (
      {stage1_3[49]},
      {stage2_3[24]}
   );
   gpc1_1 gpc940 (
      {stage1_3[50]},
      {stage2_3[25]}
   );
   gpc1_1 gpc941 (
      {stage1_3[51]},
      {stage2_3[26]}
   );
   gpc1_1 gpc942 (
      {stage1_3[52]},
      {stage2_3[27]}
   );
   gpc1_1 gpc943 (
      {stage1_3[53]},
      {stage2_3[28]}
   );
   gpc1_1 gpc944 (
      {stage1_3[54]},
      {stage2_3[29]}
   );
   gpc1_1 gpc945 (
      {stage1_3[55]},
      {stage2_3[30]}
   );
   gpc1_1 gpc946 (
      {stage1_3[56]},
      {stage2_3[31]}
   );
   gpc1_1 gpc947 (
      {stage1_3[57]},
      {stage2_3[32]}
   );
   gpc1_1 gpc948 (
      {stage1_3[58]},
      {stage2_3[33]}
   );
   gpc1_1 gpc949 (
      {stage1_4[56]},
      {stage2_4[15]}
   );
   gpc1_1 gpc950 (
      {stage1_4[57]},
      {stage2_4[16]}
   );
   gpc1_1 gpc951 (
      {stage1_4[58]},
      {stage2_4[17]}
   );
   gpc1_1 gpc952 (
      {stage1_4[59]},
      {stage2_4[18]}
   );
   gpc1_1 gpc953 (
      {stage1_4[60]},
      {stage2_4[19]}
   );
   gpc1_1 gpc954 (
      {stage1_4[61]},
      {stage2_4[20]}
   );
   gpc1_1 gpc955 (
      {stage1_4[62]},
      {stage2_4[21]}
   );
   gpc1_1 gpc956 (
      {stage1_4[63]},
      {stage2_4[22]}
   );
   gpc1_1 gpc957 (
      {stage1_4[64]},
      {stage2_4[23]}
   );
   gpc1_1 gpc958 (
      {stage1_4[65]},
      {stage2_4[24]}
   );
   gpc1_1 gpc959 (
      {stage1_4[66]},
      {stage2_4[25]}
   );
   gpc1_1 gpc960 (
      {stage1_5[54]},
      {stage2_5[22]}
   );
   gpc1_1 gpc961 (
      {stage1_5[55]},
      {stage2_5[23]}
   );
   gpc1_1 gpc962 (
      {stage1_5[56]},
      {stage2_5[24]}
   );
   gpc1_1 gpc963 (
      {stage1_5[57]},
      {stage2_5[25]}
   );
   gpc1_1 gpc964 (
      {stage1_5[58]},
      {stage2_5[26]}
   );
   gpc1_1 gpc965 (
      {stage1_5[59]},
      {stage2_5[27]}
   );
   gpc1_1 gpc966 (
      {stage1_5[60]},
      {stage2_5[28]}
   );
   gpc1_1 gpc967 (
      {stage1_5[61]},
      {stage2_5[29]}
   );
   gpc1_1 gpc968 (
      {stage1_5[62]},
      {stage2_5[30]}
   );
   gpc1_1 gpc969 (
      {stage1_6[23]},
      {stage2_6[21]}
   );
   gpc1_1 gpc970 (
      {stage1_6[24]},
      {stage2_6[22]}
   );
   gpc1_1 gpc971 (
      {stage1_6[25]},
      {stage2_6[23]}
   );
   gpc1_1 gpc972 (
      {stage1_6[26]},
      {stage2_6[24]}
   );
   gpc1_1 gpc973 (
      {stage1_6[27]},
      {stage2_6[25]}
   );
   gpc1_1 gpc974 (
      {stage1_6[28]},
      {stage2_6[26]}
   );
   gpc1_1 gpc975 (
      {stage1_6[29]},
      {stage2_6[27]}
   );
   gpc1_1 gpc976 (
      {stage1_6[30]},
      {stage2_6[28]}
   );
   gpc1_1 gpc977 (
      {stage1_6[31]},
      {stage2_6[29]}
   );
   gpc1_1 gpc978 (
      {stage1_6[32]},
      {stage2_6[30]}
   );
   gpc1_1 gpc979 (
      {stage1_6[33]},
      {stage2_6[31]}
   );
   gpc1_1 gpc980 (
      {stage1_6[34]},
      {stage2_6[32]}
   );
   gpc1_1 gpc981 (
      {stage1_6[35]},
      {stage2_6[33]}
   );
   gpc1_1 gpc982 (
      {stage1_6[36]},
      {stage2_6[34]}
   );
   gpc1_1 gpc983 (
      {stage1_6[37]},
      {stage2_6[35]}
   );
   gpc1_1 gpc984 (
      {stage1_6[38]},
      {stage2_6[36]}
   );
   gpc1_1 gpc985 (
      {stage1_6[39]},
      {stage2_6[37]}
   );
   gpc1_1 gpc986 (
      {stage1_6[40]},
      {stage2_6[38]}
   );
   gpc1_1 gpc987 (
      {stage1_6[41]},
      {stage2_6[39]}
   );
   gpc1_1 gpc988 (
      {stage1_6[42]},
      {stage2_6[40]}
   );
   gpc1_1 gpc989 (
      {stage1_6[43]},
      {stage2_6[41]}
   );
   gpc1_1 gpc990 (
      {stage1_6[44]},
      {stage2_6[42]}
   );
   gpc1_1 gpc991 (
      {stage1_6[45]},
      {stage2_6[43]}
   );
   gpc1_1 gpc992 (
      {stage1_6[46]},
      {stage2_6[44]}
   );
   gpc1_1 gpc993 (
      {stage1_6[47]},
      {stage2_6[45]}
   );
   gpc1_1 gpc994 (
      {stage1_6[48]},
      {stage2_6[46]}
   );
   gpc1_1 gpc995 (
      {stage1_6[49]},
      {stage2_6[47]}
   );
   gpc1_1 gpc996 (
      {stage1_7[68]},
      {stage2_7[18]}
   );
   gpc1_1 gpc997 (
      {stage1_7[69]},
      {stage2_7[19]}
   );
   gpc1_1 gpc998 (
      {stage1_8[35]},
      {stage2_8[18]}
   );
   gpc1_1 gpc999 (
      {stage1_8[36]},
      {stage2_8[19]}
   );
   gpc1_1 gpc1000 (
      {stage1_8[37]},
      {stage2_8[20]}
   );
   gpc1_1 gpc1001 (
      {stage1_8[38]},
      {stage2_8[21]}
   );
   gpc1_1 gpc1002 (
      {stage1_8[39]},
      {stage2_8[22]}
   );
   gpc1_1 gpc1003 (
      {stage1_8[40]},
      {stage2_8[23]}
   );
   gpc1_1 gpc1004 (
      {stage1_8[41]},
      {stage2_8[24]}
   );
   gpc1_1 gpc1005 (
      {stage1_8[42]},
      {stage2_8[25]}
   );
   gpc1_1 gpc1006 (
      {stage1_8[43]},
      {stage2_8[26]}
   );
   gpc1_1 gpc1007 (
      {stage1_8[44]},
      {stage2_8[27]}
   );
   gpc1_1 gpc1008 (
      {stage1_8[45]},
      {stage2_8[28]}
   );
   gpc1_1 gpc1009 (
      {stage1_8[46]},
      {stage2_8[29]}
   );
   gpc1_1 gpc1010 (
      {stage1_8[47]},
      {stage2_8[30]}
   );
   gpc1_1 gpc1011 (
      {stage1_8[48]},
      {stage2_8[31]}
   );
   gpc1_1 gpc1012 (
      {stage1_8[49]},
      {stage2_8[32]}
   );
   gpc1_1 gpc1013 (
      {stage1_8[50]},
      {stage2_8[33]}
   );
   gpc1_1 gpc1014 (
      {stage1_8[51]},
      {stage2_8[34]}
   );
   gpc1_1 gpc1015 (
      {stage1_8[52]},
      {stage2_8[35]}
   );
   gpc1_1 gpc1016 (
      {stage1_8[53]},
      {stage2_8[36]}
   );
   gpc1_1 gpc1017 (
      {stage1_8[54]},
      {stage2_8[37]}
   );
   gpc1_1 gpc1018 (
      {stage1_8[55]},
      {stage2_8[38]}
   );
   gpc1_1 gpc1019 (
      {stage1_9[60]},
      {stage2_9[22]}
   );
   gpc1_1 gpc1020 (
      {stage1_11[55]},
      {stage2_11[24]}
   );
   gpc1_1 gpc1021 (
      {stage1_11[56]},
      {stage2_11[25]}
   );
   gpc1_1 gpc1022 (
      {stage1_11[57]},
      {stage2_11[26]}
   );
   gpc1_1 gpc1023 (
      {stage1_13[48]},
      {stage2_13[22]}
   );
   gpc1_1 gpc1024 (
      {stage1_13[49]},
      {stage2_13[23]}
   );
   gpc1_1 gpc1025 (
      {stage1_13[50]},
      {stage2_13[24]}
   );
   gpc1_1 gpc1026 (
      {stage1_13[51]},
      {stage2_13[25]}
   );
   gpc1_1 gpc1027 (
      {stage1_13[52]},
      {stage2_13[26]}
   );
   gpc1_1 gpc1028 (
      {stage1_13[53]},
      {stage2_13[27]}
   );
   gpc1_1 gpc1029 (
      {stage1_13[54]},
      {stage2_13[28]}
   );
   gpc1_1 gpc1030 (
      {stage1_13[55]},
      {stage2_13[29]}
   );
   gpc1_1 gpc1031 (
      {stage1_13[56]},
      {stage2_13[30]}
   );
   gpc1_1 gpc1032 (
      {stage1_13[57]},
      {stage2_13[31]}
   );
   gpc1_1 gpc1033 (
      {stage1_13[58]},
      {stage2_13[32]}
   );
   gpc1_1 gpc1034 (
      {stage1_13[59]},
      {stage2_13[33]}
   );
   gpc1_1 gpc1035 (
      {stage1_13[60]},
      {stage2_13[34]}
   );
   gpc1_1 gpc1036 (
      {stage1_14[42]},
      {stage2_14[23]}
   );
   gpc1_1 gpc1037 (
      {stage1_14[43]},
      {stage2_14[24]}
   );
   gpc1_1 gpc1038 (
      {stage1_14[44]},
      {stage2_14[25]}
   );
   gpc1_1 gpc1039 (
      {stage1_14[45]},
      {stage2_14[26]}
   );
   gpc1_1 gpc1040 (
      {stage1_15[44]},
      {stage2_15[20]}
   );
   gpc1_1 gpc1041 (
      {stage1_15[45]},
      {stage2_15[21]}
   );
   gpc1_1 gpc1042 (
      {stage1_15[46]},
      {stage2_15[22]}
   );
   gpc1_1 gpc1043 (
      {stage1_17[37]},
      {stage2_17[23]}
   );
   gpc1_1 gpc1044 (
      {stage1_17[38]},
      {stage2_17[24]}
   );
   gpc1_1 gpc1045 (
      {stage1_17[39]},
      {stage2_17[25]}
   );
   gpc1_1 gpc1046 (
      {stage1_17[40]},
      {stage2_17[26]}
   );
   gpc1_1 gpc1047 (
      {stage1_17[41]},
      {stage2_17[27]}
   );
   gpc1_1 gpc1048 (
      {stage1_17[42]},
      {stage2_17[28]}
   );
   gpc1_1 gpc1049 (
      {stage1_17[43]},
      {stage2_17[29]}
   );
   gpc1_1 gpc1050 (
      {stage1_17[44]},
      {stage2_17[30]}
   );
   gpc1_1 gpc1051 (
      {stage1_17[45]},
      {stage2_17[31]}
   );
   gpc1_1 gpc1052 (
      {stage1_17[46]},
      {stage2_17[32]}
   );
   gpc1_1 gpc1053 (
      {stage1_17[47]},
      {stage2_17[33]}
   );
   gpc1_1 gpc1054 (
      {stage1_17[48]},
      {stage2_17[34]}
   );
   gpc1_1 gpc1055 (
      {stage1_17[49]},
      {stage2_17[35]}
   );
   gpc1_1 gpc1056 (
      {stage1_17[50]},
      {stage2_17[36]}
   );
   gpc1_1 gpc1057 (
      {stage1_17[51]},
      {stage2_17[37]}
   );
   gpc1_1 gpc1058 (
      {stage1_17[52]},
      {stage2_17[38]}
   );
   gpc1_1 gpc1059 (
      {stage1_17[53]},
      {stage2_17[39]}
   );
   gpc1_1 gpc1060 (
      {stage1_17[54]},
      {stage2_17[40]}
   );
   gpc1_1 gpc1061 (
      {stage1_17[55]},
      {stage2_17[41]}
   );
   gpc1_1 gpc1062 (
      {stage1_17[56]},
      {stage2_17[42]}
   );
   gpc1_1 gpc1063 (
      {stage1_17[57]},
      {stage2_17[43]}
   );
   gpc1_1 gpc1064 (
      {stage1_17[58]},
      {stage2_17[44]}
   );
   gpc1_1 gpc1065 (
      {stage1_17[59]},
      {stage2_17[45]}
   );
   gpc1_1 gpc1066 (
      {stage1_17[60]},
      {stage2_17[46]}
   );
   gpc1_1 gpc1067 (
      {stage1_17[61]},
      {stage2_17[47]}
   );
   gpc1_1 gpc1068 (
      {stage1_17[62]},
      {stage2_17[48]}
   );
   gpc1_1 gpc1069 (
      {stage1_18[48]},
      {stage2_18[20]}
   );
   gpc1_1 gpc1070 (
      {stage1_18[49]},
      {stage2_18[21]}
   );
   gpc1_1 gpc1071 (
      {stage1_18[50]},
      {stage2_18[22]}
   );
   gpc1_1 gpc1072 (
      {stage1_18[51]},
      {stage2_18[23]}
   );
   gpc1_1 gpc1073 (
      {stage1_18[52]},
      {stage2_18[24]}
   );
   gpc1_1 gpc1074 (
      {stage1_18[53]},
      {stage2_18[25]}
   );
   gpc1_1 gpc1075 (
      {stage1_18[54]},
      {stage2_18[26]}
   );
   gpc1_1 gpc1076 (
      {stage1_18[55]},
      {stage2_18[27]}
   );
   gpc1_1 gpc1077 (
      {stage1_18[56]},
      {stage2_18[28]}
   );
   gpc1_1 gpc1078 (
      {stage1_18[57]},
      {stage2_18[29]}
   );
   gpc1_1 gpc1079 (
      {stage1_18[58]},
      {stage2_18[30]}
   );
   gpc1_1 gpc1080 (
      {stage1_18[59]},
      {stage2_18[31]}
   );
   gpc1_1 gpc1081 (
      {stage1_18[60]},
      {stage2_18[32]}
   );
   gpc1_1 gpc1082 (
      {stage1_18[61]},
      {stage2_18[33]}
   );
   gpc1_1 gpc1083 (
      {stage1_18[62]},
      {stage2_18[34]}
   );
   gpc1_1 gpc1084 (
      {stage1_18[63]},
      {stage2_18[35]}
   );
   gpc1_1 gpc1085 (
      {stage1_18[64]},
      {stage2_18[36]}
   );
   gpc1_1 gpc1086 (
      {stage1_18[65]},
      {stage2_18[37]}
   );
   gpc1_1 gpc1087 (
      {stage1_19[42]},
      {stage2_19[20]}
   );
   gpc1_1 gpc1088 (
      {stage1_20[30]},
      {stage2_20[20]}
   );
   gpc1_1 gpc1089 (
      {stage1_20[31]},
      {stage2_20[21]}
   );
   gpc1_1 gpc1090 (
      {stage1_20[32]},
      {stage2_20[22]}
   );
   gpc1_1 gpc1091 (
      {stage1_20[33]},
      {stage2_20[23]}
   );
   gpc1_1 gpc1092 (
      {stage1_20[34]},
      {stage2_20[24]}
   );
   gpc1_1 gpc1093 (
      {stage1_20[35]},
      {stage2_20[25]}
   );
   gpc1_1 gpc1094 (
      {stage1_20[36]},
      {stage2_20[26]}
   );
   gpc1_1 gpc1095 (
      {stage1_20[37]},
      {stage2_20[27]}
   );
   gpc1_1 gpc1096 (
      {stage1_20[38]},
      {stage2_20[28]}
   );
   gpc1_1 gpc1097 (
      {stage1_20[39]},
      {stage2_20[29]}
   );
   gpc1_1 gpc1098 (
      {stage1_20[40]},
      {stage2_20[30]}
   );
   gpc1_1 gpc1099 (
      {stage1_20[41]},
      {stage2_20[31]}
   );
   gpc1_1 gpc1100 (
      {stage1_20[42]},
      {stage2_20[32]}
   );
   gpc1_1 gpc1101 (
      {stage1_20[43]},
      {stage2_20[33]}
   );
   gpc1_1 gpc1102 (
      {stage1_20[44]},
      {stage2_20[34]}
   );
   gpc1_1 gpc1103 (
      {stage1_20[45]},
      {stage2_20[35]}
   );
   gpc1_1 gpc1104 (
      {stage1_20[46]},
      {stage2_20[36]}
   );
   gpc1_1 gpc1105 (
      {stage1_20[47]},
      {stage2_20[37]}
   );
   gpc1_1 gpc1106 (
      {stage1_20[48]},
      {stage2_20[38]}
   );
   gpc1_1 gpc1107 (
      {stage1_20[49]},
      {stage2_20[39]}
   );
   gpc1_1 gpc1108 (
      {stage1_20[50]},
      {stage2_20[40]}
   );
   gpc1_1 gpc1109 (
      {stage1_20[51]},
      {stage2_20[41]}
   );
   gpc1_1 gpc1110 (
      {stage1_20[52]},
      {stage2_20[42]}
   );
   gpc1_1 gpc1111 (
      {stage1_20[53]},
      {stage2_20[43]}
   );
   gpc1_1 gpc1112 (
      {stage1_20[54]},
      {stage2_20[44]}
   );
   gpc1_1 gpc1113 (
      {stage1_20[55]},
      {stage2_20[45]}
   );
   gpc1_1 gpc1114 (
      {stage1_20[56]},
      {stage2_20[46]}
   );
   gpc1_1 gpc1115 (
      {stage1_20[57]},
      {stage2_20[47]}
   );
   gpc1_1 gpc1116 (
      {stage1_20[58]},
      {stage2_20[48]}
   );
   gpc1_1 gpc1117 (
      {stage1_20[59]},
      {stage2_20[49]}
   );
   gpc1_1 gpc1118 (
      {stage1_20[60]},
      {stage2_20[50]}
   );
   gpc1_1 gpc1119 (
      {stage1_20[61]},
      {stage2_20[51]}
   );
   gpc1_1 gpc1120 (
      {stage1_20[62]},
      {stage2_20[52]}
   );
   gpc1_1 gpc1121 (
      {stage1_20[63]},
      {stage2_20[53]}
   );
   gpc1_1 gpc1122 (
      {stage1_20[64]},
      {stage2_20[54]}
   );
   gpc1_1 gpc1123 (
      {stage1_20[65]},
      {stage2_20[55]}
   );
   gpc1_1 gpc1124 (
      {stage1_21[60]},
      {stage2_21[16]}
   );
   gpc1_1 gpc1125 (
      {stage1_21[61]},
      {stage2_21[17]}
   );
   gpc1_1 gpc1126 (
      {stage1_21[62]},
      {stage2_21[18]}
   );
   gpc1_1 gpc1127 (
      {stage1_21[63]},
      {stage2_21[19]}
   );
   gpc1_1 gpc1128 (
      {stage1_21[64]},
      {stage2_21[20]}
   );
   gpc1_1 gpc1129 (
      {stage1_22[53]},
      {stage2_22[19]}
   );
   gpc1_1 gpc1130 (
      {stage1_22[54]},
      {stage2_22[20]}
   );
   gpc1_1 gpc1131 (
      {stage1_22[55]},
      {stage2_22[21]}
   );
   gpc1_1 gpc1132 (
      {stage1_22[56]},
      {stage2_22[22]}
   );
   gpc1_1 gpc1133 (
      {stage1_22[57]},
      {stage2_22[23]}
   );
   gpc1_1 gpc1134 (
      {stage1_22[58]},
      {stage2_22[24]}
   );
   gpc1_1 gpc1135 (
      {stage1_22[59]},
      {stage2_22[25]}
   );
   gpc1_1 gpc1136 (
      {stage1_22[60]},
      {stage2_22[26]}
   );
   gpc1_1 gpc1137 (
      {stage1_23[30]},
      {stage2_23[20]}
   );
   gpc1_1 gpc1138 (
      {stage1_23[31]},
      {stage2_23[21]}
   );
   gpc1_1 gpc1139 (
      {stage1_23[32]},
      {stage2_23[22]}
   );
   gpc1_1 gpc1140 (
      {stage1_23[33]},
      {stage2_23[23]}
   );
   gpc1_1 gpc1141 (
      {stage1_23[34]},
      {stage2_23[24]}
   );
   gpc1_1 gpc1142 (
      {stage1_23[35]},
      {stage2_23[25]}
   );
   gpc1_1 gpc1143 (
      {stage1_23[36]},
      {stage2_23[26]}
   );
   gpc1_1 gpc1144 (
      {stage1_23[37]},
      {stage2_23[27]}
   );
   gpc1_1 gpc1145 (
      {stage1_23[38]},
      {stage2_23[28]}
   );
   gpc1_1 gpc1146 (
      {stage1_23[39]},
      {stage2_23[29]}
   );
   gpc1_1 gpc1147 (
      {stage1_23[40]},
      {stage2_23[30]}
   );
   gpc1_1 gpc1148 (
      {stage1_23[41]},
      {stage2_23[31]}
   );
   gpc1_1 gpc1149 (
      {stage1_23[42]},
      {stage2_23[32]}
   );
   gpc1_1 gpc1150 (
      {stage1_23[43]},
      {stage2_23[33]}
   );
   gpc1_1 gpc1151 (
      {stage1_24[79]},
      {stage2_24[22]}
   );
   gpc1_1 gpc1152 (
      {stage1_24[80]},
      {stage2_24[23]}
   );
   gpc1_1 gpc1153 (
      {stage1_24[81]},
      {stage2_24[24]}
   );
   gpc1_1 gpc1154 (
      {stage1_24[82]},
      {stage2_24[25]}
   );
   gpc1_1 gpc1155 (
      {stage1_24[83]},
      {stage2_24[26]}
   );
   gpc1_1 gpc1156 (
      {stage1_24[84]},
      {stage2_24[27]}
   );
   gpc1_1 gpc1157 (
      {stage1_24[85]},
      {stage2_24[28]}
   );
   gpc1_1 gpc1158 (
      {stage1_24[86]},
      {stage2_24[29]}
   );
   gpc1_1 gpc1159 (
      {stage1_24[87]},
      {stage2_24[30]}
   );
   gpc1_1 gpc1160 (
      {stage1_24[88]},
      {stage2_24[31]}
   );
   gpc1_1 gpc1161 (
      {stage1_24[89]},
      {stage2_24[32]}
   );
   gpc1_1 gpc1162 (
      {stage1_25[48]},
      {stage2_25[25]}
   );
   gpc1_1 gpc1163 (
      {stage1_25[49]},
      {stage2_25[26]}
   );
   gpc1_1 gpc1164 (
      {stage1_25[50]},
      {stage2_25[27]}
   );
   gpc1_1 gpc1165 (
      {stage1_25[51]},
      {stage2_25[28]}
   );
   gpc1_1 gpc1166 (
      {stage1_25[52]},
      {stage2_25[29]}
   );
   gpc1_1 gpc1167 (
      {stage1_25[53]},
      {stage2_25[30]}
   );
   gpc1_1 gpc1168 (
      {stage1_25[54]},
      {stage2_25[31]}
   );
   gpc1_1 gpc1169 (
      {stage1_25[55]},
      {stage2_25[32]}
   );
   gpc1_1 gpc1170 (
      {stage1_25[56]},
      {stage2_25[33]}
   );
   gpc1_1 gpc1171 (
      {stage1_25[57]},
      {stage2_25[34]}
   );
   gpc1_1 gpc1172 (
      {stage1_25[58]},
      {stage2_25[35]}
   );
   gpc1_1 gpc1173 (
      {stage1_25[59]},
      {stage2_25[36]}
   );
   gpc1_1 gpc1174 (
      {stage1_25[60]},
      {stage2_25[37]}
   );
   gpc1_1 gpc1175 (
      {stage1_25[61]},
      {stage2_25[38]}
   );
   gpc1_1 gpc1176 (
      {stage1_25[62]},
      {stage2_25[39]}
   );
   gpc1_1 gpc1177 (
      {stage1_25[63]},
      {stage2_25[40]}
   );
   gpc1_1 gpc1178 (
      {stage1_25[64]},
      {stage2_25[41]}
   );
   gpc1_1 gpc1179 (
      {stage1_25[65]},
      {stage2_25[42]}
   );
   gpc1_1 gpc1180 (
      {stage1_25[66]},
      {stage2_25[43]}
   );
   gpc1_1 gpc1181 (
      {stage1_25[67]},
      {stage2_25[44]}
   );
   gpc1_1 gpc1182 (
      {stage1_25[68]},
      {stage2_25[45]}
   );
   gpc1_1 gpc1183 (
      {stage1_25[69]},
      {stage2_25[46]}
   );
   gpc1_1 gpc1184 (
      {stage1_26[54]},
      {stage2_26[22]}
   );
   gpc1_1 gpc1185 (
      {stage1_26[55]},
      {stage2_26[23]}
   );
   gpc1_1 gpc1186 (
      {stage1_26[56]},
      {stage2_26[24]}
   );
   gpc1_1 gpc1187 (
      {stage1_26[57]},
      {stage2_26[25]}
   );
   gpc1_1 gpc1188 (
      {stage1_26[58]},
      {stage2_26[26]}
   );
   gpc1_1 gpc1189 (
      {stage1_26[59]},
      {stage2_26[27]}
   );
   gpc1_1 gpc1190 (
      {stage1_26[60]},
      {stage2_26[28]}
   );
   gpc1_1 gpc1191 (
      {stage1_26[61]},
      {stage2_26[29]}
   );
   gpc1_1 gpc1192 (
      {stage1_26[62]},
      {stage2_26[30]}
   );
   gpc1_1 gpc1193 (
      {stage1_26[63]},
      {stage2_26[31]}
   );
   gpc1_1 gpc1194 (
      {stage1_26[64]},
      {stage2_26[32]}
   );
   gpc1_1 gpc1195 (
      {stage1_26[65]},
      {stage2_26[33]}
   );
   gpc1_1 gpc1196 (
      {stage1_26[66]},
      {stage2_26[34]}
   );
   gpc1_1 gpc1197 (
      {stage1_26[67]},
      {stage2_26[35]}
   );
   gpc1_1 gpc1198 (
      {stage1_26[68]},
      {stage2_26[36]}
   );
   gpc1_1 gpc1199 (
      {stage1_27[42]},
      {stage2_27[17]}
   );
   gpc1_1 gpc1200 (
      {stage1_27[43]},
      {stage2_27[18]}
   );
   gpc1_1 gpc1201 (
      {stage1_27[44]},
      {stage2_27[19]}
   );
   gpc1_1 gpc1202 (
      {stage1_27[45]},
      {stage2_27[20]}
   );
   gpc1_1 gpc1203 (
      {stage1_27[46]},
      {stage2_27[21]}
   );
   gpc1_1 gpc1204 (
      {stage1_27[47]},
      {stage2_27[22]}
   );
   gpc1_1 gpc1205 (
      {stage1_27[48]},
      {stage2_27[23]}
   );
   gpc1_1 gpc1206 (
      {stage1_27[49]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1207 (
      {stage1_27[50]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1208 (
      {stage1_27[51]},
      {stage2_27[26]}
   );
   gpc1_1 gpc1209 (
      {stage1_27[52]},
      {stage2_27[27]}
   );
   gpc1_1 gpc1210 (
      {stage1_27[53]},
      {stage2_27[28]}
   );
   gpc1_1 gpc1211 (
      {stage1_27[54]},
      {stage2_27[29]}
   );
   gpc1_1 gpc1212 (
      {stage1_27[55]},
      {stage2_27[30]}
   );
   gpc1_1 gpc1213 (
      {stage1_28[42]},
      {stage2_28[22]}
   );
   gpc1_1 gpc1214 (
      {stage1_28[43]},
      {stage2_28[23]}
   );
   gpc1_1 gpc1215 (
      {stage1_28[44]},
      {stage2_28[24]}
   );
   gpc1_1 gpc1216 (
      {stage1_28[45]},
      {stage2_28[25]}
   );
   gpc1_1 gpc1217 (
      {stage1_28[46]},
      {stage2_28[26]}
   );
   gpc1_1 gpc1218 (
      {stage1_28[47]},
      {stage2_28[27]}
   );
   gpc1_1 gpc1219 (
      {stage1_28[48]},
      {stage2_28[28]}
   );
   gpc1_1 gpc1220 (
      {stage1_28[49]},
      {stage2_28[29]}
   );
   gpc1_1 gpc1221 (
      {stage1_28[50]},
      {stage2_28[30]}
   );
   gpc1_1 gpc1222 (
      {stage1_28[51]},
      {stage2_28[31]}
   );
   gpc1_1 gpc1223 (
      {stage1_28[52]},
      {stage2_28[32]}
   );
   gpc1_1 gpc1224 (
      {stage1_28[53]},
      {stage2_28[33]}
   );
   gpc1_1 gpc1225 (
      {stage1_28[54]},
      {stage2_28[34]}
   );
   gpc1_1 gpc1226 (
      {stage1_28[55]},
      {stage2_28[35]}
   );
   gpc1_1 gpc1227 (
      {stage1_29[47]},
      {stage2_29[22]}
   );
   gpc1_1 gpc1228 (
      {stage1_29[48]},
      {stage2_29[23]}
   );
   gpc1_1 gpc1229 (
      {stage1_29[49]},
      {stage2_29[24]}
   );
   gpc1_1 gpc1230 (
      {stage1_29[50]},
      {stage2_29[25]}
   );
   gpc1_1 gpc1231 (
      {stage1_29[51]},
      {stage2_29[26]}
   );
   gpc1_1 gpc1232 (
      {stage1_29[52]},
      {stage2_29[27]}
   );
   gpc1_1 gpc1233 (
      {stage1_29[53]},
      {stage2_29[28]}
   );
   gpc1_1 gpc1234 (
      {stage1_29[54]},
      {stage2_29[29]}
   );
   gpc1_1 gpc1235 (
      {stage1_29[55]},
      {stage2_29[30]}
   );
   gpc1_1 gpc1236 (
      {stage1_29[56]},
      {stage2_29[31]}
   );
   gpc1_1 gpc1237 (
      {stage1_31[57]},
      {stage2_31[20]}
   );
   gpc1_1 gpc1238 (
      {stage1_31[58]},
      {stage2_31[21]}
   );
   gpc1_1 gpc1239 (
      {stage1_31[59]},
      {stage2_31[22]}
   );
   gpc1_1 gpc1240 (
      {stage1_31[60]},
      {stage2_31[23]}
   );
   gpc1_1 gpc1241 (
      {stage1_31[61]},
      {stage2_31[24]}
   );
   gpc1_1 gpc1242 (
      {stage1_31[62]},
      {stage2_31[25]}
   );
   gpc1_1 gpc1243 (
      {stage1_31[63]},
      {stage2_31[26]}
   );
   gpc1_1 gpc1244 (
      {stage1_31[64]},
      {stage2_31[27]}
   );
   gpc1_1 gpc1245 (
      {stage1_31[65]},
      {stage2_31[28]}
   );
   gpc1_1 gpc1246 (
      {stage1_31[66]},
      {stage2_31[29]}
   );
   gpc1_1 gpc1247 (
      {stage1_31[67]},
      {stage2_31[30]}
   );
   gpc1_1 gpc1248 (
      {stage1_31[68]},
      {stage2_31[31]}
   );
   gpc1_1 gpc1249 (
      {stage1_31[69]},
      {stage2_31[32]}
   );
   gpc1_1 gpc1250 (
      {stage1_31[70]},
      {stage2_31[33]}
   );
   gpc1_1 gpc1251 (
      {stage1_32[25]},
      {stage2_32[20]}
   );
   gpc1_1 gpc1252 (
      {stage1_32[26]},
      {stage2_32[21]}
   );
   gpc1_1 gpc1253 (
      {stage1_32[27]},
      {stage2_32[22]}
   );
   gpc1_1 gpc1254 (
      {stage1_32[28]},
      {stage2_32[23]}
   );
   gpc1_1 gpc1255 (
      {stage1_32[29]},
      {stage2_32[24]}
   );
   gpc1_1 gpc1256 (
      {stage1_32[30]},
      {stage2_32[25]}
   );
   gpc1_1 gpc1257 (
      {stage1_32[31]},
      {stage2_32[26]}
   );
   gpc1_1 gpc1258 (
      {stage1_32[32]},
      {stage2_32[27]}
   );
   gpc1_1 gpc1259 (
      {stage1_32[33]},
      {stage2_32[28]}
   );
   gpc1_1 gpc1260 (
      {stage1_33[12]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1261 (
      {stage1_33[13]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1262 (
      {stage1_33[14]},
      {stage2_33[16]}
   );
   gpc1_1 gpc1263 (
      {stage1_33[15]},
      {stage2_33[17]}
   );
   gpc2135_5 gpc1264 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc2135_5 gpc1265 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[1]},
      {stage2_3[2], stage2_3[3]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc2135_5 gpc1266 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_2[2]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc2135_5 gpc1267 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19]},
      {stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[3]},
      {stage2_3[6], stage2_3[7]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1268 (
      {stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24], stage2_0[25]},
      {stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc615_5 gpc1269 (
      {stage2_0[26], stage2_0[27], stage2_0[28], stage2_0[29], stage2_0[30]},
      {stage2_1[12]},
      {stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc615_5 gpc1270 (
      {stage2_0[31], stage2_0[32], stage2_0[33], stage2_0[34], stage2_0[35]},
      {stage2_1[13]},
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc615_5 gpc1271 (
      {stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25], stage2_2[26]},
      {stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc1272 (
      {stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc1273 (
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[2],stage3_4[9],stage3_3[9]}
   );
   gpc615_5 gpc1274 (
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[3],stage3_4[10],stage3_3[10]}
   );
   gpc615_5 gpc1275 (
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28]},
      {stage2_4[9]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[4],stage3_5[4],stage3_4[11],stage3_3[11]}
   );
   gpc615_5 gpc1276 (
      {stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_4[10]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[5],stage3_5[5],stage3_4[12],stage3_3[12]}
   );
   gpc606_5 gpc1277 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[5],stage3_6[6],stage3_5[6],stage3_4[13]}
   );
   gpc606_5 gpc1278 (
      {stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[6],stage3_6[7],stage3_5[7],stage3_4[14]}
   );
   gpc606_5 gpc1279 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[7],stage3_6[8]}
   );
   gpc606_5 gpc1280 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[8],stage3_6[9]}
   );
   gpc606_5 gpc1281 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[4],stage3_7[9]}
   );
   gpc615_5 gpc1282 (
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10]},
      {stage2_8[12]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[5],stage3_7[10]}
   );
   gpc615_5 gpc1283 (
      {stage2_7[11], stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15]},
      {stage2_8[13]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[6],stage3_7[11]}
   );
   gpc615_5 gpc1284 (
      {stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19], 1'b0},
      {stage2_8[14]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], 1'b0},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[7],stage3_7[12]}
   );
   gpc606_5 gpc1285 (
      {stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[8]}
   );
   gpc606_5 gpc1286 (
      {stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[9]}
   );
   gpc606_5 gpc1287 (
      {stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31], stage2_8[32]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[8],stage3_9[8],stage3_8[10]}
   );
   gpc615_5 gpc1288 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[7]}
   );
   gpc615_5 gpc1289 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage2_12[1]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[8]}
   );
   gpc615_5 gpc1290 (
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[2]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[9]}
   );
   gpc615_5 gpc1291 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[3]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6],stage3_11[10]}
   );
   gpc615_5 gpc1292 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[4]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[4],stage3_12[7],stage3_11[11]}
   );
   gpc606_5 gpc1293 (
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[5],stage3_13[5],stage3_12[8]}
   );
   gpc606_5 gpc1294 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[6],stage3_14[6]}
   );
   gpc615_5 gpc1295 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[7]}
   );
   gpc615_5 gpc1296 (
      {stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[8]}
   );
   gpc615_5 gpc1297 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[3],stage3_16[4],stage3_15[9]}
   );
   gpc615_5 gpc1298 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[4],stage3_16[5],stage3_15[10]}
   );
   gpc615_5 gpc1299 (
      {stage2_15[20], stage2_15[21], stage2_15[22], 1'b0, 1'b0},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[5],stage3_16[6],stage3_15[11]}
   );
   gpc117_4 gpc1300 (
      {stage2_16[11], stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_17[30]},
      {stage2_18[0]},
      {stage3_19[5],stage3_18[6],stage3_17[6],stage3_16[7]}
   );
   gpc606_5 gpc1301 (
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[0],stage3_19[6],stage3_18[7]}
   );
   gpc606_5 gpc1302 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[1],stage3_19[7],stage3_18[8]}
   );
   gpc606_5 gpc1303 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[2],stage3_19[8],stage3_18[9]}
   );
   gpc615_5 gpc1304 (
      {stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage2_19[0]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[3],stage3_19[9],stage3_18[10]}
   );
   gpc615_5 gpc1305 (
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28]},
      {stage2_19[1]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[4],stage3_19[10],stage3_18[11]}
   );
   gpc615_5 gpc1306 (
      {stage2_18[29], stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33]},
      {stage2_19[2]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[5],stage3_19[11],stage3_18[12]}
   );
   gpc615_5 gpc1307 (
      {stage2_18[34], stage2_18[35], stage2_18[36], stage2_18[37], 1'b0},
      {stage2_19[3]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[6],stage3_19[12],stage3_18[13]}
   );
   gpc615_5 gpc1308 (
      {stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[42]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[7],stage3_21[7],stage3_20[7],stage3_19[13]}
   );
   gpc606_5 gpc1309 (
      {stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47], stage2_20[48]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[1],stage3_22[8],stage3_21[8],stage3_20[8]}
   );
   gpc606_5 gpc1310 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[2],stage3_22[9],stage3_21[9]}
   );
   gpc606_5 gpc1311 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[3],stage3_22[10],stage3_21[10]}
   );
   gpc615_5 gpc1312 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[3],stage3_23[4],stage3_22[11]}
   );
   gpc615_5 gpc1313 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[4],stage3_23[5],stage3_22[12]}
   );
   gpc615_5 gpc1314 (
      {stage2_22[16], stage2_22[17], stage2_22[18], stage2_22[19], stage2_22[20]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[5],stage3_23[6],stage3_22[13]}
   );
   gpc615_5 gpc1315 (
      {stage2_22[21], stage2_22[22], stage2_22[23], stage2_22[24], stage2_22[25]},
      {stage2_23[15]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[5],stage3_24[6],stage3_23[7],stage3_22[14]}
   );
   gpc606_5 gpc1316 (
      {stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[4],stage3_25[6],stage3_24[7],stage3_23[8]}
   );
   gpc606_5 gpc1317 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[5],stage3_25[7],stage3_24[8],stage3_23[9]}
   );
   gpc606_5 gpc1318 (
      {stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[6],stage3_25[8],stage3_24[9],stage3_23[10]}
   );
   gpc606_5 gpc1319 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[3],stage3_26[7],stage3_25[9]}
   );
   gpc606_5 gpc1320 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[1],stage3_27[4],stage3_26[8],stage3_25[10]}
   );
   gpc606_5 gpc1321 (
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[2],stage3_27[5],stage3_26[9],stage3_25[11]}
   );
   gpc606_5 gpc1322 (
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[3],stage3_27[6],stage3_26[10],stage3_25[12]}
   );
   gpc615_5 gpc1323 (
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46]},
      {stage2_26[0]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[4],stage3_27[7],stage3_26[11],stage3_25[13]}
   );
   gpc606_5 gpc1324 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[5],stage3_28[5],stage3_27[8],stage3_26[12]}
   );
   gpc606_5 gpc1325 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[6],stage3_28[6],stage3_27[9],stage3_26[13]}
   );
   gpc606_5 gpc1326 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[7],stage3_28[7],stage3_27[10],stage3_26[14]}
   );
   gpc606_5 gpc1327 (
      {stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24]},
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage3_30[3],stage3_29[8],stage3_28[8],stage3_27[11],stage3_26[15]}
   );
   gpc606_5 gpc1328 (
      {stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30]},
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28], stage2_28[29]},
      {stage3_30[4],stage3_29[9],stage3_28[9],stage3_27[12],stage3_26[16]}
   );
   gpc615_5 gpc1329 (
      {stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage2_27[30]},
      {stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35]},
      {stage3_30[5],stage3_29[10],stage3_28[10],stage3_27[13],stage3_26[17]}
   );
   gpc606_5 gpc1330 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[6],stage3_29[11]}
   );
   gpc606_5 gpc1331 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[1],stage3_31[1],stage3_30[7],stage3_29[12]}
   );
   gpc606_5 gpc1332 (
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[2],stage3_31[2],stage3_30[8],stage3_29[13]}
   );
   gpc606_5 gpc1333 (
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[3],stage3_31[3],stage3_30[9],stage3_29[14]}
   );
   gpc606_5 gpc1334 (
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[4],stage3_31[4],stage3_30[10],stage3_29[15]}
   );
   gpc606_5 gpc1335 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[5],stage3_32[5],stage3_31[5],stage3_30[11]}
   );
   gpc606_5 gpc1336 (
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[6],stage3_32[6],stage3_31[6],stage3_30[12]}
   );
   gpc606_5 gpc1337 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[7],stage3_32[7],stage3_31[7],stage3_30[13]}
   );
   gpc1415_5 gpc1338 (
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], 1'b0},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3]},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[3],stage3_33[8],stage3_32[8],stage3_31[8]}
   );
   gpc2135_5 gpc1339 (
      {stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage2_34[1]},
      {stage2_35[0], stage2_35[1]},
      {stage3_36[0],stage3_35[1],stage3_34[4],stage3_33[9],stage3_32[9]}
   );
   gpc1_1 gpc1340 (
      {stage2_1[14]},
      {stage3_1[7]}
   );
   gpc1_1 gpc1341 (
      {stage2_1[15]},
      {stage3_1[8]}
   );
   gpc1_1 gpc1342 (
      {stage2_1[16]},
      {stage3_1[9]}
   );
   gpc1_1 gpc1343 (
      {stage2_1[17]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1344 (
      {stage2_1[18]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1345 (
      {stage2_1[19]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1346 (
      {stage2_4[23]},
      {stage3_4[15]}
   );
   gpc1_1 gpc1347 (
      {stage2_4[24]},
      {stage3_4[16]}
   );
   gpc1_1 gpc1348 (
      {stage2_4[25]},
      {stage3_4[17]}
   );
   gpc1_1 gpc1349 (
      {stage2_5[30]},
      {stage3_5[8]}
   );
   gpc1_1 gpc1350 (
      {stage2_6[24]},
      {stage3_6[10]}
   );
   gpc1_1 gpc1351 (
      {stage2_6[25]},
      {stage3_6[11]}
   );
   gpc1_1 gpc1352 (
      {stage2_6[26]},
      {stage3_6[12]}
   );
   gpc1_1 gpc1353 (
      {stage2_6[27]},
      {stage3_6[13]}
   );
   gpc1_1 gpc1354 (
      {stage2_6[28]},
      {stage3_6[14]}
   );
   gpc1_1 gpc1355 (
      {stage2_6[29]},
      {stage3_6[15]}
   );
   gpc1_1 gpc1356 (
      {stage2_6[30]},
      {stage3_6[16]}
   );
   gpc1_1 gpc1357 (
      {stage2_6[31]},
      {stage3_6[17]}
   );
   gpc1_1 gpc1358 (
      {stage2_6[32]},
      {stage3_6[18]}
   );
   gpc1_1 gpc1359 (
      {stage2_6[33]},
      {stage3_6[19]}
   );
   gpc1_1 gpc1360 (
      {stage2_6[34]},
      {stage3_6[20]}
   );
   gpc1_1 gpc1361 (
      {stage2_6[35]},
      {stage3_6[21]}
   );
   gpc1_1 gpc1362 (
      {stage2_6[36]},
      {stage3_6[22]}
   );
   gpc1_1 gpc1363 (
      {stage2_6[37]},
      {stage3_6[23]}
   );
   gpc1_1 gpc1364 (
      {stage2_6[38]},
      {stage3_6[24]}
   );
   gpc1_1 gpc1365 (
      {stage2_6[39]},
      {stage3_6[25]}
   );
   gpc1_1 gpc1366 (
      {stage2_6[40]},
      {stage3_6[26]}
   );
   gpc1_1 gpc1367 (
      {stage2_6[41]},
      {stage3_6[27]}
   );
   gpc1_1 gpc1368 (
      {stage2_6[42]},
      {stage3_6[28]}
   );
   gpc1_1 gpc1369 (
      {stage2_6[43]},
      {stage3_6[29]}
   );
   gpc1_1 gpc1370 (
      {stage2_6[44]},
      {stage3_6[30]}
   );
   gpc1_1 gpc1371 (
      {stage2_6[45]},
      {stage3_6[31]}
   );
   gpc1_1 gpc1372 (
      {stage2_6[46]},
      {stage3_6[32]}
   );
   gpc1_1 gpc1373 (
      {stage2_6[47]},
      {stage3_6[33]}
   );
   gpc1_1 gpc1374 (
      {stage2_8[33]},
      {stage3_8[11]}
   );
   gpc1_1 gpc1375 (
      {stage2_8[34]},
      {stage3_8[12]}
   );
   gpc1_1 gpc1376 (
      {stage2_8[35]},
      {stage3_8[13]}
   );
   gpc1_1 gpc1377 (
      {stage2_8[36]},
      {stage3_8[14]}
   );
   gpc1_1 gpc1378 (
      {stage2_8[37]},
      {stage3_8[15]}
   );
   gpc1_1 gpc1379 (
      {stage2_8[38]},
      {stage3_8[16]}
   );
   gpc1_1 gpc1380 (
      {stage2_10[18]},
      {stage3_10[9]}
   );
   gpc1_1 gpc1381 (
      {stage2_10[19]},
      {stage3_10[10]}
   );
   gpc1_1 gpc1382 (
      {stage2_10[20]},
      {stage3_10[11]}
   );
   gpc1_1 gpc1383 (
      {stage2_10[21]},
      {stage3_10[12]}
   );
   gpc1_1 gpc1384 (
      {stage2_11[25]},
      {stage3_11[12]}
   );
   gpc1_1 gpc1385 (
      {stage2_11[26]},
      {stage3_11[13]}
   );
   gpc1_1 gpc1386 (
      {stage2_12[11]},
      {stage3_12[9]}
   );
   gpc1_1 gpc1387 (
      {stage2_12[12]},
      {stage3_12[10]}
   );
   gpc1_1 gpc1388 (
      {stage2_12[13]},
      {stage3_12[11]}
   );
   gpc1_1 gpc1389 (
      {stage2_12[14]},
      {stage3_12[12]}
   );
   gpc1_1 gpc1390 (
      {stage2_12[15]},
      {stage3_12[13]}
   );
   gpc1_1 gpc1391 (
      {stage2_12[16]},
      {stage3_12[14]}
   );
   gpc1_1 gpc1392 (
      {stage2_12[17]},
      {stage3_12[15]}
   );
   gpc1_1 gpc1393 (
      {stage2_12[18]},
      {stage3_12[16]}
   );
   gpc1_1 gpc1394 (
      {stage2_12[19]},
      {stage3_12[17]}
   );
   gpc1_1 gpc1395 (
      {stage2_12[20]},
      {stage3_12[18]}
   );
   gpc1_1 gpc1396 (
      {stage2_13[30]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1397 (
      {stage2_13[31]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1398 (
      {stage2_13[32]},
      {stage3_13[8]}
   );
   gpc1_1 gpc1399 (
      {stage2_13[33]},
      {stage3_13[9]}
   );
   gpc1_1 gpc1400 (
      {stage2_13[34]},
      {stage3_13[10]}
   );
   gpc1_1 gpc1401 (
      {stage2_14[12]},
      {stage3_14[7]}
   );
   gpc1_1 gpc1402 (
      {stage2_14[13]},
      {stage3_14[8]}
   );
   gpc1_1 gpc1403 (
      {stage2_14[14]},
      {stage3_14[9]}
   );
   gpc1_1 gpc1404 (
      {stage2_14[15]},
      {stage3_14[10]}
   );
   gpc1_1 gpc1405 (
      {stage2_14[16]},
      {stage3_14[11]}
   );
   gpc1_1 gpc1406 (
      {stage2_14[17]},
      {stage3_14[12]}
   );
   gpc1_1 gpc1407 (
      {stage2_14[18]},
      {stage3_14[13]}
   );
   gpc1_1 gpc1408 (
      {stage2_14[19]},
      {stage3_14[14]}
   );
   gpc1_1 gpc1409 (
      {stage2_14[20]},
      {stage3_14[15]}
   );
   gpc1_1 gpc1410 (
      {stage2_14[21]},
      {stage3_14[16]}
   );
   gpc1_1 gpc1411 (
      {stage2_14[22]},
      {stage3_14[17]}
   );
   gpc1_1 gpc1412 (
      {stage2_14[23]},
      {stage3_14[18]}
   );
   gpc1_1 gpc1413 (
      {stage2_14[24]},
      {stage3_14[19]}
   );
   gpc1_1 gpc1414 (
      {stage2_14[25]},
      {stage3_14[20]}
   );
   gpc1_1 gpc1415 (
      {stage2_14[26]},
      {stage3_14[21]}
   );
   gpc1_1 gpc1416 (
      {stage2_16[18]},
      {stage3_16[8]}
   );
   gpc1_1 gpc1417 (
      {stage2_16[19]},
      {stage3_16[9]}
   );
   gpc1_1 gpc1418 (
      {stage2_16[20]},
      {stage3_16[10]}
   );
   gpc1_1 gpc1419 (
      {stage2_16[21]},
      {stage3_16[11]}
   );
   gpc1_1 gpc1420 (
      {stage2_16[22]},
      {stage3_16[12]}
   );
   gpc1_1 gpc1421 (
      {stage2_17[31]},
      {stage3_17[7]}
   );
   gpc1_1 gpc1422 (
      {stage2_17[32]},
      {stage3_17[8]}
   );
   gpc1_1 gpc1423 (
      {stage2_17[33]},
      {stage3_17[9]}
   );
   gpc1_1 gpc1424 (
      {stage2_17[34]},
      {stage3_17[10]}
   );
   gpc1_1 gpc1425 (
      {stage2_17[35]},
      {stage3_17[11]}
   );
   gpc1_1 gpc1426 (
      {stage2_17[36]},
      {stage3_17[12]}
   );
   gpc1_1 gpc1427 (
      {stage2_17[37]},
      {stage3_17[13]}
   );
   gpc1_1 gpc1428 (
      {stage2_17[38]},
      {stage3_17[14]}
   );
   gpc1_1 gpc1429 (
      {stage2_17[39]},
      {stage3_17[15]}
   );
   gpc1_1 gpc1430 (
      {stage2_17[40]},
      {stage3_17[16]}
   );
   gpc1_1 gpc1431 (
      {stage2_17[41]},
      {stage3_17[17]}
   );
   gpc1_1 gpc1432 (
      {stage2_17[42]},
      {stage3_17[18]}
   );
   gpc1_1 gpc1433 (
      {stage2_17[43]},
      {stage3_17[19]}
   );
   gpc1_1 gpc1434 (
      {stage2_17[44]},
      {stage3_17[20]}
   );
   gpc1_1 gpc1435 (
      {stage2_17[45]},
      {stage3_17[21]}
   );
   gpc1_1 gpc1436 (
      {stage2_17[46]},
      {stage3_17[22]}
   );
   gpc1_1 gpc1437 (
      {stage2_17[47]},
      {stage3_17[23]}
   );
   gpc1_1 gpc1438 (
      {stage2_17[48]},
      {stage3_17[24]}
   );
   gpc1_1 gpc1439 (
      {stage2_19[9]},
      {stage3_19[14]}
   );
   gpc1_1 gpc1440 (
      {stage2_19[10]},
      {stage3_19[15]}
   );
   gpc1_1 gpc1441 (
      {stage2_19[11]},
      {stage3_19[16]}
   );
   gpc1_1 gpc1442 (
      {stage2_19[12]},
      {stage3_19[17]}
   );
   gpc1_1 gpc1443 (
      {stage2_19[13]},
      {stage3_19[18]}
   );
   gpc1_1 gpc1444 (
      {stage2_19[14]},
      {stage3_19[19]}
   );
   gpc1_1 gpc1445 (
      {stage2_19[15]},
      {stage3_19[20]}
   );
   gpc1_1 gpc1446 (
      {stage2_19[16]},
      {stage3_19[21]}
   );
   gpc1_1 gpc1447 (
      {stage2_19[17]},
      {stage3_19[22]}
   );
   gpc1_1 gpc1448 (
      {stage2_19[18]},
      {stage3_19[23]}
   );
   gpc1_1 gpc1449 (
      {stage2_19[19]},
      {stage3_19[24]}
   );
   gpc1_1 gpc1450 (
      {stage2_19[20]},
      {stage3_19[25]}
   );
   gpc1_1 gpc1451 (
      {stage2_20[49]},
      {stage3_20[9]}
   );
   gpc1_1 gpc1452 (
      {stage2_20[50]},
      {stage3_20[10]}
   );
   gpc1_1 gpc1453 (
      {stage2_20[51]},
      {stage3_20[11]}
   );
   gpc1_1 gpc1454 (
      {stage2_20[52]},
      {stage3_20[12]}
   );
   gpc1_1 gpc1455 (
      {stage2_20[53]},
      {stage3_20[13]}
   );
   gpc1_1 gpc1456 (
      {stage2_20[54]},
      {stage3_20[14]}
   );
   gpc1_1 gpc1457 (
      {stage2_20[55]},
      {stage3_20[15]}
   );
   gpc1_1 gpc1458 (
      {stage2_21[18]},
      {stage3_21[11]}
   );
   gpc1_1 gpc1459 (
      {stage2_21[19]},
      {stage3_21[12]}
   );
   gpc1_1 gpc1460 (
      {stage2_21[20]},
      {stage3_21[13]}
   );
   gpc1_1 gpc1461 (
      {stage2_22[26]},
      {stage3_22[15]}
   );
   gpc1_1 gpc1462 (
      {stage2_24[24]},
      {stage3_24[10]}
   );
   gpc1_1 gpc1463 (
      {stage2_24[25]},
      {stage3_24[11]}
   );
   gpc1_1 gpc1464 (
      {stage2_24[26]},
      {stage3_24[12]}
   );
   gpc1_1 gpc1465 (
      {stage2_24[27]},
      {stage3_24[13]}
   );
   gpc1_1 gpc1466 (
      {stage2_24[28]},
      {stage3_24[14]}
   );
   gpc1_1 gpc1467 (
      {stage2_24[29]},
      {stage3_24[15]}
   );
   gpc1_1 gpc1468 (
      {stage2_24[30]},
      {stage3_24[16]}
   );
   gpc1_1 gpc1469 (
      {stage2_24[31]},
      {stage3_24[17]}
   );
   gpc1_1 gpc1470 (
      {stage2_24[32]},
      {stage3_24[18]}
   );
   gpc1_1 gpc1471 (
      {stage2_26[36]},
      {stage3_26[18]}
   );
   gpc1_1 gpc1472 (
      {stage2_29[30]},
      {stage3_29[16]}
   );
   gpc1_1 gpc1473 (
      {stage2_29[31]},
      {stage3_29[17]}
   );
   gpc1_1 gpc1474 (
      {stage2_30[18]},
      {stage3_30[14]}
   );
   gpc1_1 gpc1475 (
      {stage2_32[24]},
      {stage3_32[10]}
   );
   gpc1_1 gpc1476 (
      {stage2_32[25]},
      {stage3_32[11]}
   );
   gpc1_1 gpc1477 (
      {stage2_32[26]},
      {stage3_32[12]}
   );
   gpc1_1 gpc1478 (
      {stage2_32[27]},
      {stage3_32[13]}
   );
   gpc1_1 gpc1479 (
      {stage2_32[28]},
      {stage3_32[14]}
   );
   gpc1_1 gpc1480 (
      {stage2_33[7]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1481 (
      {stage2_33[8]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1482 (
      {stage2_33[9]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1483 (
      {stage2_33[10]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1484 (
      {stage2_33[11]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1485 (
      {stage2_33[12]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1486 (
      {stage2_33[13]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1487 (
      {stage2_33[14]},
      {stage3_33[17]}
   );
   gpc1_1 gpc1488 (
      {stage2_33[15]},
      {stage3_33[18]}
   );
   gpc1_1 gpc1489 (
      {stage2_33[16]},
      {stage3_33[19]}
   );
   gpc1_1 gpc1490 (
      {stage2_33[17]},
      {stage3_33[20]}
   );
   gpc1_1 gpc1491 (
      {stage2_34[2]},
      {stage3_34[5]}
   );
   gpc1_1 gpc1492 (
      {stage2_34[3]},
      {stage3_34[6]}
   );
   gpc1_1 gpc1493 (
      {stage2_34[4]},
      {stage3_34[7]}
   );
   gpc1_1 gpc1494 (
      {stage2_34[5]},
      {stage3_34[8]}
   );
   gpc606_5 gpc1495 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc207_4 gpc1496 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6]},
      {stage3_3[0], stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc117_4 gpc1497 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8]},
      {stage3_4[0]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc1498 (
      {stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[1]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[3]}
   );
   gpc615_5 gpc1499 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[2]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[4]}
   );
   gpc615_5 gpc1500 (
      {stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15]},
      {stage3_5[3]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[5]}
   );
   gpc1343_5 gpc1501 (
      {stage3_6[18], stage3_6[19], stage3_6[20]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2]},
      {stage3_9[0]},
      {stage4_10[0],stage4_9[0],stage4_8[3],stage4_7[3],stage4_6[4]}
   );
   gpc1343_5 gpc1502 (
      {stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_9[1]},
      {stage4_10[1],stage4_9[1],stage4_8[4],stage4_7[4],stage4_6[5]}
   );
   gpc606_5 gpc1503 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[2],stage4_9[2],stage4_8[5],stage4_7[5],stage4_6[6]}
   );
   gpc1343_5 gpc1504 (
      {stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[3]}
   );
   gpc1343_5 gpc1505 (
      {stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[1]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[4]}
   );
   gpc1343_5 gpc1506 (
      {stage3_9[8], 1'b0, 1'b0},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_11[6], stage3_11[7], stage3_11[8]},
      {stage3_12[2]},
      {stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[5]}
   );
   gpc615_5 gpc1507 (
      {stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12], stage3_11[13]},
      {stage3_12[3]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc1508 (
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc1509 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[2],stage4_14[2],stage4_13[5],stage4_12[5]}
   );
   gpc207_4 gpc1510 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], 1'b0, 1'b0},
      {stage3_15[0], stage3_15[1]},
      {stage4_16[2],stage4_15[3],stage4_14[3],stage4_13[6]}
   );
   gpc615_5 gpc1511 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[2]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[0],stage4_16[3],stage4_15[4],stage4_14[4]}
   );
   gpc615_5 gpc1512 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21]},
      {stage3_15[3]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[1],stage4_16[4],stage4_15[5],stage4_14[5]}
   );
   gpc606_5 gpc1513 (
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[2],stage4_17[2],stage4_16[5],stage4_15[6]}
   );
   gpc606_5 gpc1514 (
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[3],stage4_17[3]}
   );
   gpc606_5 gpc1515 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[2],stage4_18[4],stage4_17[4]}
   );
   gpc606_5 gpc1516 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage4_21[2],stage4_20[2],stage4_19[3],stage4_18[5],stage4_17[5]}
   );
   gpc615_5 gpc1517 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4]},
      {stage3_19[18]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[3],stage4_20[3],stage4_19[4],stage4_18[6]}
   );
   gpc615_5 gpc1518 (
      {stage3_18[5], stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9]},
      {stage3_19[19]},
      {stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11]},
      {stage4_22[1],stage4_21[4],stage4_20[4],stage4_19[5],stage4_18[7]}
   );
   gpc615_5 gpc1519 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24]},
      {stage3_20[12]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[2],stage4_21[5],stage4_20[5],stage4_19[6]}
   );
   gpc606_5 gpc1520 (
      {stage3_20[13], stage3_20[14], stage3_20[15], 1'b0, 1'b0, 1'b0},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[3],stage4_21[6],stage4_20[6]}
   );
   gpc606_5 gpc1521 (
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[1],stage4_23[2],stage4_22[4],stage4_21[7]}
   );
   gpc615_5 gpc1522 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[6]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[1],stage4_24[2],stage4_23[3],stage4_22[5]}
   );
   gpc615_5 gpc1523 (
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15]},
      {stage3_23[7]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[2],stage4_24[3],stage4_23[4],stage4_22[6]}
   );
   gpc615_5 gpc1524 (
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[2],stage4_25[3]}
   );
   gpc1325_5 gpc1525 (
      {stage3_25[5], stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9]},
      {stage3_26[1], stage3_26[2]},
      {stage3_27[6], stage3_27[7], stage3_27[8]},
      {stage3_28[0]},
      {stage4_29[1],stage4_28[1],stage4_27[1],stage4_26[3],stage4_25[4]}
   );
   gpc1325_5 gpc1526 (
      {stage3_25[10], stage3_25[11], stage3_25[12], stage3_25[13], 1'b0},
      {stage3_26[3], stage3_26[4]},
      {stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage3_28[1]},
      {stage4_29[2],stage4_28[2],stage4_27[2],stage4_26[4],stage4_25[5]}
   );
   gpc7_3 gpc1527 (
      {stage3_26[5], stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[3],stage4_27[3],stage4_26[5]}
   );
   gpc1163_5 gpc1528 (
      {stage3_28[2], stage3_28[3], stage3_28[4]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[0]},
      {stage3_31[0]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[3],stage4_28[4]}
   );
   gpc1163_5 gpc1529 (
      {stage3_28[5], stage3_28[6], stage3_28[7]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_30[1]},
      {stage3_31[1]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[4],stage4_28[5]}
   );
   gpc1163_5 gpc1530 (
      {stage3_28[8], stage3_28[9], stage3_28[10]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_30[2]},
      {stage3_31[2]},
      {stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[5],stage4_28[6]}
   );
   gpc606_5 gpc1531 (
      {stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7], stage3_30[8]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[0],stage4_32[3],stage4_31[3],stage4_30[3]}
   );
   gpc606_5 gpc1532 (
      {stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13], stage3_30[14]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[1],stage4_32[4],stage4_31[4],stage4_30[4]}
   );
   gpc606_5 gpc1533 (
      {stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[2],stage4_32[5],stage4_31[5]}
   );
   gpc1163_5 gpc1534 (
      {stage3_32[12], stage3_32[13], stage3_32[14]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_34[0]},
      {stage3_35[0]},
      {stage4_36[0],stage4_35[1],stage4_34[3],stage4_33[3],stage4_32[6]}
   );
   gpc1_1 gpc1535 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1536 (
      {stage3_1[7]},
      {stage4_1[2]}
   );
   gpc1_1 gpc1537 (
      {stage3_1[8]},
      {stage4_1[3]}
   );
   gpc1_1 gpc1538 (
      {stage3_1[9]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1539 (
      {stage3_1[10]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1540 (
      {stage3_1[11]},
      {stage4_1[6]}
   );
   gpc1_1 gpc1541 (
      {stage3_1[12]},
      {stage4_1[7]}
   );
   gpc1_1 gpc1542 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1543 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc1544 (
      {stage3_3[9]},
      {stage4_3[3]}
   );
   gpc1_1 gpc1545 (
      {stage3_3[10]},
      {stage4_3[4]}
   );
   gpc1_1 gpc1546 (
      {stage3_3[11]},
      {stage4_3[5]}
   );
   gpc1_1 gpc1547 (
      {stage3_3[12]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1548 (
      {stage3_4[16]},
      {stage4_4[6]}
   );
   gpc1_1 gpc1549 (
      {stage3_4[17]},
      {stage4_4[7]}
   );
   gpc1_1 gpc1550 (
      {stage3_5[4]},
      {stage4_5[4]}
   );
   gpc1_1 gpc1551 (
      {stage3_5[5]},
      {stage4_5[5]}
   );
   gpc1_1 gpc1552 (
      {stage3_5[6]},
      {stage4_5[6]}
   );
   gpc1_1 gpc1553 (
      {stage3_5[7]},
      {stage4_5[7]}
   );
   gpc1_1 gpc1554 (
      {stage3_5[8]},
      {stage4_5[8]}
   );
   gpc1_1 gpc1555 (
      {stage3_6[30]},
      {stage4_6[7]}
   );
   gpc1_1 gpc1556 (
      {stage3_6[31]},
      {stage4_6[8]}
   );
   gpc1_1 gpc1557 (
      {stage3_6[32]},
      {stage4_6[9]}
   );
   gpc1_1 gpc1558 (
      {stage3_6[33]},
      {stage4_6[10]}
   );
   gpc1_1 gpc1559 (
      {stage3_7[8]},
      {stage4_7[6]}
   );
   gpc1_1 gpc1560 (
      {stage3_7[9]},
      {stage4_7[7]}
   );
   gpc1_1 gpc1561 (
      {stage3_7[10]},
      {stage4_7[8]}
   );
   gpc1_1 gpc1562 (
      {stage3_7[11]},
      {stage4_7[9]}
   );
   gpc1_1 gpc1563 (
      {stage3_7[12]},
      {stage4_7[10]}
   );
   gpc1_1 gpc1564 (
      {stage3_8[12]},
      {stage4_8[6]}
   );
   gpc1_1 gpc1565 (
      {stage3_8[13]},
      {stage4_8[7]}
   );
   gpc1_1 gpc1566 (
      {stage3_8[14]},
      {stage4_8[8]}
   );
   gpc1_1 gpc1567 (
      {stage3_8[15]},
      {stage4_8[9]}
   );
   gpc1_1 gpc1568 (
      {stage3_8[16]},
      {stage4_8[10]}
   );
   gpc1_1 gpc1569 (
      {stage3_10[12]},
      {stage4_10[6]}
   );
   gpc1_1 gpc1570 (
      {stage3_12[16]},
      {stage4_12[6]}
   );
   gpc1_1 gpc1571 (
      {stage3_12[17]},
      {stage4_12[7]}
   );
   gpc1_1 gpc1572 (
      {stage3_12[18]},
      {stage4_12[8]}
   );
   gpc1_1 gpc1573 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc1574 (
      {stage3_15[11]},
      {stage4_15[8]}
   );
   gpc1_1 gpc1575 (
      {stage3_16[12]},
      {stage4_16[6]}
   );
   gpc1_1 gpc1576 (
      {stage3_17[24]},
      {stage4_17[6]}
   );
   gpc1_1 gpc1577 (
      {stage3_18[10]},
      {stage4_18[8]}
   );
   gpc1_1 gpc1578 (
      {stage3_18[11]},
      {stage4_18[9]}
   );
   gpc1_1 gpc1579 (
      {stage3_18[12]},
      {stage4_18[10]}
   );
   gpc1_1 gpc1580 (
      {stage3_18[13]},
      {stage4_18[11]}
   );
   gpc1_1 gpc1581 (
      {stage3_19[25]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1582 (
      {stage3_21[12]},
      {stage4_21[8]}
   );
   gpc1_1 gpc1583 (
      {stage3_21[13]},
      {stage4_21[9]}
   );
   gpc1_1 gpc1584 (
      {stage3_23[8]},
      {stage4_23[5]}
   );
   gpc1_1 gpc1585 (
      {stage3_23[9]},
      {stage4_23[6]}
   );
   gpc1_1 gpc1586 (
      {stage3_23[10]},
      {stage4_23[7]}
   );
   gpc1_1 gpc1587 (
      {stage3_24[12]},
      {stage4_24[4]}
   );
   gpc1_1 gpc1588 (
      {stage3_24[13]},
      {stage4_24[5]}
   );
   gpc1_1 gpc1589 (
      {stage3_24[14]},
      {stage4_24[6]}
   );
   gpc1_1 gpc1590 (
      {stage3_24[15]},
      {stage4_24[7]}
   );
   gpc1_1 gpc1591 (
      {stage3_24[16]},
      {stage4_24[8]}
   );
   gpc1_1 gpc1592 (
      {stage3_24[17]},
      {stage4_24[9]}
   );
   gpc1_1 gpc1593 (
      {stage3_24[18]},
      {stage4_24[10]}
   );
   gpc1_1 gpc1594 (
      {stage3_26[12]},
      {stage4_26[6]}
   );
   gpc1_1 gpc1595 (
      {stage3_26[13]},
      {stage4_26[7]}
   );
   gpc1_1 gpc1596 (
      {stage3_26[14]},
      {stage4_26[8]}
   );
   gpc1_1 gpc1597 (
      {stage3_26[15]},
      {stage4_26[9]}
   );
   gpc1_1 gpc1598 (
      {stage3_26[16]},
      {stage4_26[10]}
   );
   gpc1_1 gpc1599 (
      {stage3_26[17]},
      {stage4_26[11]}
   );
   gpc1_1 gpc1600 (
      {stage3_26[18]},
      {stage4_26[12]}
   );
   gpc1_1 gpc1601 (
      {stage3_27[12]},
      {stage4_27[4]}
   );
   gpc1_1 gpc1602 (
      {stage3_27[13]},
      {stage4_27[5]}
   );
   gpc1_1 gpc1603 (
      {stage3_33[12]},
      {stage4_33[4]}
   );
   gpc1_1 gpc1604 (
      {stage3_33[13]},
      {stage4_33[5]}
   );
   gpc1_1 gpc1605 (
      {stage3_33[14]},
      {stage4_33[6]}
   );
   gpc1_1 gpc1606 (
      {stage3_33[15]},
      {stage4_33[7]}
   );
   gpc1_1 gpc1607 (
      {stage3_33[16]},
      {stage4_33[8]}
   );
   gpc1_1 gpc1608 (
      {stage3_33[17]},
      {stage4_33[9]}
   );
   gpc1_1 gpc1609 (
      {stage3_33[18]},
      {stage4_33[10]}
   );
   gpc1_1 gpc1610 (
      {stage3_33[19]},
      {stage4_33[11]}
   );
   gpc1_1 gpc1611 (
      {stage3_33[20]},
      {stage4_33[12]}
   );
   gpc1_1 gpc1612 (
      {stage3_34[1]},
      {stage4_34[4]}
   );
   gpc1_1 gpc1613 (
      {stage3_34[2]},
      {stage4_34[5]}
   );
   gpc1_1 gpc1614 (
      {stage3_34[3]},
      {stage4_34[6]}
   );
   gpc1_1 gpc1615 (
      {stage3_34[4]},
      {stage4_34[7]}
   );
   gpc1_1 gpc1616 (
      {stage3_34[5]},
      {stage4_34[8]}
   );
   gpc1_1 gpc1617 (
      {stage3_34[6]},
      {stage4_34[9]}
   );
   gpc1_1 gpc1618 (
      {stage3_34[7]},
      {stage4_34[10]}
   );
   gpc1_1 gpc1619 (
      {stage3_34[8]},
      {stage4_34[11]}
   );
   gpc1_1 gpc1620 (
      {stage3_35[1]},
      {stage4_35[2]}
   );
   gpc1_1 gpc1621 (
      {stage3_36[0]},
      {stage4_36[1]}
   );
   gpc207_4 gpc1622 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1325_5 gpc1623 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], 1'b0},
      {stage4_3[2], stage4_3[3]},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc615_5 gpc1624 (
      {stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6], stage4_4[7]},
      {stage4_5[1]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[2]}
   );
   gpc606_5 gpc1625 (
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2]}
   );
   gpc606_5 gpc1626 (
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], 1'b0},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[3]}
   );
   gpc615_5 gpc1627 (
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10]},
      {stage4_8[6]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[1],stage5_9[2],stage5_8[3],stage5_7[3]}
   );
   gpc207_4 gpc1628 (
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[2]}
   );
   gpc606_5 gpc1629 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1]}
   );
   gpc7_3 gpc1630 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage5_15[1],stage5_14[1],stage5_13[2]}
   );
   gpc615_5 gpc1631 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[2]}
   );
   gpc606_5 gpc1632 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[1],stage5_18[1],stage5_17[1],stage5_16[2]}
   );
   gpc615_5 gpc1633 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[2]}
   );
   gpc615_5 gpc1634 (
      {stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage4_20[6]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[1],stage5_21[1],stage5_20[2],stage5_19[3]}
   );
   gpc207_4 gpc1635 (
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[0],stage5_23[1],stage5_22[2]}
   );
   gpc615_5 gpc1636 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4]},
      {stage4_24[2]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1],stage5_23[2]}
   );
   gpc606_5 gpc1637 (
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[2],stage5_24[2]}
   );
   gpc606_5 gpc1638 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[2]}
   );
   gpc606_5 gpc1639 (
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[3]}
   );
   gpc606_5 gpc1640 (
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[0],stage5_31[1]}
   );
   gpc606_5 gpc1641 (
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[1],stage5_34[1],stage5_33[1],stage5_32[1]}
   );
   gpc606_5 gpc1642 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[0], stage4_35[1], stage4_35[2], 1'b0, 1'b0, 1'b0},
      {stage5_37[0],stage5_36[1],stage5_35[2],stage5_34[2],stage5_33[2]}
   );
   gpc1406_5 gpc1643 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage4_36[0], stage4_36[1], 1'b0, 1'b0},
      {1'b0},
      {stage5_38[0],stage5_37[1],stage5_36[2],stage5_35[3],stage5_34[3]}
   );
   gpc1_1 gpc1644 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1645 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1646 (
      {stage4_1[7]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1647 (
      {stage4_3[4]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1648 (
      {stage4_3[5]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1649 (
      {stage4_3[6]},
      {stage5_3[4]}
   );
   gpc1_1 gpc1650 (
      {stage4_5[8]},
      {stage5_5[3]}
   );
   gpc1_1 gpc1651 (
      {stage4_8[7]},
      {stage5_8[4]}
   );
   gpc1_1 gpc1652 (
      {stage4_8[8]},
      {stage5_8[5]}
   );
   gpc1_1 gpc1653 (
      {stage4_8[9]},
      {stage5_8[6]}
   );
   gpc1_1 gpc1654 (
      {stage4_8[10]},
      {stage5_8[7]}
   );
   gpc1_1 gpc1655 (
      {stage4_11[0]},
      {stage5_11[2]}
   );
   gpc1_1 gpc1656 (
      {stage4_11[1]},
      {stage5_11[3]}
   );
   gpc1_1 gpc1657 (
      {stage4_11[2]},
      {stage5_11[4]}
   );
   gpc1_1 gpc1658 (
      {stage4_11[3]},
      {stage5_11[5]}
   );
   gpc1_1 gpc1659 (
      {stage4_12[8]},
      {stage5_12[2]}
   );
   gpc1_1 gpc1660 (
      {stage4_15[5]},
      {stage5_15[3]}
   );
   gpc1_1 gpc1661 (
      {stage4_15[6]},
      {stage5_15[4]}
   );
   gpc1_1 gpc1662 (
      {stage4_15[7]},
      {stage5_15[5]}
   );
   gpc1_1 gpc1663 (
      {stage4_15[8]},
      {stage5_15[6]}
   );
   gpc1_1 gpc1664 (
      {stage4_17[6]},
      {stage5_17[2]}
   );
   gpc1_1 gpc1665 (
      {stage4_18[11]},
      {stage5_18[3]}
   );
   gpc1_1 gpc1666 (
      {stage4_19[6]},
      {stage5_19[4]}
   );
   gpc1_1 gpc1667 (
      {stage4_19[7]},
      {stage5_19[5]}
   );
   gpc1_1 gpc1668 (
      {stage4_21[6]},
      {stage5_21[2]}
   );
   gpc1_1 gpc1669 (
      {stage4_21[7]},
      {stage5_21[3]}
   );
   gpc1_1 gpc1670 (
      {stage4_21[8]},
      {stage5_21[4]}
   );
   gpc1_1 gpc1671 (
      {stage4_21[9]},
      {stage5_21[5]}
   );
   gpc1_1 gpc1672 (
      {stage4_23[5]},
      {stage5_23[3]}
   );
   gpc1_1 gpc1673 (
      {stage4_23[6]},
      {stage5_23[4]}
   );
   gpc1_1 gpc1674 (
      {stage4_23[7]},
      {stage5_23[5]}
   );
   gpc1_1 gpc1675 (
      {stage4_24[9]},
      {stage5_24[3]}
   );
   gpc1_1 gpc1676 (
      {stage4_24[10]},
      {stage5_24[4]}
   );
   gpc1_1 gpc1677 (
      {stage4_26[12]},
      {stage5_26[3]}
   );
   gpc1_1 gpc1678 (
      {stage4_28[6]},
      {stage5_28[3]}
   );
   gpc1_1 gpc1679 (
      {stage4_30[0]},
      {stage5_30[2]}
   );
   gpc1_1 gpc1680 (
      {stage4_30[1]},
      {stage5_30[3]}
   );
   gpc1_1 gpc1681 (
      {stage4_30[2]},
      {stage5_30[4]}
   );
   gpc1_1 gpc1682 (
      {stage4_30[3]},
      {stage5_30[5]}
   );
   gpc1_1 gpc1683 (
      {stage4_30[4]},
      {stage5_30[6]}
   );
   gpc1_1 gpc1684 (
      {stage4_32[6]},
      {stage5_32[2]}
   );
   gpc1_1 gpc1685 (
      {stage4_33[12]},
      {stage5_33[3]}
   );
   gpc1325_5 gpc1686 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0], stage5_4[1]},
      {stage5_5[0], stage5_5[1], stage5_5[2]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc1343_5 gpc1687 (
      {stage5_6[1], stage5_6[2], stage5_6[3]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3]},
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1325_5 gpc1688 (
      {stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7]},
      {stage5_9[1], stage5_9[2]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[1]}
   );
   gpc135_4 gpc1689 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc623_5 gpc1690 (
      {stage5_13[1], stage5_13[2], 1'b0},
      {stage5_14[0], stage5_14[1]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc1691 (
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0], stage5_17[1], stage5_17[2], 1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2]},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1]}
   );
   gpc2135_5 gpc1692 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[1]}
   );
   gpc615_5 gpc1693 (
      {stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage5_22[2]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage6_25[0],stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[1]}
   );
   gpc135_4 gpc1694 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4]},
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[1],stage6_24[1]}
   );
   gpc1343_5 gpc1695 (
      {stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[1]}
   );
   gpc7_3 gpc1696 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage6_32[0],stage6_31[0],stage6_30[1]}
   );
   gpc1343_5 gpc1697 (
      {stage5_31[0], stage5_31[1], 1'b0},
      {stage5_32[0], stage5_32[1], stage5_32[2], 1'b0},
      {stage5_33[0], stage5_33[1], stage5_33[2]},
      {stage5_34[0]},
      {stage6_35[0],stage6_34[0],stage6_33[0],stage6_32[1],stage6_31[1]}
   );
   gpc1343_5 gpc1698 (
      {stage5_34[1], stage5_34[2], stage5_34[3]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3]},
      {stage5_36[0], stage5_36[1], stage5_36[2]},
      {stage5_37[0]},
      {stage6_38[0],stage6_37[0],stage6_36[0],stage6_35[1],stage6_34[1]}
   );
   gpc1_1 gpc1699 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc1700 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc1701 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc1702 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1703 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc1704 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1705 (
      {stage5_4[2]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1706 (
      {stage5_5[3]},
      {stage6_5[1]}
   );
   gpc1_1 gpc1707 (
      {stage5_15[6]},
      {stage6_15[1]}
   );
   gpc1_1 gpc1708 (
      {stage5_18[3]},
      {stage6_18[1]}
   );
   gpc1_1 gpc1709 (
      {stage5_28[3]},
      {stage6_28[1]}
   );
   gpc1_1 gpc1710 (
      {stage5_29[1]},
      {stage6_29[1]}
   );
   gpc1_1 gpc1711 (
      {stage5_33[3]},
      {stage6_33[1]}
   );
   gpc1_1 gpc1712 (
      {stage5_37[1]},
      {stage6_37[1]}
   );
   gpc1_1 gpc1713 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [38:0] srcsum;
    wire [38:0] dstsum;
    wire test;
    compressor_CLA128_32 compressor_CLA128_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he5c4167438c050291b6b163ca447b2f52b3019b9fc9670a13450099358433a38e5c6fb495de39de5ab60e379ff14c02e64aef95bbb8e856b8443aed2cadcf2b7978f25fc3a062b785d46a93b96e9b6818786b38a8e05435df9aa726acb906e8a118c43dc20dd8f136ee2f2a2ed86a0ba98d19e6b88d77345862206505ea36e8981e12a19a684ecce13c02e57a5f67f945019b1bd737010f82847d9b1b1333b57a0054d5c5ff80327956446fe1e595c97ed76aafe7787258ac091927a3b49c96d1f60cf18fd083cb4961de45b71b8b82f97751e344bde058293aee3ebcc519e9329df523b876b70b4f318302cca37ff8ebb5d1a84bf5a4ae9a17b004e09b8f9f0fd041521b8f958c52ff5a597d9aae7505e7b204cb4582f5edabd4cf7c9776bf12539c73bdb27f46553a770f37c033a40a564c01371e24ae8dbb35fdc72503964e28a3d933ce4c8e44b440abc1858a6f4057d2c454acdb1a53315ae04af062d4ae415707cfd65f91f1f783f02836213acccfe7249bc9b8fa80fb920cd70e012632287e2864a0be93db91798767fd6491d817360fbe240e4dc6d0b87fa21b2d2782b81bcf9b76a8efae7e879e91c9f03e1835e77fda14d8c151db5e08d60e5327231c7d03f982b08314a3a08445c6bad7d373e988a6249657425f68c4e7d9633c9597d8b94723c99cd2567adaa39031c484971d46f6489c176d74d96ac5126dc5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7f5bab994ecc05107b9bed9e66c38f3b1458a358427f943647aa8c1c37eced41c10b50cdedf703b6b1d11815bf844b801de2c95ec961d2b5df7dd16cadb566fbce1961fec9b44a448e2939cc5e8c97d4adc80af1982187044eaf6c67f248e0fcefc0d248f5eff9dc84518c9b50b33c888cdd84d407707e5a468783dd907c29500a425e0d68ff604012194780bb164d71c1e88e5dce20221b27139ea12824497fb21ce962edb70b695b0dc36c6b724a9adb6961a839dddebd0a8f7299d058c0c42a588f81f498d02a2e8d6ec74ae988c1cd07258c52bb8ff47bb4f4cae03586e514640ca7912c2a351c6f6c1d9074c59f5546e2314f9e7c5c31b078acbae8276300926de3d7d6fb5434db7805a662bd23ce4f16fad3473bf8ebfa825af2e3fa0ecfe51fa906776350d842e77cc7c90173462b274f147c441732e82d702ecb143527c3f185050e1c0fb971dc97dc46be254a8c3e0d6ff0d8002f8bbf1043b7369edde70a1d8c83647b9df92e084ae80902d92439f3c0e4cce4550ba71caa025ff7f9bc03f7b5c268dd1df42fd2bee5167bcf46d924fc9f0f1450eb27d8d09897605475944a1a7e8e72449f04faa75b5944749ff30088650eea4e314e9abc56122b253b8705d012b483ac42ac373abdc29913c815b72bcd172dde9fe1098d457ce2b969be9c3bc704050c698cc787e7c2d483d3fbb0cb914de880814b7f559e93fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbc2839c1e522800073af3348594f30b5dc760eccd4d05cb0246e33e8d766001fbffef1b42cbff16e7c463894122ea97d28bdd53b0a13cea3a410afed074e70789b22a28a3a1d5623d9f1fd5522c845f8a929a03ccbb559a78ee37bbf9fc0a643ba9dc41a4321d1a90016516fcf8fa8711651582094701a24f69f92b437d3d9a73ead49161d4fe2f0ccb7959f2907e04ca8b875bb56495e70b391fbe8e27a77bc46220a9c2b9cf7fbd9c0f43697c1a6e32d3db3e4304387490da734b4e4231231019222e6ad82bfe64ae18794479797dcb009f5f563889d0e639c8010de0d1f16e7e194aa4c4099128e60b15582d2b55734105110226fe381557e07be5185c0c06cd4f9fd3dd83a5118d6d6684fd185591b8ae3f4477541746f462c88e97c95a3ffe84f77937c218085d37df43e78805a48c9abd67fd6f3137309ddc7b5bad63fe9cf3f8e2f0c394a5f56a76626bcc78efffe5f7d52900684cade17c2e6ce93c2e3ab30fbfd8ebb9b6a60b1f8c1c17c718497a62223ae1ae3141ce800c9bf6e6dac435a10c4da7e4c555480a02a8bd38bf8139ac93508711adeb3a72fd1f5873e4d718fea920e6b8afa8e228270bc7f2410038c66a990cab4c53c4dbc693cbe2586ec36256662ccdbd886ef86ea769447437fa0e03ad5e8fe6c693b5e97d531ecb77d2d0c27fdb15affe02b0e66f99dc42fe9bfe823a0666aee266b948c35f17b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1c150e39cc2f34f1384f206759d8546c7b5fdd4bcd9277c271b1c15932de69edcf30113f05411bb95005b2413a81f9ee35e89290f9d163fde92f40e60c5944fb35dc4c06442403716633827cc8da1412d62353c2af792d5d071ba29e410476e178acbb2ea6decc76eefb2e1ff94016100ef0856bfe9e73c5f8114d23b0b162c208385aa14d5543c73aba17512f1c5e437b88810e66e512731cb8df6537f3433d4d29aae1c660e76b785742cfeb1c74352306bc2e1bb8793cf29f68fee04a0c181b9f76fe637da347823e2879bb76b39ed8f11bf10d6921eab710a188ca0086cd1410ec90afc4be21138f3a9e6409c0e1d88e7196a88623283e8112e911c070989d069f42cf87f8648dee59b335f21f50eebbdd2784be2625e2dc25bc5653ad426965c3bd3f12edf5b0ffbd855b16ec83ed134d958de24b787aae8983a5d1c59e6accdf4e1adb176363c322da3f6b9f5a92530f478fba9768086dec20790455df3af3a884bc5509934d8ff0d66128fc48976a57786bf8a45f361743b093d9446196830763f73fee0e90f5db6af9b8a5b1b48945e1127dacdde7c979c9b9aa28fb67e44097dac5b3248eba23f6481a5a4e8c8ce418256282d707a23ae6c8e0c76d7f3d2921477ea14c8050a20905c9bb53a8e8dc7fd9e03fd177e0aec7a6cb221e56eaf12762b6a21edefdc1a7c0d3dacae789482d70b21619d0c3474be9a1a743;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h33eab25b6c19468ce19ae054f958dc9bb5a24a4ef70e0817bb8d8e41ef97648618d64d4263ed02cf7c00490b66dee875e7fca26c9c7c087720a9856cd565bc4e2c27664f59f16bcebf71c7e52e4904d0f809271103cb65247cb61057b82f4260d2846705caedc689005be6372f921e8c8ec163b02c1bcaf01b043cf70d3199222dda104e85f2d1e6d04d7c66d14831fc5aa555fd14dbfc8e29768aa7862eeb94d87785b6a6eaa68d943d0db1c98c7cf14cef11fa1347f58f363fb1b1ca93883c107ecbbcee134dff7f790ceceb653ba52653b6e04319eaef8a56882871b2a367787c3f7d4aafca524a9f2aafc12521f411d75cf65fd8c4dec7c4de1003ffdf4096986312894068089670ede1ec16bc754bdaed8949f18b99432b78a3b8c2d7ebc9c324dede55d1672feb12cfd011c0cb53f2c376a8a7fa80b1f9bb51f8d4d3418d6643dc3b938b89f61b4d4686af560847ef4b3ed2c6fcea8128bab55a98d4e43ae152e3a00a291b116d7b4c10be62a6229643a478cac20820715e9505c996d582dff16f09859f753c6d1394cd336397fd790f9219c0ff2a87ad9a24ae73d1fe66032033df5762cfc64581820234a5974650cec22d91b0d16bca26116add1d6e9abfcd1d60831c06bb508ba88a9b290a7bf8c071138db3a4612ec8f6b06c9ad57c1f86682df7993532fd2884c993d4f3ad23d8319a31cba818f0ef5568f7360b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hde5c5f83e89497a2ed19161567c76b216b2bae2b1cd188fa95010ce5e119039048c24908a01416cf89e0dfa32af487648ac06eacb0428f939a63aa729d676bca1fade33608abcb88f979f61d6d2abc0b9b79c6fd41c7261d39195a0cfe6f37c77e3db074855e4c6cbbe9a28014ec9d5dadf0c8c6124db182169608ac43f967b5caf83bdd16d181fb9816161be120e55289862176041e07ce70df2a9863f38dada46bb4c05e0b1f1178b6ceabedb423101ca0dc9145f11b17bdfd9580eafb4d97a9da4fcdb89acfe188faac83420b3d97a747a27c360143fb7248b97e3a53072566b0bd820ef6f0cf087a4367ce576909a6e4432e15a12cee569c67a8a099573b9a050cfedc93879c5abf5a12871182900935999932b0f03137dca1599f5d2bc171b6edddc520e767600bdea2ac9ed9dd8a40b8226d15323ce5a11d04d87ebb49506a7879aa55f6782e003d82480bb403d88042c6b875c391ac85b5848c0ed387484850eb9053f803ceb46fb026d4f536a7ec406bf0dd19793cf4e1b58f0fdb46f726038fc70c2646bd59c22a87079f1de2d708e421ec0831adb5758ba450065a08f838d79038f9489976e69b3d4fe8b529df2b47665e12c026a250428f2dcadc7b9f80d0fd0e30ee75e28ad4baa32544303ef6709e182fcbce8c73ff8c9f984505d4182d2058bbb2fe190f309772a59c0cc7db7ce7b9597deca1816ec1333978;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c6de12dcbd09e06cc25c604b9134e36d1bdee5c40a0febb38a7cdbd84feb7bd926ac6985f7634ff632d6f17b4efdf4aac289695fb95ce985ecb18b52777da2432b9f919ee94550a455c88f094cfc0f45795a8fd570f3c5cab4baac0f3697c22b92a7b68fc5bc210ebb8ce9a7a3ddb1c5bc57cf5fa06964ce8cd9e0867a8e3a802c2aeb6583ad45bb015c4f88a1d0e828445c59350af4473c9ed00e63fcf4dd00ea29e8db0aa17899852b1d8fd8dbf57150488edb5002f0c8ba1420a7c1dccd931089e7d24363a8b533f8e747dff3f4e9ea5322a9cb5f134f61a86766c7a80359698808c8155b4dd5c80abd9cb6f425277af4a92351b277040bb889163a1041e94fc7a135a3869eb0f6d00733b0af6dc0e0eb51422259567d2c36655c90b22f8af430184eef9166639eb7735ebe095c8c5ecb64c52352c593ba22150f163e5adc9393e3dbaa7de6de14d77e87dd18d661f9f74dd7d442139f477ae86562ea1dea3f89f56cce535db2aaa24044845e2e0247a6e84a991b10723677b8f1a8663b424084ef45e0eee55d695f2adf9347a07d8ed4a36c82f9e68e2a7f6b8231abe2baf99c5b8c901cd1cbf5153b244165a5f741f2d3748cccad8f81e6f62d03c9fd80b337033295122c0035caaa23f9dd62f0521379af20bd782a0af5c4d83409d66428d545f1ad039955b2ad7a71395035cd430f1d7c09c40d6495dd983c6acf55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf06d01b8b51b811fb787aebe970117d593c6792d42881ba2596bb7ad88a212ac73b5286f64e4220bf6b046892e3daae47d60fc4a4db539ea7c27f1614c6e43ba1088fb0407d63f55a94f2373a78c47a306f0ab68927b7b3bd9f62f29d255f2b6e66a3097880ee2504224bae4262fbdc7151a2631b66853d16435690c7fc1570285864b2a15a1553d7a5dc858212d612a673f1ed8bf6c8f6cb0981568ecef041efa242990d379955f6292d0db098902cefa35c6e4727344916825735ca94fc0a9d73f55d411c3efac46cb65dbe2bd27755db9c5f83f3ab01393ee7f0978ca3a00f2782ef27166fbd908fc891ccbc93dece7a3ccf12f6559e7d22a9d2416445d6a6e35efc6f1d6a3b8552baf350a4c2d9aa22006ff605e6e1e4850c8d7ee450cebe00ec564282e599959884497ed6d7924a2b858172572a04e9c00463a3ebb8de8ebaa68a21ee7218d6ea4a299b384059602d551ad5c62dab59c456b86da468522c3cbd21ce5ca9bd54382300938f913d756840ccdd7acb3d70b0cea845b14e075ad13a74fd506850aab56d458b3f833c1cbe462962ba6475cda26b1499b2ac8b057ea58fdb06fe43d3c8340019d2b9b31c26d776870799450fd595ca0a38e76bc490c36d152f192d668237a7a489023d11e40a9baef8548c785b8c17bda071bb3405eca1e8100f32992e4b46e37d25d4162d2a2584828226ac939d78e609496e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'haf027f5109feeea8110b693849f15bf128af1ad581527e60b7fd1799ff16f084eee673829e7f39c981e1dca91c71abe0cbef0b7d506eca2014b733ba006723a6ac2632510644f310b1dad737c703ad77749d014b02be1409bbed2e534346718f6b34c58d1dd62e8ba51e2635c8218adfd6f42c9148f98fdf2bbca926fb216e054f5a7b09385344e38d27fa0c9873981908d68e5acb9e7925665b278bec476684b262cbd32ebf60281225bcfd188f3f05ccb89eabdd49499a32c6c779c787eff43ec38808fc0b50b18cc732a9d5fced1b8845f5252c94accdea9a1a27cd38bfcc8fffcc9e9c60cc7ceeb5eeeda6f3411d69286727fa5958caa01b0073964ca7831485ea680917d647e6df64691f3319d24818ed1d0899c485c992a297c8b740e8c43e0385085017a0a9d9ce1b98b30add6d08cc6ff1e2d52df90616e14d203dc55977bc3befdd43092ec6316af216de2f06bfdff6f4474008d3e596bc87232fb0304193c9eb545a4636e9149f8fa543544cbb407542832874cdd5da02dd068953e93313518440da58bed1f8dd2d6fe698a7e3b594f4608e91bb6b03188b3195b33b391a077236432feea46da20ae2245250fd3df9451000aec7eb63bc2c9e714fd92a9a8284c8f921558f947d50e3535a471eb9794f4cd4e17714bef153e1d9954a0e999ff4e2110b482ae219f7bbf315dced2af25774223bfaa6786467fa5c01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc2e5250a63e33aee04a7c6a4961ce5e09ca1cf1a4f7b15a6e9c1763fffaf9d2e8be4e5b53faa774d95e483b76416a82a02e06b7842ff39f00b9202eb62f3ace04cfc4ba025715e90c7c034c6d56bb3bd3617ca6bdc2070bda5ec13d55967c1c6ff7c53eb39cb4a423b2cd64ff87cbe9d3125a1671a536f2ecf8396152c727068bd50e9ae2f77740b8a8e482026d1dd02b82e5b83afb0b30334d5255a4b79d6b457360a332b5b00ae9da55344c51a5fbf95b241f2f2079b38f2a841613fd099b805d6294965cfb781acb7aac74687b305e867487bbb59e51b21f7c01bfd2513ee1d1833379f67d7ef15a80cbfce5b399e04e0db07a2f1359d795d21becf2e0ed4bd56f92874eaf5010ea24978caebd66914278e74f8a6d3e079c1e8b188fee457e84d1b8a5eb75c13ecaf8e9bcff60585457c44610e4100c07fbe9a6da4db5efe17b236a3c4dc7da89cf1cfd37fe63d8ee104522780d9da79c16d1426c0bdfe5b481f87348b18732c1e76d7d602f0d396927be85c7ff2b402ff8c7c6299eb5eadc305fada8ec3eeda63d2b27a1b8c1104394843c71d4a848a5bdfbf8a4c07d6bd55181b733dfbcd1a0a05f8caf2a6a90b093cf841481fb6ac8cafe5d36e2eaf6f598065d027f64da7e3515ffff20ff4b4cda0cc7ca26ea29544e4c4aba2e6fde293c7efdc20fdfb74af52e701f89aa891583ab829afb684bddb588df026cbcac5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5ac7913c1e5b45feb3fd1994300ff9f40f95d3e9111c1ce8f23d0acd30e7829b07caddeace334ce08990b08567d454ecc610f69a36d61f6d9a0e952483a5c71b938cca8a308859021480c2b61f1a8ee0e9905fcf3665653a81845678b839e5d0f29825eb755860536d3b5d8678d84563af0b074b8b53dd41a232b2b09e251e4d2a58b64a6f6ccf13fe22542fb8870947475ec85bfcb6c37c1a7317e06de98985cf09eab0a5185011577769b9a9fc58f5bf9d4572c148f4dbc9bae54f742d158fbb120bf9d1380326fc3ec369bd6f17d3689ada6762431f3f7ca59603feee726437c2a3e83999aff563bc4cee0fd6542f989d0ce3918bca51630bf14954048482c32b7c1e8a03dacd940fbf14fb15681a44ef090a16c1db2053e544b59c64497e5f0b87cbbbb5a81b3e53c9a59d706713c656e9fa0c88619a43ae7defbcb3cffc6819d9c21659922f8f6d61a490f4787caa46cc5619dee91ccbe386ab70d6bb78f78a04607ae2feb0f2e026b058f0e9bd3b56605cb7bb42f24b3d1484e617f4fe232225f85acb3d41070d2d86b658a141e44749f9a1c408e1884f265f7a8e690d86b76e88a0dc3f1fb25924f928bd1234a6ca9d994fc88a0b17f86c965d92128e11e6878563f0e70242aee817026369cbdfc1be0436d7e3da552386b0b91d77789f74d39181163d39402dc938394284660377a6566c22b51eff617a241d4ba655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e50122e76621a79dfca92c0437530fb98974840d89b257e89aec46f8957690b78f1048a3f1e122b76fb249fd79f32e33ceb3839eeee6dc3ffbd8d3565cd2a1f77373dbc97517e098203d4f4887ca60a795e573957e5059a329357a11e1506234d9db8f5825f6c34c4d4c673c84a6f529aed4927eaf6ec2a8c5fd74cf7c927ed9c1fc52108f98d016064b4731eb60cdcc86d453b5583bc37750e845db7e98d66dd4dabe412f5314f79a6710404a3efd1970d9601862a4f3f06b5090c04fc2fc1fee93048f9ccae33b11bbcb9505cced485dd682d19ec474e46a415012c686799e50f6ec3445bdb3b239cb65c19c87e324a6f2e426c8405d0f734bc6c3e8429baca2680bee6ab36f07db8ef03279ae4202a5c4c3fc3baf4300a087023a2f0638ef5fcdc0832dbbd0bbd77c9014239f2023bdc37344b8268b2fce95384bdb21f23d724243227f168b3058116842a0a2894ea6f83b05ae48e95404208d325ebcc95c4e05fd0abbb38a3a62ad5db574a6a08dd1b4673826d681b42299204f2c93ea32bdfb3863ebd7b2fee4fea5910a9861939786a551b48e231ea07006581f65451e7670f05dc184195bebc2aeca07a72da79baa86c1bf1bf3e04af869fe6a69f79904423937ac4528421ef53681d93c2fcdb60facf60d5c55165f35b478c3cbd4a778359f1080bab747d6bf959006650d476f7f55d8d45fc0caacd3784556e0202;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h84b4e43926ed2c72170ac1281a6d7201844ccf94258050ad81a13d9171c8021854e95940711e33f8f1fcfcee30f7bd17310193425d28e074d9575abc34aabc0752276aa70bb160f6c3a17ed19109014ad226442c1d43f094b616d07e05650bc42879bf481765a5252bbb208c65abb513afc3484bbd59f46899c1d3f6ed567e3f6d487ead5aeacc9f48111a0b9e8198cf9f1843a09a85980d3721309adb63adac6b148f273a697f6b6af79eb61e3e535f759857c4af4e40197a7d1872a7e5850402cda773143a819780727eca9065b46d7a21907375f970b73ed38c2168ce309ef040834f35172ee28222aee057568b8c68e79e1376fa1a1cf7e48af222781878c7d9d358a2f6cac43c1e76039ff350a5744ca67d697797f79d4b182c52082f884faa9edd7bf3a1754467ed0ca7ed642d405285eefc3faaa29c43db434f9ccdbde9e0914ad78ab99431aeb08c7a2b6c25a245203eae4fddc10a345b526ca64238abfa7825ce9f610f772a3e98783bd875bce5b1d5f6dfd9355977c8913894acd6dbed3d13b99f681b18b7f082a9473226d51b1c48d877090c07583e0d4cd51a748e6521cc1815745caa51100bf9c2f94c1a3713435141cc8401c34ffefba00d284dd102f87146d4704a1d55fcc21690656a2becf95a7a8c1182070f8ab5c4d1f3a92f379f809cb7319a41f253688eabca3afffd8235fbc4f8a2927e2b9632dab2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4bb74c8f61d272d61ef93e0c73994f43e8f6aada2cbb3e91f34de9b0b4cd0e343639223145a2bae7b82020787ad3a6d5ac02a5d18cbcae805842816b213e4037435b1f36b1fa8a522d4a7ae398ef634af65ba3dee0668125789949933de014278ee1d78df1da74ea9f2924fb6bf4390a8beedd406123bc024de17054c933cede012515f645de468ed7154982f58c0448faf49ac10d13bb53c07da1b799eaa3147cc558a9c6273c8a9a021bc80a38417144426bd35df99a5f610748f06dc4604241168528ddd4003fdcd81d94bcb1b33fa810c93955b393050993a5ddc968bec3fa6309af0bd926b32e67074218ed28a89cd8cc3d37091c458d39c0d71343f95179d537e115c4fa0255d1845247121d9191ab2a556b5a92a6d807b1213e3e935b56cd4019c7fb1bbf724ab25ebe7e7d1dd0dd0bce0e80b4cf74cec52b0d5ca3327dd0203ddd13b9db1e41b4789c615afe25f5879698682de1780ae4fff295d50d7b1cfce3eed7e4b6ec3eabd91b978cd5c6ccdc28bd911588962f8b782acdfd2bb09a2aa84cf6c6457d3b9b8b6f7211e4a62c19eb26962183b8355766dad395eb83425786e7f9de4e0a25b56842adf90b781bf3d54006ed857a4d60746a2026cab70f780a6becc6b211a862372a5051aa9c092c27711f43bc975b33f59bb801cc3df4757331f96c7c501061a1d1631f450f7980cc27754acc27d55dfe77215382;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8a98abbcd792a804b8c680d0035da6da5f33899ccaa676f2d2955d9ce77bc15d505b19fac0f4200a65e9a992319809702c8c2a75634607897f5142224331ae47630092546f71b0d5f04f22f0cde4f10bfc3d52b16cf54e9ca891f63cdd33f0b7fb6883d6cb997085e8a7db60207934e1f83d84ad31f4015f713796969a1ec837e256b70b9717d338e1871139793f60f974e6c0d5fa05021692c4b55fabd1045e384c45ca10d3088ef4ff0ecb4490e813f7932e52d0cf7c525f5c5b6bf17db60881b0631aa5de90da2b14ee9ae10e1ab30626e8b8b3f32d62cc1bf8a03c7efc33d1006e29031c45d0d1877b0c53e189cb57af697d8efc24b89330256c8831eb471c26167048710eb33efd6d7d23be7a5766f75aedf04afd151e82599a480ff766812d90f0765ecdf4a4cc36a99c7738d48e920ac3cfd7afd22a2f75922453b588a73790c3b750f660a1836906d0a4e60d439398b6399937204f4b8fa63e26ac13de7c41573d52c325f20fc80881eb82cab8e412e410a7cf3f2da115db9c1e76c397b237ffbe7561a8facd40cc3b34397ccac1c4aff09119d769a63079b1df92572003ff63c80381c1988fc5e93c86b344d3a680a5491cb910da3a17327b6079238f08f4ee6ccbad4fa327b277b98318e7f168f3bc0d1f3966a26cc49a171b3be0b0af708a14958ab9ab860a1a73b836a92e68654f44e64c149447e70c71cacf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3cad31e7f38e1419dc99616fb05479d92ccac7b27647a13231faf11b742e3637ca529b2dc780e8a41163c8aee7a46a81438ecc9a70644167a185f561929174021e27ae4dacf61d6cae04f4d89f77d26d3a05a7addb654bf3e5d0c6acf59752d283d4ea6f53c1274c7d6bae3bdaa9ed4742727501064beca824987f6efe317015b6ea6ac6feb2d235bca39c7d8c7797e500e4b2352758051d5ecca6e0b67c3cf748a9551e9b1a02c42ba14f1a7d0f2beaefe0d590577f017b8cf69bdf46a0e94765f45b75b7fbc3f7a79e6ef68b47b002b4a42ed5a5a4251905383eeb7e9de9a2177fa16b012f62e1dee2f0b0aaff1d8a884edd63ca9591f56dbc9e35a87203c9193f49624905a1aa9e4489f28eb0dcd763aff2abc131e7b350fa2de0a98ec2e63b9f0769473c5541ec8cf234a446b6fd2774c9b97ceeeb4636b1b8f0199bea968b87055a923c082caf627369c0e81feebce870c065b84c1f1bfeaba279221091c15bd29a7d16e8cb518d2a0030b53184f6a680fd0e242ace969d6956ce169bbe57fabfe88c230ee370a88c5addc15a832e36d20228fd0e4a8e2030c78f8b95924a2487e6396ae866e1595007fed6c82ef66f038595e1284c9e892dad317028a5d19ec56749f93d4244e72a5e0a6cfc9928c3df3a745d207b780ee9422d8e953432582bcf06b1e1dc4e1314d999fa71344b0bd13d7c65e905f57be13bdecde71d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd113bb310c117025149c0819caa8ffc52dbb1b6233e3eeca6bf0d708f202cc3e447ec1ca09a527836393906f77dfb5a6ec8504f01b647e73af7e25204d786caba713114707060101289669ac735dcf8010103d9faef4daca72c7a947d55332e9914e79fbd27b195d9482acad8bc7695a8b23daaa17d0ca0c193778780e2ed4100af22c4753ba2dc2186329ac359c335e789cfe89547e70321ef213fdc3b01802acf36e5044e384b5e55be2a59638be0fd5f02cad53545478512d274ae48453cdb8b8c6a1a03fcbfa532505d6318d32a7f9380e2dfcd553a819706455d2c9e3975e867153dade39c2ce94d4d8c8462132f966564bfd78e5dd451006899788f5b5e84a74117df610b9a65ef41c139b49b27521f217ec6380e860916e82173cd29ac9217b11066d2f36c7f487a6cfb2e0e3bd24849aa342990dfc7b16f7e2dd473f2211ef132313404022f13c2b7a90cbbcc861f631f5275bc2b82cfb88f5b6863a0814f105a1168c079d0cf89b97394ad5028d73294641c79a9a0b8403b0f09463e12aa1cb019f6eb0303f92e4c7c6b824c069bc869d978900dd302af5fb1acc328d607952a69371e8a48673a614dfe09a150bac958e15311071d63ad806c3392eca292b53d4beddf523c2d1b23582d504c7f2719ffae7b1e59d18e517f62d5b5bd0181ed1cf3010fae7fcd2638f24e0491805e94ecf94a61a9709b9502c43e066;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3edc1fd5b897eb81eaa03f334edcb428d0013f26fe0fbc5ec3e4336a6765a70d5cf4027c99941845ea354994dea093b06e7b9308c704758e0bf553818d076325629506bd16927c28a56ae1e382c3959cdabe80e3954474a4df75b36ca1092389ea2f9f3ae927a22fe77d45997c755c7396c86b9bc3445670e8812faa2b39a8092d49d5dd686b94a21d0ee281ed71830063c62d34ca1e881a7f09a9b556b9b24078dd5fe94c0354923cde34556a90889d365c7fb85ec1201d3ab51fa2e5c53d16a12798fdab999867e6dcb08d291bb5e5db0b33bc1dbb564a7e8d261dbda9d058871a2b22a86c2af7b90e194bdd39afcb884e0c0a91291b85a1a76c1af870a1317061f3bdb15f2f5947170b493181c7f94312407f37a37ba79aeb88c09af6604a20b636cd284f27a6b7da1458a362de206dadca9d75bbc5eb50df04b9de4129416534f3f2b226fea5e29fc9ad9fed62caa8747cb468def20b3c55af3bf49d286167909a84995294eef89959e3f852087ea4c80ba1441889e65efc2cfe49bee7608ad07ee1147338925cf2ac3f1abcaea512a9f9ad9b7c766824a1c660813fd74bed4c04e45c041bd13f8d1edd1c1b16ee58ce00393ca9852c1da291b6a0bbeec36c9464fde48cbbebd88abe75156485f1d7f110e1f19d88ff2be84ed2d33568076fd8c9b203213eef50b41ccfe13abd47941ec6338a44b57ccb2db9459ef65325;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3eaed66849c18f1d90c731e2128f1fc58db20c74924644505c9dd6ab1d665c0d04bdc8d2daaa7b4806fb5bccb1b44a8a15778326076bc75c0d9c5f24eb76025204d504c0d0e8af69c68be997e43f69bd85cf7481581e1d96b73526ae53297deb8b0b32b8c2f449e7e7baaf590b177416f9f5ffbd7160858ad0edcf2383727cde1f27556f514cc82e9d5bc0fb36105af75630f0d55d8f4569aaa2a1e7b32e1b25f8931c24bcc6078d729e8644a7c4919d1080cffb9c7f393996db32fb20ec8f5f5a5fa03b838f2d376c699fb599eaa2b16028fb8d5604ad7d55b69ebb30ef9009e2844605caa8632a85acbbc755feab2bfd8d107a30611a88e81d6085acf0660a7b38bdcb822deac4471729559b02a94b9d1dfcf12a32676fe83ca2f54e7ba1926d611e7110fc824ddc52ee598a7884aaf926660d0dde2ab1c963948bc0d11bc2f7c93795d201249f79e6cc77bd1bb08871871155ce95655486a1d97dca594c01f12d5d3abd95017d7d70cb031c55ad7abe23bc4a293702a2a348ff66154d0876a938d4678d370ca7fe597a351185eee95a20e62a3b56c962649b25a2d398e6d5e98265db34ee5cca867774f6dad075e9c0d1cb58b78d39898ef1601d63c84f3faf3ba0e3bb6a84e6c757bd9337099860bd83e79b57f8008da98c19d1a910180d7b830959ae6a8d34b29a1e6a015d709047864186a1c80d8d09dc0142e059edca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf23017f094589bfc0c0f7fab378b050a559a4564f23de35942130fd24af57f6d3f92faf4b7e97656c60558431fb293a74a5c031720348a22a4eefe0d0b046d7adf526f1b0a60115d640cc6c70b22fd72da52ad1da1df8c7cd83a8da126883f1b83ee79f8dd33f1d4e4ee742dd4946395086f57ed7434045b09d8efc619434088dc92afc6f599af35ea4903704f7bfa00f7a2da5f8653c12d5166a769c4db463ef596221da77fbe195496af074ea594233b4b100a2758364205c655314a344e13b23987928ddbdd6dc54ef0b350044d81248407c0e7ef5a9829c7ef2e858e5d5d6811313452b35a7e31bb7d7d054d8127870f990eebb5aee86ed490681dfd726b8d7b5dbb21847d08bcc3e8f1ea0f12eb1fb1a07c580d2d7e89c8bfe66b58fa4c4a09b38e21e99d70d2dd4849d659b01892e8ac0a0088e6a474b1ba9ea45af3f5e69eff9c673ce6bd18058fb92f5dd556cc619408f097f8f8fc5ca340f5975630a5cd7e6ec75983f13e1821e8846d28eb8e3ca3254c84c7c56a34e43ae52cb00a2efed049dd63e676dbbea9c677b258c71d685cf6e1b14cfab80f7e3013e798f0bd2e15bebd3be5c787bad6b0d7db8a1bf377c814793993ba966bf3b812fca67f187c82e68e896833af7fba7416d8d957b6c9ce9838b9c95f49f411919713fe11193dedec7ee03a842d91d6703af2e94f7129df917a9d349371d0aac4b1cbf362;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha3f2ab1cd2a53cb7f20e129027ac17ee6e0cb74a29a45288f62cb666f2058e70263cfddbfc067b57e2b58b5265ec636a2a73592f5598f66e17707d7ba53bd405dae301e1961bc908bd90380eee3428331a944b6ef1958ac87e6ef687f149a73c84d5fb5007e7bf0f7eca99d2235ddafe6daeab8b934f8db6f67a915ecc67da3ce7d98f99687330b87ff6239750ce829f2745f6f01f09a1a6c42e029eda789e4837c23e40445a3e0b764cc3fe415ca124b015b57b7497ca7f819fd1445dbd4f5abd8d93054ef8e104bedb0a111e5772459878bd199fef5cf72477d1230bd265e20eeb120a467195a43c41c74b4878caaf355227b02d4299de9940b5e762e892581934d12fa2aaa15d1e14fe8ccf74d3b507cfdd4478dd16f4714a4b497c5ad96e277f9604854ed92908ed5a8e4307ef8b6561d7935cf3252cd00254ec2a3e98e5b9d48bea804ef9b8f32a834fa6e43c3610672cca9f5b3116c6adf307b8e01046e28bda36b1f229aa6738bd273588ea01302e53b380cd401c5d14452173fbb9816a05cff67ef69f00cb035a9ade60a84370938e9eafce2d4f2e0246cc83a3e1f2285e2718be279dafa8c459e2a938dbe07a54f4cd23b6747c39b2cd3f65ebaa9c7d410280cb7b6d9acbc22cb1b577fe3dd164482d9af574e4c36795afbf9052f7ac4d713c46bbbe0c305a9aa56c686b625871a015931260f1ffe5e4a3dec2de2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd6852c09140f45436186d7c9f408532db9f5c4dddf615fc25d4fba83cc536af94b85d8ef684a1c74b32f9dd8ac3726ec07112a108244cd5cd17cd399f28bf25b0678411e88edf489373e36dabb8441a281e444ae06f233845dd9278ef0340b230e9dcf9e6de7770d38b50acaaa9aa357068eb5ee1cf66ac52fafa62e9c0fbbab2e63d7612b11a3050908f32c6992ac1d671a7ba72abb35fdc66985ccdfb05342476b0f87b3a4d3acddeaafe42f9bb09615514e53e00125e3ff2bde49de1cbfa98d31d58f959d3f84db80e0415dc2aeb9aea5df896fec1fa2a4b71ea050877dce56b180a24f7ad36c83a2a51c6df2ef602d99b35862d7e717c7226bea9fad0c49285db3a68de016495d3441b0d41d6084c368b7b974c6649004d8d98c7a2dc91711f7d37e324b9c998b192cd84175d0daf8875b51ec0dc6ae569e24be366578f00c837785658c52b6676ad1212530a1935a3a752d910101899ad8480f972eb250d21863fb70b085eaf297cf0892b0167289f03a120f709024e3369321dc6fd20e065fab21669ec2458f9c8564b7f77e70ab345800e2050b4e926537328e2fc87e7bc58dd1cc11f4f71faa1a4735deb6fcf62385ef7f850b88cc77ec70f66991d8825dfdc765f35ab4a5502057c634b2d9592a4a4b302c74dfaa0c80cc9c42d9666547f6737a6de6d03896ef9bd2802228fe9657d7241591c6071fc34451387eb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h523d6ff444d9e56833d8842ed50e3a9f37173793cc91cce6798b8232ada131b804d8157bd0cb923c4676bb66ad5fc4f681f1673959afda6e365855d7a9c5dcaf7fb5cf3803de295431aeea1fcc03e0d91a49f4d4671107241e26d15baeef8736c94fe024454d29996005e31e82625922bf9d249bff36900d2a1b39c6618182681876be9c50f2fc0bec3b20856d3890eb9f4bf96c317962a7a348cdc4f08e6f810817377b6114ec9045e03b152ed95df27c48b77d064f2c5af9646f6dfc197682a028100ad27d921b32ab2cbd5f1909bd9066f9c155befa8db0840dc7e2f7a5090f891dc97fd08a4e4c6d091de2afeed0c7200e65a48cf1c12b73522ffd7e67d4113128d031dd7aab7d4e04183b272f7a789780788aecfbc3083399d621859f044bb093ca05b71e80d97a02efa5a360ca78018f84b711b5e550c18046ebc15574e15209e3e1f6b19d43095f034c43fe0192aabb5b9733c2cda8ba8a872ddbf593bdff3ad93f9866f85e1e5a4dce9d71961c54cd31c8bf9abc964fb9cf7852f6a00b0d21361fd50e446d94de97304a5e969eb74948943a855c449c2f17e29b60f7173764d7e3c0cd58914440c907b72acce3d96621e2e8e1813b1bb1d06792dee56d774592557ab003d2ed7c074cca062f5e5837ddfed6975079d799012538db2bd26e0cd4a092eaa02582d02ac4de074c851635000d023598485efca32d84f83a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7914ac98984a0be96ea03afc3afdd5abaf00c5bc23cf1ac6593d8995497d72c6bfef80a1fcba7d37effc316b6bfd85ff16c80a3dac80b96fe1ffac6d352bc8be47c7bcef90b40b46266685df43fc3d765de47ccdc45758bf97ded2eaf95aab0d83a7b34a35e93a7897400bd1535307c2ada6911550211459fba6075ae5d5e9914b3ae85bc125163697a82d5dbfd29c73d99d8d39a60f95022aad79296e7b35e5e368047113d60677b02958eee60c60d5facd6b0c139530637bead5cb041dd439d9c2324fe293b31842ae96b1707ca285875af41b1b9e7abd20b064fb943e8861ac3c9f3911ebc8e0cbe26842ff5cb25716b276edf85749264a415e576cff6b49882f0408d9fe47841d916af4a9419b15eeb8c965c0bc2783e7bc9a07962adc5552812113a7cd1e62993a4a93005f0ef66e926c171b5bed4b391747157ca8b102d233f3ce106cd1fe58098678795c33f07562e7e811c0c1e30e605e029e1e054bcd572f8bbad7e4eabcaca2d8cf246bd3b2522c7f13d228aa8dc633db667059809075ce79dce3853a8d594874787720542a521856317e0bfb2895ba7fdcd995dfa5ddf094cd112c1297f786792d90aa327fff169959f0402867617464becbb6ce58c40b249590922262316d2d6e0aa24616590a4557887f029f1c2d8ed1ee0c70fb28265c4d8f6da73a50e974af2029f147cf4b480427cef2ac1a0c6844072054;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3a7478ba869dfa1de31f4d380079440540cb66c9b7c135b16e8413a65474bb439bc091de548fba35a5c6297d4b852052eebf34a8a69a0fcb5e0713385b8169b0a6d6a219ff007bf4a48e2f1817d78e94f5a63e5c4437cafaf7cdbb7412d71ce79e575feeb5faee6a9d0cdde1f8c0ed1db3878b88e6a3b100ef21a8ce04eaa714c5187f53bde131aef4138f9b6dea61de05e8aa7604b6d364ace8991aab1be53de7cc0cfe61bac13c20637b1f64d5d3ab578614921f12ad551a8d7dd4a7fda2797579490a13190431f8bc49fbf30dad6ee72381a00030a005c90eaab7214eefcf0073320724a0f36b18f49dcc36cc212ddcca937ac6de2947a7f187a5db358a6315e42d13569293a9be3ba548f1cfcfaeceab47b79f98830041065e43a79ee2c9c42a9764e7b06abcd3b1bcb045e76e02480553ffe92648e0d38775b403d5a09d53ee1423e80a34abfd302fb3dce803249c2e9c8061669fcf06856cbd6334cebf52780e2b0f414869c0cd5ec3a1a791b6e108e6a4317eb6b57f427351432faf6aa74ad4893c2f218aca73bfc3652635b8541ce630f467c803773d925b4e78d422c5701c35486043e4b91ac49669dd0235be489188a9a4f19009290af44e1758985c0ea5eb249ca8583c4584b09c3ecd39486f599cbb066cc18a80643cfc355fdcfd75d528daf834ae30d5d04a830bfcb1b8af1c433e31165fa7c8f12d0e9bd45e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h30d27d7a384c4044afe67532f8485994426d6712373de1a1f68760f465f1547772431f1bc6f9acffa54f01d73da25a1e07be7fff045cdb58f76f2dd13b5d47d66bc02ea21064c0344fe41cf2dfeb1e5f1b0cf3a5fefecf6558b30b19826d25352b2d92e5f34960db7fbd11b1f0601991013dda288a80b742fc5462417c42f59bfefb1505e8d7fdf4ab1fad5a7bd97f12139a4c468a5f7620c40dca0bd7e61263feb7d220bac60f9943ddb129d7bf2ddd9c76b3c21cfa2269543d1da86e67eebd17ec6ddc66dec134d4645ba1b64b99ce77528e897231ebd73933419253ad420c76c4802eefa6c4b99ee3006826624fce9baa1042ba23058350ccfa2654239f745c1942e736222fa8e94b8223c78cc92d1b3354bbd5b8f48725d78ddb8543ad48da94f4a498586f8fa6cc2fea4f9db61c5c2d9ee558661e074540319f933163b31912056fe1361d86a7e7ca393988c7cb8794a71592eec4d944eb3be041d84925a1add0c748baf8e3aa4fc977cbf2726f590d3068b345140d24073bc7f43b8d7a9d9219dc62507e5222554077cde8a164e1dccf4032475582c7d60940c1debc7d2fb7e616cf06aebaeeb4db0c2907d316e1542afbd1cbc91eeefb715ad04837347bea2cdd23e3b265a86a42ce73923b64ce51c226d52b24810d55826ec7c2386cf8c3f49ecf3d1b35d24c4bfba19ea64ae7ab90bb5fe7e9bebb9b78112280a6a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h417668e62baebd4867e74262ae6c43005e04443bdad3f81611b8998b48ad4a09aaec8e3ce827e6039fd217287f28c8cfdbc99064ec2834c7a16587edc4b2a7c8a10a6c59c338f83344513f28d0bdff59258c6b1551ac241fd009282f27c8bf64b6b99017d7f231dd9a3a2b366861a2f8514cb23cb06ff33ca0b0094612c85f1aa963a6a935a0ba624fb3acf1795ada358f26d839a02f4418c63408ca5920efa8fa095eec4c5d220f33a6a5238b0b7e7dcbe3c1da4495f2c0d655239cf44cc1065690b53c48cbc555d83bdf41d412745096eb7dead5d738170094edac37748669be0ec2cf4a979120988628cc26f9fbf444bfe603806b817f81fa437188763c17c46134fc220161a0866d74b8de0e2ac72231782ea307b5450fb8fb74286827243c22d9923871745766ebc12952a376bd7b4e4423d6253bc7d0d2c17df9dd48a2f61ea8a672446804eacfdafb9e2ccc834f75401ad07d58aa9eb74fc18edf32818e32198b5fed898ec08a25d357c2a8dcdd31fb5dbec9d332139db4955d3182ce4fcbe13e1709b26b027ebed7a7c4afe07a7d8d2a6985db4c01a27abf962cf7fb750e9700038ec2fd744295406cd31285e15304b22dd58e3caaa225a9c6e7e3911f57296eceb3a2beb8127a39194e7c6a1cf51a5231c2e0463f8a7e4871f39f6dd7eff84e6c857014807516bb108b9c0d994772b043a31f55afd088ed419dd984;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfdf24fe70fe896e99b667ff9681157c633452542fef2f99f48e3a7b27d609b5211ad7e25b92fa5a55a42cb5b9e88df9f7b4fb9376fde9c0234ded89402c7627c91f65f686698096b9f814b49d59bacdd9f33aaa7702db33492c016738673c43a60e8f45342573b9c3f4908663e218e0df63f483bf1fca8ab3806871dd9128457b6109bc3996d8ca93a95f7ab465b189f1a2224c966c0810122b00a4f7c0bd6679e528f1703856226f1997e13bd4fe4411ade80a681d8f902f367d2e18c4c7400929a1b465048421a3799a2638e3914b9d84e7e228a9c609c3b814de7ac061606aca408e660ee8f743e2c8d86b6b855bc54549cdbee15ce9f4ddb3a72421166cfb644eb53992a7abc809ef982d272c9afbb1b34496cd92b551786ad8b642431a39c8e3db9ecfc8d63e6ab7632c8025a20c166b1f6a4b73f7d8d7d788afee87fdad6769155c779a26499d9257cde0fed63173c01d0f616c3d205a810ec72f6febef040ff9f17878741f842edc3d4c5d8d6cb89624757f87d68ee47143b865e9654bd4b0878d22433e238ce22aed9288d53abf45e53245e85742fb582bcb9db88d41dc1945890b422c75bcf307e8a547ca0d759e32298a1694b98c8f9edcad30f0489131d76fa14f90422b9d297d600bebd1cbe606ad3fae1842421af64b6f6d4f794d40b7e34f696e17531763c2b01077c0f7fbbb54714c3d792196331f932488f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h73bc3058f30f4d17ec7f9f6ab4bfe9c5e607ea83a42839be4293229b1a340b276f2f71cd287b7418f7af35ba3318e1a12214dadec4b009c7090065fd1237ef69699327708596a21722f93d6534f7c9b6d1e425096936e2ad4c44f4ab6d0c787616d4d69553bd5da7cd18a8425ed8010ea0490419a52781048ca633c8f4144f75d662b7a47de3c5f640c414f82dc74a821996608d67a767a4940b71816eda3c3cf95d11ef3ad4d9835b75e026332d642f9dcc0448408d2e06b147983440ed8924dcfbe9ef587420ad6911ebfd748a0a34e4db27a0fa3681ae09571637f9175b6d18b455baa58380d59bcc3f6b3145e2be77f3ed3d03877a801703fd37394988ded0b2caa63c307fbcc58ac401a6a2623ef38c50424ebe5749d344ffbe948127b818999fa6908bbc76c08385a75c35503c03f3b1a667ebcc0cd28c486f7481a61ecc7bab3d327d5e1cb2e06605aa1909e9bdc1175cfe4f0e3808f8788dd054a1491839682baaf7b60292e07ee4da4f0ce5468daaa661063c7580536f81da66e3f013c230367b96e764794e3e51cd79891a2597ee3caf6cf0ee7f72b9d4673a1b1fe8c17378f40bda8c3a3434af2419bb7ffbec475bd15298032868af62f7ec97f92fd59fba6ac204e1e7e0687a3b9803604b355984cce715d0a3c2dad30e44391b5f4e71abcde04e0c1a19494b7bd91281e7550c634b40e7f6a56cca46e4ac519;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd65e058c1c22b6926775a8d1fdfa66f59a6716452d280501e369eeb21b463781a16faaab331d25e86af2e3ef5493063562a41467a4c21c3d21142d7a2ba81d406ca7e3d2d82ebb466557f1e8ede37a86818e5a47ec388d6c4eb9e95412c93c74c7ac7c1a79f592376d8cdc2c308815e8e7162d0fe6d196e7c324250cb782e4541a36d93c085b786d3f4fc170e8d49efafbb0bff4d9f116d5c7ff44e67089a038bfbb014f5365a5c4ff36e121150930617416cea779f32bf536c481a996fea3ec69c7f2b5bb1537d53c1152d1a112d512721481d5142a07b28737a78b48885df2622afdbbdca3fb7e167bec8a9d0c29d7d45e3dbb2895d7ced2632dada016c4560ce1335a4e218b3cf14b4c72145964780ad4931ba9e51b33302d36fda51b1bd77dbb7aa94efe437b0667760e2497583f064d3f3a43a2ef25dda93383175370ec807d3e2062039f9243cd1e387605cfc1dbb66abbda3f2ff55834f1f6a730219fc46e86caa1d13e1ebc2f0ce7d42fee7401b73e0b867b026d3f535a131e160532d3558a8b9727b4c08cb7d41d0f340e902fe8dacb868b2a29fdeca38444ea079c69993153cc4c10aefbf4304bf6e43bfc79d5a471751f4f42b94de98a858083edc9fd67519c7d4304831d63c9f7e6321ff6fdc6ca0e4003c95db21fbd82a7100a9f03a6a469a416b4b100162ec58c034aa79e50e2b63cfce8bcea7c33b6743559;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb10d0c60b89df5009cfa297ef0b80d8a89ac9905d53225ba758315d54d3ef1aeb4c30b58f5a5ac87434b49a2242e913881cccb8fa42f792a4486a9a86d6c43b122aaa07aa3bbe3bd440387fce139d60c63d33b84f2f74a3c0f09d2ba2eb900fde7f0aa4516c6ca00a0c6ea5f5c725d3ae9455160edf3cce52688297cc50d16360ee0d3f5da0bb3e2d534742a32ee4fb3f974048fb7ec0f98d908ecddb3900a6a91f00f9a32d4dfbf3160fe7c3a7b43b726c73ebcb4d0a87e8f3a3949b66ba8c988d988b8637d4baae46727cbf0c9a2543060e3acf8a634cac7075f3df9f649f55652b54364f818f8ca710942320b407f6fb48f2789d693c2678371bd94a6bc727a681ced62210fc27b485f785bdd5648525b0a5fb9ceaede6224b585cdc17520b3b065ec0545fcf62ecadffd5e2d514e074832e4f81816b98ffe4f7ddef550d3d7cfc28b599281acd870eaa92210939dc4c36177bfbe3e4b3ccadf5251d6291fa4752f87d241739ba1b880949c67d1738ad4c4064aa921dd66496e2a830484ccfc3c12c5575cbc8af3264eaa46d1396a3b668d629e154a672e214fdc79e5e341635af4c5307a90c2b1a4a5ee964b455e3630490cfe49a507b0d8a74491d45228ad259b96968a2eafe8860328c9de7d79045e675f0b91d4b47a28a44e9a4d317f56ea4889d8bd4521487fab737fff1b3a5c47a776476a765b5f43a944a0028b18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h777c1f9a708824f300ccb7a4c334321914118c5a4b00d3a173da60da0590653b390d51e35a7c1e966c5290564b09fce93313678fbd1db350487fce5436a453a6ee92f31263a9b62c715b7d4eebc62aa92f22d2e304388be44f78a729ad3d7608215ed5aba69dfb03eb835a8efafb12ee54e211e9f54d09872a59fb43f312b0a88fd9ac493016ec57a1ccdb0a3892f50bfa08c791882c810c85a59dbacb02a9168878606c4a6ebe9cf1f0911831c5bae0d15dddb25ce4a955256985cdce89ebd421bf6bf80a466bae01ce431eb66d28d52d0b69e75053466e71279b2573d36db5e153dc50c2a4c66bc396dd061778510c29e9bc98848aa915b161b16d1e8578b350052749c5165eef3007cf86166bb53829f4d1c8269533f58e7ef875ec10ebe84d35e19beae0c746413ff87d198b0d54aeed0b38ca1cc1dc70c5da45e549ebf11cadab340284b0b4d8f42b453d622c05494cc5690be0da124aea0e8ba750df1e00e03cb56e3b358aeafd6de5b0628445da2b729dbb030b207da7daf7d22d9f8e9dd27c0cb447b468ecbc861f15030bc6156cccbb79d6c9fa0eb8535bbb53ee4ecfc5777967e2bb1f51cbb7ee2da97f280f904023a9327f6464bd995966b13b8a5861796a1bfca70715f0762e17b29d38b8791d78444428823ec209bf3dbb168370111960fa8524811dbccfc7f5f5a8a33f9f9cfc2f66a5cf9f4971b8ffe06f1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2be50d9a451a068d12c75f73d5f741504c870a84563e3ab75a2fdaf8e6ce0a91d00977f257c233a193b99ad73ef1d0cc317216b70cbfa8b366e136e190a6bfe620f2618434c44a888d6f4514f6cb437999354fc79697c1461bccb3e23ffaac38e71c5f97a90cbba9933a390ce3e2342238d1aa5e9ef1a15008bab057898255dc5108cddb085a15f4554918bad81edf5a0ec1666794834c7a94033120d34282fdc3eb9d40e67be6b640a54e3c04f02c7bdc6f87684f4e4dac39c569b10d77d9b2a89276ad12a00a6b287fca7acba1f2bf359ef3ab915158a4fbb677bc85d1990ec85e9217073780d6387855d62dd390f9d063b92c71312dab5d850dace24a308f1c641c07adb2955d6b4b768ff091e40d9bed1037803c8013418775fb9bcd37b567cbea877842075af655a1e579180b038241662c2632bd4fe95e9a08ae6e0e9c68960750f701d861c7eb1882dc0263212e8104359565dcc41cd62c39e8cb7107772da1c1b76a3a8dee045ce50824fb20d09505e66e3e1fe1e804c468960abcd9b67152277832ee0194431b899ae1b0c5610d594c3982cf2869777352f6d8c5b48e6f26bafd767a312543d422c14338c9b895cd72975bf186b58e231f922d719a329cebe5260678e3bb187a4d33198732b5d78e7794a68b741f2ce10d062e794e78f6bd963610eb243715593e02da0b0b9430418d152c0971d4ae9a3350fca29a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3228007138284475f09c202323a7ab44f2be05a64ae0dce40c1590e9cea996c1cadc44ff6085450b24a1de1398bb371fa935b4a07705d162e3fe19da0052a0886d59abc0985df0212b376df52f5bec4ff0b232c16022be8630bb5e207e3a22a90d97957da4110c575216089c0668feac87e063b10ac336f8c7b50ab3df3859325d3b93d439968a50f92ff14df4589d467916eed95ba4e21a70f0a7cb0cf9100c4ed4a952466f3efd0f41a4b0dcb198206ea6530a20ee58e01dd16a2b3e15d730bfdd27e9e04830364ede668fcf3f31efb31b0a62a299460261c3a6af15947304f717070e68a8758b40fb479087767dfe9a5ac5af8994c9c5548c74f2fdd4a1faac93ce48d49e8099728d611c64db341dccfff01bfdab76784c6607798771a4db8f707e96a268b3060874e971f76a1d462a6a949c3360f4afe557e0b60d68b80980846792e2baae7d4dcc01f21fe1f8473a8002dd06cddcebc07967e298fff8379fefcb127f983b5060ae031cb9677f1c0277917123407cf86057dfcb9a80046a921e0e8179b7905a52eb44d22a36f6579b97c31a252158f23fab7f475e165dc7119feb0ce80a1cab7d1d6f30d1f4e4bab69345ea6a40170e87c7c7eaa90a7c781c272dc7117f21341ec7fa7da90ef09833ce5825c8719a4f45c7a71da28f1eabd6c962b6fe921b656d4b25750586776f6bef7b62872f1503b15cb618c4543951;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8a67f397cf991835e7b41418022b4809374c731098c9a1dfb849a5bf33db569bfe2929fa6bdc3c5def67acbf464f706f20d81cdbdd26f6638c28f1c346e3b165d0068fa692d41f9d1454f70a10d88366be6a8c7a8a47290da3324305f7c8f0379a4f547b8f8139eba661e56f1be905d7314fb06142e4811c9cc247291f30fdf8ef1af12d668d7ae03dd64cbfe1775a3e947ea031861c5be8addc2da153a560ff7cfec07098ad456dda3208a78106791befad518ad06963e963d12cca81629f45c2fcb028e951207ee127a92e67b40647082cbd4aa58a95a92ee85eaddd6005bc627966e5598e9d4f39160613a19ec150138a5cc24407acbcf56200bd408774763e4a4e064f023930fd4a0217a30f42d9d8cf1d65028063690db5a56bc4f881456fd3ea3f1f44a7a6eb4bd874bf5967b0413c9c93f4a7090178510f6ae7ab4381f42a824372c6fe9e5aaa2ee236199036b160643bbd5b24ee2d76e6dfb8596f4c0f9de7a56d927cd24ce8a9e0084e924bfd58ae4a91aca3ae3e6ee4a5a2ba2ad229eb9f0989d4a225bc9d601a2238c5ad33c836da5f2d5184743b7bdef42e497716ce8b5c166760c9f68bc6057c0f5ccbaa7cb16135989dd0554aeab41fa15c612338d0d0d01b8d01e28d3f78b5c73a944aa2c55fc63816191406849be099f9a1ce8d936c0681152abffcd20e1bad27641d8f50b24888ce9809d163f5c4e5c755;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc8b2b114843fa293a488d79e5ad153a7c688558bc2dbcd99b45735ab4010cce3a0da3ee060130a8f370afb5b346440fd3037f26407c1c2397892d44fb95ac1a3694cefe6131a52d9b2620a0b1111f4aae6071c4592c2c6fe63d743e38cf76401097353956f8fe6e736b2af884e0db2a5668943639474a9cc3413312b836ce22f08634c44228fe3a7764d93d272e25235c6b1984c302b6777941c75a234043519ac93ff714baf7eb91ad06080473004643f72b12f9dc38f54f955ec2e206b5592c6042001426e724349c44ce633f767e04bfecca7743753cd58a97b3684d6b8951f56a97c590d9102cdf13d169a202e3e6d6b0616f84e1da77f881833a59c34345220e21fa365e4e9767d9576dd41b7f7369c9c17d10205f40a8b1ececd238fbd644625b0a26b21f86a2da449eca414071ea1870c3ebfbf5bd7b42baae3a832269c5ce411bd0a48cc98dec9851475920684c901e069468a1733474876d232eebd58d3e8c7ac59ecd4c481f0fe96bcf92f0923dd9c041cdaabcffecfd3d56b48119b0b206133a0f8d5f484848ff6945a3df76355a914bf44d0ccbb2ec993addfbd3d3db620c30f874528709d84f1675f726c627905841374c0ebbb485f7ef054d523e879072112b11c3d8821b57809ea7f634ed915530e6634880130f3794bb5a9c77885aaf4bc085600fb6b564e430a5ba1002bfe1d9754a220cdb09ca4a7698f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9eb49aae34628fb6876df938334e9e16dbc613db6ed15c2438c30a1c8e25432265ad8908bae37ba8b71319d28253845479a6cddb4bff983189472c204efa885e4e3fec5f1d7a0c8bc34cb3c8d149636c54d530b90c233fb53e9d742776ef303d822991a9a511a819b1c5530bf6d81c5f2049d502181c399d301c8fce7c2500209a182a42b7f9bd94e303dfd6b577faf684e6c82db020c1f1594703bf0a9530f2c800a34984687cbfd65bf695b34a6fa9ad4ccb7e1b6101bcae09764e10492ac3efa31eebd5c9d23980cb0660a405495a7b7ab3956448d300af05aab5ccd2cb74dbd4fb0120221e0d1c3d37f3c1acc48e8e06753d59ba9f93e9fd5ecf17aef52a1145a8889784ebc8e48355f03f976a40e268abd622d72f501607749de55533280dfbfea84723fd71813d264c182fcb8152dbd3b33409bd51e820cc58533d2c892b33b8acf37cab76a570380a3d2961e525fd8c616bca13aff44080e79746d830ec6dc5ed29ab3a1299e6029a5b73add9c5b0ae671806b78603ab16aee0e2a94eb5a64854cbc2c86febf1b76775a7303fa701bfd5e5d24549cbbb0eae5f5273cd5c83f32c2e9d58f06790280f2a037d6925a9234ace2045da8014d00ecbf9393ee47fd6cac22a1533a43c4e63d2bd19aa6d8df65bf5c5329d5643f574dc78f6eae489a4d8d3aeb7ab174faead0d066fd4609010e89089b93f3ec71766665905a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5f1ecf250ff19b73940fc8efa01a78b5af38f30fc21c5488bf1d295dbb0e6490a127a5d87c5aa6a9aef8ebd2b622c716ba55f1141540eeff86b885f15282db38a7a0f6153e54de4526ecebafcb914e7badccc9640c7e08b59c01d67ee56e7da9002ad6ff222fd8b2b2fd85f1e7bf8332bd07226f31f37d43c85d28757927a1f66f93cb4cf9718b1c4da5aba1780d8424ad23ac1d24626e4373089b1388800acbf5b005263e1c82cc5dac5654d9222ab2586a9d6b9e348be16c11ded504dfab43cf03f03fe01faaea6d289fe43f907a9a70b51f7847e2c08d02df6127912bb59ed706c2a678beb3c6c7001542bd3f7472a87b934ea910b1500ec8c128787f5538cfa07a3e25452ff863e70929014cbf449a59d0b34224a223700ec6871b5508033287e3c8d6dc222f06890e33c864092f28b02088bc8eaf8bfc9cb56c5509a9ff335ac3680c0214a2abb8f8dab3a83f1831b14a4b438ea61a71f373a559ba8b43e4b621504b67c82da43f0782d9c54110a9f199dffdbe3e109a2cac6568a13ed24ba211694cf250cb5a7fdfa458067445e9141c4cad54f419fd711ffced61403eb49a66aa5d8cb7afff86be9b2013f24979d3c1ddb14b7e79621579c4ed1760fcd4c2df6af60f15a751ed72746e9aeff0cfecefffce73cca7a30431c90512896509020b870aedef1f6346b9ad30cb81ea5949b9a4df0d8b184fbfe1260b05104f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4fa38bb9728843bdce84bc58322c73348c0005d2ac898fc7a73868ffc1326d975077ffd2c44839d23e7be3547dff373af9666da9175cfc5e2ec9133d2b519c6c013d19dc2c96bd5d17691622534f7ff9ea2e04e13747091608ca236940ec17c08a27098df8327123be5a8ad24b856b3c24eb780593f9dadcd4441638151857b3bb847002a44d53c89c6213996fa4efc89d3753932c77fa9b3bbb7329e670f91a301b7bed66d6e04422513d7f1fa70f378f6f0b2166f74075e9f1356a31c00f1067cfeaa19a300490b3f143073b79215a1317dc1ba272fe41633a1f33877448201d2c3e52679c8c0d66ef2c0e238b4043437af31669fa50857169c60283a9432c657a5a90aa868f7560c064e9d6f062e456b29effead05794e8027fa2512a00c8df641ee347ef55b641b7e2df24dabd2d9edd3bc6b1aa46d9223a59e72f331d274a117b3502671fc31268b25a022e6d8a959754a6d7669242ae25e3da2e22d8f13f5799912c6b6f5259f21a1a716229ae48fa9ef3c9240adcc50a768a29b113aadca5431cecf351e34826cfdd415d1fb1910fda3b1591634bdac57d90f64b0e85b3a133e3135797ee90fc518427ed8adaaaa13fad4fe108e79052a0aa3a659ed4956e9a8dd621785b9d95a194d60e41994a19ee1eb067e801cfeb7a7846b20bd89bd54226baec68b98c90f394e87c0f251a83abde921fc4f37e8a9de2cfc725eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha0a73296491c80b783916a264e6670f9a8c6d36ef3c74f43b559e86ca31208194fba217f14c094d1fbc3dfedcd0ab521465e4df150fd8d5466e669bf8e367c8a12aedc02e44028c9059fa5dc1e9d7348a79cce5c89eb38fff25551dad319f48858e14f2c0b5da698f685549814305601f4195e909835d515ff14e8d525e12b62cdce99e0623d2e36f52fefdc17956a4467f9a57c4b8e4f772adcd32e382f53c89470a18173e18ec4bc3c6b645d2e2ac53ed9f26ace809166cafd64f7e5724bd350c515a9efd6965d164adf50d99cd64409d8e8918e29a9687675526a9d24bdf89380412ea035cbc9aaac728a013e5fe668ce20370edfe7edf9f5012049c3233c359fdb9cbcaf3df010549cfdf6a166ece2e0c9d87f10b7f4997c835bec14d32a7f1128de2bf6e1af9e4450dd6f8f6fc0161f85a1523a18e2f0a98893821338dc079a36ca732f756dfeeb830d0b27b97ef2cb5ffa08c0e21a4bde6a67ac8cda1058410d7911e7248c4d242452793cc0215ec59cf83fbe732afb99a96a9c0e3aaabe99476f2d193c8515b99f758609347a67cec9ccde8256f27933f9c37dbf8f69df2e472eedbba0624fadbcd92461cd62949f36ac7d9243251992a1dfe38652daefbacd60bbf529976fb68b1768a7d556e9538f5cea9be24f684752721eaf3e3cb4b540cc590974e199d6ff42513c2bb3022deb84a76375f73672f4d3b445b15b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd55359dbad1c38c2ee1a30cdd836e3d9a9b805fcc7af1dff99967fd0d830729287609911a48896e877d0a79d3caa9e8344435a8bd6ad3790f46a3ad111d8b5b9639dc335726ef039307b755c6dbbc0deb4738db27157294fec5ef5a5b55697f9af4a5ec743905ebde8540daaf9f08022f1f2b557343ba1988ec2e33377923731667fe53a3618bb11dc09264c9bcc602e854c33c97da9249315cb399246101726b2ea8c2033b1a47b9aa7b7b8037de903c05edc564cfe03da3df4d1ef1579a35d9f6e7ed7e35b919559430fffd30165ebe4875f42056f7ae8eb7f5c0ab34b974087bdcb804fa78387ad25ad800b30a435986a46907bf905bedbc0ac0167f0413bef969f0e2139dd746a42da6d49da855fe3e7f7af8743cb378208c2a77d09c5753320173976afe4f642c4b768324dcc94345308a21a54e0f4955d6f8195df1c65cfe51c52969ae17069e093126ea215ffa973d19b9a3f8a2662b222ed85ca21b83ae9b59f23e3c05ca12447f1d383ded4a10171ba34a40b474268ccf7a1ea3301679ba7c8aa757cf5ceafd29e100f87802b49257bad8b6b7eacdf4976769c7e439d364d2d0a13f3c4a5257fc6f491ca6a67252ad5e923e9b0fa414b11bb77a10002dd65242ba15bfeafff38165efc1f8d1aec24097d8595a6fc9ab2503db1f9c3c395532b7939bd490ece4dde0f81f3d03109ffcf607f42179fa3d1c2f447d0bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbb01ab8e80fe7164106515ea164feab60429fcf84007e6d89e2bf0491e6a4598a0f6e91ed696ebad08b5297a9dbfffd98bdecedad01e1ae34bff393c6611155c703d45c79c4e3ed8e82700d9cca81156cbad9b3e1cf0faf49cf760495008f86bfe02710f90cc2a3c550397b301ec22ca294eb3c87845c8b962c58b0206da8c109e7c27b67ce9645a1f2987e61f0414d7d4a094bbcf228d21545f4cc9d38fcb1646005bb677a55a9574e85e6fac9e265623146e93c4efbc8406dfb1b3ad4fbed6e17d0216ca117721160b0b6df2f56b82216544972ae7f0311a715ec8ea1ae63efd96be757c39afa88911c6bc9808366ab68abb5ee9b3bb2c4867dbf9238ad4ffb8c78fda082da2aa2512322d770a06f53e1ef675cdbc8376ac9455e7b0f798a95e37542792b79637c33100ff36654abf06ce4fe84b71a5f070f1c2f32c67b5290316ab55b3a34c1e813470820e8c5c7d37ed8f64725d6f68fe1fd4725bfc0e33eff981bc51de385b4f97847586103f9e978fa1bb1d326235f50c3d9986e0163574b1c88667dba7c6e435c915ce53101253417b8a0c79728e0ba8f50c8bd5e2293f839dddfd51ce4ddb7e1ef94bbbd51cd720034007778bbe2b4a3cab20d750f365a0c20df3a4d2f884547864ef510c5029852065cd19f4644a0250595a670d13af77f8935766515b7425c1484e1f05e341530ea3879801c0da68c2a45ccc0c40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2acbb3412eb37f86b728ece154dc4227e09cf9223c6ac75c468e787738ffe92396710659eb86c58abf16b5583b768bdce45c31f3a0d1a7050ab344c5a6f68bb06c963d29fa83036bd409a8e1192fa2e305a6da58eca2b91f125c820f906bc0a9bc8f6683f42b9797ca48f0438197d51add2fb8219ae038e59999ce52f496b039cf951b231293b8b34d8b0b120247fa8a62566899521717c6698f8546f565dcbe8398d3794a02b16e3e31f261e95606a53d80e173d49957da1c152e884ac561eb0b818c7883d072f36496c3c0810c4a7dc5f5ddb881c11673fcd99af49f3533d6cb9acaa226a7551be3633e44af5c9c6371163cb6ddaae517a0ebcbed6c81b639c0691e4798714956f48c4560d80592b98058de4a63639290602015081332dd20335baf8f0f7b8cc83a1724c76ac1ee0b576a6b2594678c59444f5482371d3be759aee5f4b6b6dfdb95bc74f3435a6105ff6300d1aefbeb440140c234b909bbd382bb041e84a2f176b4f7d16dd71edfae4edd2244e3dcdd10e8bfbcde3bbc1a9a318e953db85bf0031e60f9d2a121949b867e12db8b87fa51052f79273527a47f162134707a08dbf1db91d8e20fbcd97221a5712dcf53846556ceb096cf09815813e11f201c372c04c0d5c5a1e330760a3f8155e6a4eb0d21fade51821cbdc61b978fc50caec1df270ee5d0d9e917dbd322ee8dd298531ef2feff6f409098c430;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9ef48a38adb5bc0c1eb0c6a2da614910b68c3f1343656ccdf0a9ec24c05923085eba5aa5312f04e0ecbde9c609848f2c3cb496cd6a2b0dc51f15f28dcbc908b35c7957a8696ab8e5663130f70148aa9e89a407a3eb764f459a7206a6440f36e9f52d9c3afaf098746f396157a19a4264ba7288d782831c67f7ff665388d5b4a33bfecae85efdd600c40b871fb3099553d7207be255b4a0d7a37756a8c9139a19126117d26c4d00562a9e76711aac050b3eaf1e0ae71cdeb19bdedb30135031b41a5bb80bbc96f86929b357d8c26c18610584369e00a553d2f9c72dd079c6095a37667e63e50418f7c145e8e3294291cf6928772e567e0333a037d1dc339520e1c0e3f5aec7a57d3ede555ea7b51f99306634844ebd4343b45b419ab13f588d614648776b186eeeea724a7edac3c92ff80a04131ed0f971b31878b9b3e0b367034d429273740288d952d96e4d410b2127272f6ef0905abc773a3e50212e7255c5348cf9e6f4361845f4583889e164f4193a1851e04b0831ce70a835c24891b5976180a5cfeac3833066d95255ca5a87ba4b35dd279001f1091fa201118e44026a45e982590299180f49ab4af27d606afae2acbc8b8d5a5622afcd7c482543e2d40f02aa6adb5d4a1839b4afc3af780e60fb737c1917fc63af7ab888e1210e4a8ee6c7a17c0f307e9dee900e590d85979c363b6909084f19595d2afb4602373173;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h175f0404006d5b3aace3cc6a5038e67bebbd74bc41b725642615c9ee9022b910903286565f3e232630502325e7e779a11b936953269e8f4df159973d3f65ad76153236d00036b708f0fe67690d2ac7cc921716fae0d4982f0fc0260ffbf2dd2932566cb679584d8aaf3dbe526d3e2aafa8532098bddf95b54819521529cd5d56afa32a90503a6fceacc76df8cf945f3058e4a1223bf893cea4c8ada2f7c1b404628c2d6ac4dc7daa64a0b2fbeb4bfd868522791611833057ce21a6b413bfcb8d8d09d6f7a2068c098d3842368b56eb488b3517a6dd8129ce9de668979b1b02784a586982744077a36e5808ac2382ecbe6a2e5bcb7072a6b473aeecf3075e2021aabdaa91a6695b6b435604468263b73c1a9bb6bcb45c322b654143ffa3e7d5ac0dfe459b30d1276df2aac68bf2e24e983195f1db229fc5ca8b104792722106720254fe98fb9969e0b9bfcd6633daf4e47929ad8a429e74e8deccfd1cdc393c37eccba0aac90ad3c119433e9a4e4a3c2db7d1fe25d451a29c8a98b849d301d949d564266dbb567b1a85e86a4d4afe0a9022a8582179eb19d473b5aa3e79c53a48ada41a2806a9811a7da3e6b7db8ee0281134713b27fb6845a014016e09c0e3d677b494521bfd8e27ce533b99821ca948675f4131c4f467d7704955a3b9067c7a872f2e1b061eccc4f6c1d8b5b3d0287eaa1ab12a42b8b515757d724fd884811f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3bf9e9b4d4744bb701f79e73ecc2c0db34588dc7fc0b21089e603be14378bf8135972a9722b34c84e6ecabcc6f2a5fba09614395e51867c297cad23407ffe83c57882bbe16e5fb8094a0437afe21b55b18fff1568d756c4622e915ea1143f35d183a04ab2223c9b463853af74cda48797ca164e4a33ef18c697f9ad58cd8f7e46696acb6b1db520d7c7ae43b886ad7dedab7b5d809e16e2f5efc3c4abd322b5057e481f91631cc70ff9bfed2e952ef189ca9d7881196d77c7a4a75346478365c5c90c176ddcb493e0bf4af863c41408f56e3e10fad43505ef9140561a721d4c894a049d4ee9ea004b0c2aae9dad57cc0d9ee8f71d1e155ab9c201d1d77b2619e6399b35c8ad090de66c30fad1de60d7fcc044f6e352aab39943ab0d7a327ab01c47d492cb92429a4284c41b46428aff767c9fbfb9eedd9bdea9e7e86a4f2d8b59b6eec6fa3c2309bfefbec20350ab2777fb5a81a8c8bb05b7ceb1a6ae5f5275841313f2a19143701d26a084a6ff644f57c6aee3dd325ebbe2b3dfba9c7f5b91cfa0bf7fca4a57c9a2a5a33e94086231abd1a38de9ffd14f24cda2a113cb539a5ba6a9814f1526f1aa8c82a62dfec402da6cb826b9daf934d21792ef7d9257b92f62ac37c73288aac4f0e66fa13ad8df9e0f7a2ba9959a56bad17ac1d4d4e72c0dcde7c0d75ba36f215b70ae5fe91401633dea953f3fe1179893f44a1f2e31e90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8f4d61093b495ad26f8c252faca57451f6731de8ccbfd9f18015b3aef87f1d5e6c12db3acc3704615cd9af1ad6b5691311a1f2556204a6b20fc7eb66a4692cbe57964219b03381c8baefaa210bf9724bab30bb8b54ef44ae7baf425334cf40166b9e3468531461fa073354795a5380186412966d9b151dab0526a00b6cdb32f6317b3f9fcba9f0d8d42ab6fecfe8b6a6630f4f017a7b3632d192707c1b82c35171d0dc39b322c750b4c230883fc21d36115d55282dfb60e7226e6f56a021f799dd6b57790914e861fadef43637c94c74b116f1c3ab849d57a91b2ac41d458d7622c21ad833ef6187fddc4c8ec38304bad5f220ebac0f7b959b912c2e4054ffd85340daa91643a347d883c672e5026c4f90e3bb36a9df3290e2a45b91941d683069bed9994f45afe5a30fb8d9458a05f97ef38bdecdb33e46e868599c36f1b2ca343411fdc4aeb7de46ff761ce436971222a18671e3153cb8e05424b63bbe7ea09a13478449fefd62e5d8dcba58365026b3683b8ae02acaf24d6b15698f0742c6a0676d8c5f94e7fc3e75acbe939c8fd7bd568537648db5ccf17429060716f28ff8fcd98721211c854c56fa9ea4bf1e406584f10e7c7ea63347eb0db4ca9172c6d255f171dab985aa1e1210a2093b3d0449fe83a989abeeea502e4a64fe203053aecfeead818a68cd4ded186a1a40707c00c9fae0369e10c98863817c2cc67875;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfb2a409479a0b4e780301466ef55aab44bd465f44dc5c397989e6b09473506e4f44b0b5e388001a41bd4fe6abf00b647f0be33862039a087b20b33c1cb6fef29d6d0df8c1cc34fe19e0dbcdf9e0b895056eff6eca69005ff361bc9f819295e7cc7f7488c58e6f1e62959636dc24a0271bf96813dbeee833afa7bc438c6c6d4cf8bddf2ccc20fcfe8766bc92345503f394e4a75a4310c1de4cac3346864aad15374132107dc2f33f61e6b325cd9f8f677fd0afbb0a6392fab511ce555d40957b0f37e4d68af18f82d142cfed7785dd1d603a21e73510ecbc16b163174918d6b26d66f92ca78e7ca4c98d44237147b7c4a3546b25ac11fdc7e8db6bd1b11c7926c4a5ab88ddffdaf396cbb020ca634c86acddcd8be554654dcd7ab866c20e83b3727b1acac0dafe3d13607eff1a61a7ff31e115fa3d2a535992e435c583bcee138e134d65549c8d8a636ce328c1cd7539fca20358a1d46510eb41a1d99a93736c0f44e7d70d16a1051d87ca0e7f2cfc727733ad98a17e3614eecec5d3bb370b3c3ec2fdc31edbdc92b2a6393c1e0e8dba386f7e0e5735c38f393b92c2949e08048a5cc6a137e572cbbd23bfedaeed00f13e4d8aba7a69c845aca9ebfab5533eff9d30e5504f339b54f6c69cccef68d2190291318c3c7ee576686d5ae4398fca7374230bcda9e51ebdabbda597be56e222bbfbb3f30cbc37dca48a02760d5d4c51a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h671711b7f35c14fc54fd1ae0b6da6321519f7a71f6201522c9ffe1d5f59407611eae0d54701e9a131b992c1a6f3c38a814ce9e7c1e99fb66941c197c140edd8f272466ac5015d199ea85fd4427fbc8c072c6ddd23fd49ab07a0227e304ddb6c74b502cf9dcb17e427b419a63dd492f71a75928da03c1410c2b09e7a06df39d19dffa15179b79d9d1f38e0954aabe057b5d0d9807f19fb1586a565aed0f1605d92e9e6d9b1c6aa025e2fed5902f45031d6e0a750ccecf93a7868ab95284af12e53fa57c231115acbb5d640b7536c1a66cdca34ca7567f80181f8fd48698231a9c40659c857296a83bb1cf2bb4758b9d8a4aa8f94295b331297673f7cfd3405433201f310c748aa7c4a596f988f166f7b5c4f675dcba034f27f03b36c4f05471381ba40ab65298b88a78bea8576b5e0b58f3e6d4a22f6aff84339946e5a0ae0c1d3aea7d8737eca36cd633e4b59f02c75b37cac7ad58dfd7e7167987668307fe0935a9d87067f76f61ec481a3d328cc349845e8aa7054a4c1edf3d3b35f02b74906252671563743da8d866f54805e027199410fed08127237f492ea249c996f16138eb1c4b0dabc192df510580a37ec9ac4a0a11c7cd8588cd6b245e59a59a95255663e2ea08fdf9448585ce5b52f7009b1155e5b94359ac62de5936baabc4a289c54f2c0f897f36a9dfc6a53c4ac0ced8b88119d55c4bb24fbded93881417baf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9df022f7cb1f8ce78ace2790395cdfaed6b7a0fc07e0a3df4ce2508045924d76e449a99fa51640b58bdfc2f59827f297ebedaba6b97a04ffd138349bd63661394fbcad6d28487692d46a3feb8009d61230da4cede36a24411a8d8e126e54702a393bb2e5591becdbedaa54ec7bdb7b44cdaf0e8ddbb068fbd0405823089ab4930b2752700fe07eeecff6f14ceafef9497fa5a9afd3bc705521e93e2dfc3f91de7b56c0073cd90b3314c0f52c443f855ba16ece9772294459b9a3b7b1bb6b792556e415ec83d525813a05c061b4b9b268228e9dbc14d7cb26a4ec9163b97bf3e75c0fa09e59939ef4d2953468ca9daf967a74a9bfedf1cc68cfb9d187565e5b066f0bbd3e6671169b59f1a5de25fecb879fa54f166587b3b365dea859d9d3acdd5116d121a67c25edf0a12bc79fefbd9ed3fa5898547d340f579c0b9c666872a2703f9a74913a3e16ee61cadf677e1cb38fef78b34509c028e8decb3a379c3034cea69eda627a44e96b5acb5f65fd2242b5ce6e1b25d70d91eeaafefcc8708be4446a9e35d675d9678f1b8e95990f264756e1cc8e257091ac1492d7ef6d50ef276f32bafeaafaee1cc12e4740bd5e3897eaa92d94a3e794f3c171cceeb0924a16227d4ef7f6d173a808bae569d6f0071ebef6c476f85c1c07994c173dc093e293f93b48427de4b9c3ab3bee4785244ed20813e953c53201070d56b4d0de5439ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbf305dd12c8e4f6354736d67a057368757f955fa77ae04126544324a6257a62691521811dab74bf171c721d35a1da7b648f4dfdcfe2f80aad4fddfd28d41d76035bc7b9aa12a6522bee67ffdec66ab567e0188e0704c1ff668e693d367e83e8e6e6bdda64bb6cd8642f9a0297e91fe1c0a5d0f4c2749311424694f5d4a647c29a3e1795cc6a9e63f05b0d526e116571e06f7d676ee19af1c52c257a8cb798809eaa8f159c542f845e1ae9f6745d8a8d41a6105e7b7406579ebe4f7c443158cc69068ec9237d71ee8abae88b9a333bfaf63b58c32c30bf3d7c15f437a9dbd9e37888f5818f16543d50e2ef07a08be4230a91cdcd783f295e21c203fac6b40a707f0bd2843985a53e56060bc7c309ffc78a26d99adf4a135c031cbaa3c924a739bb573828d60ca42bd00e5d631264f685c797d329af04772031a2c92ad8c7387ac2ab0459a74c6e8b7ed077a91e78a983160d40a40c3d10ddf5b678ec9d95f92615d9eb2a1c1841e95207fad53aa2575aeb8285745df1ea552e4b8db6d5693253b3e3d5851548906fcab2d64f44ca89b531682bfe31e062a6ee567d23118d08f488ebf289522353c206e0e490d3188fad66e8af2730e3e13c3534128170d8f429bd3ceed18ab4cb6699826f53060d64db11b26215041216db68fe4422cd64608a9f4e726005fbfd605a1dc8678de6e5270a96227fe577689763542e9331b2f7c14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb7c443b167db1f9894c6e1bace43f82a7cfa92958e9341ca643b103b05ede79f5a7ab0c7613788f4d57b83ad7a419098be1dc64084c8a68d22deb2ead820fa6767e9c82ec6d512589cd7b81bce71113ed3696fabf166be4842e821fb1f8cbcc9fe819cf4c92a0b0d81040de51888e493c74f51f6e351684461bfb83d000060015d8f2d6cb43f5ec85ef5f920107d17940f6add5dc4b6d72d80a2725b2eef4d9f7a2bc6dbd90fdbed4bf4d0fd27e9858257aa837c4e7cb6380b703e3122d2243cb56d862c1db1f2eeb9a423dc5fdd074cd57605ea3a4ef82fc1471769b29f8b4d3b06ab51c79a1cd3d41bf409e5b16bfe2f73e708f818450da6fc5b064b8316654ad2353a1cf7f210cc6ee62996e412766bdcd4463793664d679cd481e3a2ca969dc0eeeed87f38d494e70550342d378d721d020dfaf973f5e62393245b5dfe28f3f3a547982a9acf07c725d31a5bd94e39168ce6ebdbfe9b933ef960f26fb3067de1568d3acef77dcb3eae466eee6af6f283200914eb159bcc64959d87c94591e349c74442e3c0edfa34185f83a6614418a94563ca130196becf17aad66c955fb6777650a6bc2c7d884c1b5101d659bcf19f597ca9cb836d3004bd00a75776d2e859c2bfda5bc3f51d8f6c9119764f22f47f0894c86f2d0cd2dbd1200f0d8adfb32a20c0d75093d5a646d081525c198becd784b4ead9e5b2f208af57642e6517;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha58ea12a2f24bcb2d2ac475fb9095a300e3207b1efc501dcf78f6566e63c5e97ce6cee5c74f9eba9cfa3ee026c81435a363fce331b4befa06e706175819bd4ef3b8adc239bbcf245a600328ac7a1ca94773e4b0ec7725992fcdf318a34ba3ec650dfc664fe7b9eca10f3f87b27f7fa5e8e8332def9169f361e61f910a662ad37820b018389677944340324472bc5f6405cb41e12bb74e9ea47c8109eee2cf66bb6404d29bece85e68ca8c4b5ecec596981bc5c881a43dccdf0418b14d7deaf505ae39561fbee9591443337daba4ac662b07f3a8aea8e0998f464486e1c9d028cd005d1ca4e46677e6b298f65877dd672071b1f920b9ae7249d24c6bac472f41163cbc56bef3a10e299b0f2a0f37dd099e6db1e34c9b7c7b6dc24178a3f61953a6b6c3158c1c94a0ddd49243a3c3e02c4485f13ddedeb010bf6035576a6c1b6a5428e7e2e06618919e833aefaba97476b806cc1d8008fac20f42587f1290c5c79dc87b7129b402dd26edb450dc8b22e51af7c8534742f9f6890e1529152aa89b600caa12e7b77091126ea6f0c1034417bd1dc12fb806fcfc135aa2764e79888b3a5551cb94b271c859b8a94ea7f6a39f7ad9ae81282a7fc2f6f57b4f9cad20de575fd04573c327a7087d3156d120c14ddb33485c6fc5469378fcee22bd4e095cb951c2721bdeb10ec9e95bdd97d5f547fd9c7747991ea0414320c1d39087d382;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5d920eb9fff20d32be2e2ba5c883fe8f6260118468866bc226f57bbe972e637f0cebb04e3b9d6588782edb044cafc353a1f12c5d79b03c16bc21c9e298dd4bbd0cb75b9308efdc8125648f5031a50800bd3996039925b17a6fa267e44b498a7c7e9f217d93ae7291e088233c56ab182cce6fa30b93c3371af57a40d436787ae3caf90266632ab6f21879d4c3bb1029f2e36376c4ff9779e1595aa02209bb863d0b53034b1dd42ab68f41e9df40ccb5eba5057e62f54a0fb2f7acf36939570c2b3c30b732abb96facc7d79776c92639208db2cd32e06c99f1939528cd3c7665261a653a575bda2c54c15fc7f4e82629e67091a6da70f3a04d60581dfe204cf54732584ba039c963140f4b22bfae6dab4717522c187a0846056ae6c2faea513bb64ed67b5a1dc4846cad7ede8d9e817579d48a3bbbaf3ed711a2633ea9dd6571b363af59db5c6f20e718b4822c01767417107065f99a406c964037263dddadcab2ac69c771dfe979ce029bed14efc731ccd269f3bce5fbf21299b421a8922b6fc9ed3376df8a81d6ed9910da8ece73361ae68cc26e4b2b4298d36a26e85362064f02f0fa2b43a9b9c658bcad8780f840c6d93457b6fd6f2163d3464d050f7133b63ee4ebd10012752b6be9b61231b20432c3322cb8e105f0d831475ed13249d451c658200c4663329e7bcf291db5c8b30d17698a0ef04dd53f8e9e48c3b513d138;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h928172d1374aa750565272042da1d5f994cdac54be1523bf7ac22e465590bf9bcef9a76fbe4e1ac65252239ec8c1dcad45fcfc972abf0092a8de76a26d1748ff112607b2601eb9d2ba642a22121c5df9cb381c84bfb165a82a53dcce60df9680666c1bc7bc0831e27ed8f65ab7f1dbfb75afcceec6ec9da83052ab862f65eeb2c47336a08a61a2a324275aaffa3970709fc459badb44b9e2b7c6b22edc43d13589c184a0f05f35ee282abf4fce24d44dd71fba156d7a76587f68ebbbe8b68edf7135b2dedb5ea5882d8d9d4c714369df7b0503e5bfdc5543a336a9942e8fcbae718088685174d503fd7c8a133fddad02d96969553454b086f63d2bf3737ae513f03e2da51d39dc3aaf3c9ca5d7948097c8f6ccbfdd35a31c18bb06b9418196ad8c9ecde0a10f552fb53ef76493d6542b1eac293d30fdaeaa43f8d6d8203e476c00d38e5da32013c2f21ff207f25645aaec76a123c3a85002d8d2d11d975c99df093a5f7fba046ea1f85c0cc3f822b25d1db1887dc6c84678b20855500a7dd880b8887048ae3bb7cc10469eb4974d655c2aae8e9eb65955c5bf275fa57bbac8fdece31fe2e9766a9191e6b1d091d2549aaffd66dea67f1838a3fd6bcf997bc690e30357e1681d588e6bac8fb1d2b05e2d39e47b83348b243d2a77b2fb155f6c648adf39f0a0f78337d555cdc6ace5ff7eea4c5ec82a6e296368980be6fa24c655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6910aee08c505dc90ef71668ef7f33b2720d9db5a41db0728b9cce00e4e69f4d502f2ea629ea22b35cd7c7660a6d43c1e5a0a29f5cb1fb266fc7b778fe18e35636f5bc1bb90ac29cae7aa4003351154d310b9c09a64ef5b1ba483fba281ba4621d014700d0c6c1f5159cc966c0d37ae2545fe7fb38a40f314434bbeae9b4ba934348cd8ce703199a8825c4033acdb26a38eba7fa739d7b656ef63c5a48980be90ae4d4c5420c63adcf922cc96c53074552c841f0649f6cfb9c648036ddbadd8c8ee8810b62fcede43f7fc3ebd7f87789a14ce35e0cb2fd3c9b0d87133c9030f68349d7f257e60a6e4f4870c199fd8689b42f309c60ac9fae83c92f9da83d81fe93e611ac7bdbe9850296700d97590134dfdb132b0f1cd8de23633eee0580d3862c5e8e346c02c852a3e1174df074aadb2c0d6e49d3ec72ef2c9cf66bc0fa7ab20d4af5ac27f0913fbe516452ea443fd518fe8a5ff3b9013a9c15893b52d19004aae6a1f9d72d4b93ddd11e8445c276fac2f0d552ccc9ffe8f7c9802fa84ccc4f69987eac0e3cf58b6597f974bbc3cc770f98fd7677bdf0956483e69aa69715a10a97f2a4f40b0315c192a3ffb9f6d82ccb5d488de312988b39638b52c32a964b736bf4408dd535f33b051c2664239388c568992319509415bc54baadbfdcb83d98fa9d6aee0e237c0181e848bc3ff1496440cf7943ba499b1266a631d328fe23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1bb1818db9cf04df51d3a9e1a514e88f5671c84daa69562eded679bf99baef0a1d339c0bc3a759293301a03be254d64fd0667f4902787315f17c40789402205078f356b8c8d5b3f3785d724a41a79b3ec1c26e11987639574a94f4cfcd9d3e7904a716544d0082980f59436d24ee2b1e7ac539e857321134f80fe9170ce455d6b8749653f992eebf45f540dbdfbe98d6084952dc5c096b6d175a88dab3cd78ce192edd74ca475a070e7f2e8bec533cc92b499208389c746660c2daf55ffb54f323b9a895b463038f8fbd195db83ad646333ef1b690ca9dc2bdc7670703b4ed89a7abf74227c5c88082fe9a0659a274832b4b1f8476e881aa03bef68752d664676bd71a285e4ffce44517135ec4035cf8c065339235588fd3b916dc1a1df4e52429489c4028bb21521e280e25b1de78d180f1bb9258cffa68b686fb9149c1943d841faf8e770836bf50cbb46cf08fc5ddf66793fb3e825b5137cf8ccb211f531e341cad6c530537011c04c0c6597ce1c74fab3aeb997d2fa5f1fdc576027d88a9146b9ff2b77313497cc428907020a59c2819e813355f81ffec6034ad707ee8fadae2aef66378e82ce72158ecdd59cddd7e1588ff6a7b3151aed453f9f7587376c90e52db828621cfcb9509b8d0503a7f1b9ecd103fc079ef7e9578c9e777d40337be80b3811083c10a52c58ae729f1ce811ca7cd371bede0c6c4e973427870df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e5406d9a4fede8e66a328363bfa2503fda66d3a106df9b878a02195021bfcd49f3ad095b7e2652b5c3a095adc62ceeb6a543cff6a663a655ac8a36f25a6e0410cb319306d1e0f8a257cfcd10759c64b12451d0f396722b0dd27be0480f5293b202c5ffd32d018e28af426ad29fa255a003835c169b36233dd206ef786807fe7e51239f81f7305da55c632b6b533caf90c32497e7ad0f62a5d67114e07408da4f1ee7589e844f4e8e07bf3e59eca08f7dadb92420e21858b60f50d05eeec2a0ed4e701e154a9a24b9fb8115685af9afa90576d8a9a780f666c6aab510b0ddf6e84a7b9e8f865a5b70f667e18aea4b5f2c4fcc337e9eb48ece82ff313b605efe1ec86a62e93b8b8c90884145f2a8e176277f4b8a87a6a4967f52a6a40c68ac77d51ee106154d9a9e41e36ddd3a7da900aa26eb99447a3f1b74ea513ea503bc94b983b215745e59d4f31cb96ebf37aea4ed0a43f5bb0f81a51ef9a95234e4078f5d39accc94a955a08476fe9b083d8346fe5d24691884ca4ba54e9f112dad42b8af43e94984df240979d3635bcd6ed4259771eda21d1869d531a88b7f71408e0a4a58fef2a11c37cfc8088b757892241b00d4924a199fa9569a084cf890f01130f53d3291c555323414d26a8c35a99d0ab21dfd544e60fa3b4f18c5595510663a70eed6f55ce4a205850f25ec88a4817074ffa62576551ddc1715e22fb2c763624;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h48af2fb5acfdb4382985b60656f364d1e671a95997284258699648d27d8a89ea601be41216f2be51de44a13c05355531b87a956e9cfe72962700ce2092eebf23f802c63f1cbf65abc1999c16ab02246fffe30751d95d54d51003ce140bbd93e832c4b04e76d402c72e753ad133199f8de22a282114fc4e6e97ba8651d4b25f2c833dead092e42c16fc750ecfc5c25f1b55661a04de7a1f412d623769925efde6829746adc74e254d345537fe36eb0291c4060dd3bc7bca1e48ea587b189282c0dd431da225c512967cad4e222758cb9e72f7b1d5c4a14ec2debed620eb8abbc29cc4a8eeb6ff9d785a960e1a61d9f76c08429c5e1568324d8f671ea0576f9b1bfb933a51021103f4b64478368f65f6382fc4de4b5059453e7b99cec14582cbfdbeb5bc6e4fc57fe10c9fb3888b5dca60212683569a696140c65a0afdb104c7b89e394bfe07af075a267ed8c6bb23bc09eb326704532a2ad522e1c9b41b9d7743c41841ec5f83fdfc47c8b2b42fbc1531c6a5b9071adbf6c5f1aef4554be7e2dd1bb15b611a6801d1b3b38a378f4a3dcd2cdb979134e2f5d4df030a7c8938fd0ba5eb902935b12b6b2dbcf8b4ead26d1acacc3ff79a6a19d16ca349d4e9aa21326dd9d901d0c647db13a0f8fcd6d8279bb86788246fd1e561bd259f6a755d9f9cd88ea2f48c8770d3de20af32a532f74d41f6ecc55fb85407b2d6da9a7e26c727;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he9722abdd3dd80b253ec51a9d485e74990351024a241a7ac06c751a6dd27aa5551ee58b5ef583819f8ae9e9a3e63c8fcf0ad44d91eb0af74b5219ea80456de31562675597ad1acb447b7ee5b9795a694a7c9617cf69b01052734f7036bc90b9ee9ecc9960b91b9f12d635d6eb347b2f7de30126ea2f8d92c1c1b11d352c5173570e615bd64c39fa92e9f36c92c07b8e77fa51bd4e2e3c1d6d926aafe8565a725a0a1b3f8b96a78aac23e2c3fad92b05a2b30b58d2db26af4420284f1841345b2b66309889eb7f4aceccc6d0d7acbf492a098e8d1837b2ef6c49fe4760d779714499cb8bb1bb8ec43562e4fd247936940e31f7c414b8ea3108ee973bb22865efe266066d532d0024e574323e57b26175e73e37abbb05719731d8d76e934dbf37d773ab12d7702e250091d405a8befbdfb7deb40741479016ab29960db2eeac03a580d1a343bb1ae6232ecbdb7784827dd40ee7e3d04eba2fd33e39c342985299e77bdf14161c69f11ff1ddb03ab9d935e70887d35cd4f1f7640d43d02b19ffb3e89e03050634ca6e175376e6996bee7d306f5e14733006c270b89813d80cba9bb0d6be1f71fc10fa803c1673ea51c28c160c7b340dd5d96f00bdab130a2d8a51cec70d3c3b2698a6c71e521b20fba6ab9c6b985960b5e6e8a6fd769f338300294caa405c097d791d855dc61b710f5706d07b1b1673084ec6cc38602faa4c2d59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h61a596dec8056d1be7b9afc623493ffae0a1660ccab07f315f54dcc83121e823c8d1eef4f3d6299fc0a150508486118dfe5ec28dc2ca7e8f324e229ce7655cf01d2654de68ba42b71f174115230a7faf05c95e328a9ed298da1551295808bbd464a8ad0f1a24f844f944f2f53fe2920df0df0df5c6f407865ef137c389e780e6fcde277bf46740c97c100182a7ef60abc5ca5126ea160d7a624c8b83b497591c223aae2e5f75c2710a6737fae687f59fba618a673e50b3abee3fee9504999dabe926d318dcdfd342620110da3ca9c60df33134b799531415dc07bff244ba1704038ae182e84164ffb678d1425abb22befcfc5e23e917f7fb88c82bd6184e6d5f04456a3c9cda4d22f53416433b2d1fc0cda844976e8832578760b47096f4401a1e7e68c7eb6aef5a8ceb73299bcd1b07cb46b2d911f74f3066ad92edeffb7602bae4ac071633a2bbb869aa6157031e6aea6a2067384e4372a5e07a18f26f54649ac3e01decbf1ecbcaaf93eb4751ee35e629f867763ae9eecdbc8d1dfaec0e43b5868f0e9e89b3e0c7878731217c6b9663567c1d2bae482ab453eba1b1027b9017bfbbe8fd4c13f2eaaa3a91c3fb7143e9269cace89698ab2d01a35e309713daed46158cdd32d048f4a0459f7d9065079454fad5abb8db695bec29a352a02b4ed3efbbdabbc70fd919ecf1d5fdfa1ee817a85862d4587242e6c65d6abee0abc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdc25196c7f236671515e4cd42f7b8782a8b2753ec2c654dca58b292f200519e5aa503da0096514f45ed6518b7237f7785efc289b58155344a3937f5c12732eaba53edb3bdf4ae86c0e76ee1ea6333b1488d6baf8e5eecf524a98f33e140c4d34d88a5a067daffbd10586e641a2d429f24c775043351161c3711221414feef6156e64eb29bdc575805fed1f759fd0fcfa864eebfaa4e13a91be9f1e7d9c2d66a4994be449d1a64a09341adb49b8f39696a6d16c8cf24c21ebd61c5bc2f069b7b2fdea798e4f9d444ef607ae5a46ce7e0e04d32c74b6e791abfde5efc81b838d73b32aee2892b72e123671d59941a489c0d72985551c22013b0c5c5f70125d348de9fce59cb5faf94ff7ad4f713bbe4fccd849bcefa5e69874846978c98fdcbcc1503620bbde13472256e802f5b5d7fb3084e78a9b495ed1ebc91ec75891a882d3c51a3d6a61edc4ad465b91564653df93cf50e40250c6fd8d610e396073c69b6eeb7be8f033cd2faadabc1d69280b6b01e2414e290438d162ca7fe13a2a2b298992c5a8006a7a122e4d0e16c4302815ca33fa34b04c093a7c785f97be8ae8d48a54671e065d194218016f1e1a662bb642d69bec34402075231607388587a5ed8364e82111f194e0b97bcb75ae0951fd807b05d970c06ff48c7ca07d2af16540993bc1e45fdefed439480fc49b06a284a44bcbbeaa7134f0e5dc8b9ff049666f82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4d8654b1eb4574b3748a9f40cb6a5a93189b036a36692751cce479537769e6c77d122153a2ad793d7c643c81ad5d6be4d87e0ff7342f9eca37d035ef4cdaaf377af03aa0c8b34aedf9e9807fd5eda33bc670164905f70ca7f7e888f34f8a12b5783ce091bdf0e2ce5643716883507a6d2063271d65025b7b4d53fb0121a2b6769700b5b93a5eb886fab4d77915277613be46b8eb0caa21eacd608a7462f7df5bd9213865cc8f209c564c1939e5474a7fc5eacaa1c67fda936089fe39229c91d2845baacef26924d8167739d725d7dfdabcee6b52461e68c8c5ab64ab414ff1bc6fb972490f4071ee1eb276a9696faf1f3f9a9f16847e5a5af56912f555ea760a3a8cca4ebe7982b3cc1f952d383558d1d6f71197ca803163da50ecc154c9c52bf3020b7908a17b8ad9531b65aff432b7d99de2bdb23d8b4a26d79c51ced0abfb69d690a07c256cbee8785f74d921a2f8e2657f1d583567ce910a0d2f892da4f8a64e61c3e1024f759674366706e3c353e2529e2fa8504d5f9ae29e3053e04075f0a9fbd8f8d9e18f9ee31ff4870b46993e1d43da52d61eff49e2557a6ce3bffb310910ce27d216af2546b8d5846383e7cf2eebed981134f958dd0e1c6202e26188f194b7003e5f31d459580ed0d3b094259d6b5b8542c4264e28bf37fb555c0439883ebe92b9469feb800a3bdc933b99e7d4353655666531481424d05d53fd34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h240d50b84b0b0560988b829d651ab8a6747afa2f3541b4d035a053a01a412c2d05668c09ad1a7082ba0da0f30b96b8cdd27821e8a92979b8170301a1bc45876964524f8fed2766a279d7e8fc6cd3eda81a7031bb95d14845165a3065936b83713795f81fb7dbbe632b5fc244f42b3dbdb289304100195adc8e619a2a4a4e47147662143fc0237098c33e6a81dac5a5fba7074b15ce3776d77451f64fa251145af26686322c95bf668a73006b149a8dab5b2a84b47476fb4447689bc47880f7a4f00824b2d98c055e37d3011be74c74839e2e93a782f762e1543edf5db49738860ac9516bfd7c39b889f0bb6d3b8353aeb43b07107ab9ff08c49711ec06a57fee3e02d8fd1923fccc0a5c487e80b71a1b89e96dd9d610254d9f41181ffc4ad3a78c8132eeedc05a0bcda576c962bed4ccd47e59f98fecf10b7854b63fffc998b6d34b110256ae03ed75ff21f4cad56493895684d3e1bc305ccc5c25cbd84ecc03f937e44bf8df713ee8e4440620d0b7a6faac6c62684354048e1f6b59ff12aa95908e9e17cf5b544df5d38e19afa5fe20f0c8251bc5b38765bbc447002ac26d446882460a1386031ef0eca148661d874346b624a7aa4166e26ea540030e1877a139ee81ead278fef9a19bc79e594f12369ada3b958a345953a9372da6f1999c4e3ee858df25bd020f1a1d4cab671e66b229aed73767f2c33825f4c92c8e7ce36f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h745c099ee3266549d50fa3761aacba691dfb4573bc73a974194f0117caf4d5ec3fd4cd253a833ffc0dcb04bacc494ee17ea21f2b4da39bd8e950a5864e64c3fbc763dda6ec04fd486d4a582571a7875ef87253daebc4eae8e0e2708f0a7637b92ae98382f32d4563b27a82995a027a83d3e6212fbf13f088bd37fde31c41402c8ba90e5fdde476b697e1586848df7acfb848f759c34651373501efb7b0c0b2fb7b8b84149f6b5328068b0b6f4414cad5413e910af14e449218cc88f9a6c32b25525adda978764799b656b41b0850ea11f63ec18e1689cff729c70e6c4b3bda477f18fc4e5b1be6c650ee163078cc4a42f004b0ada31a326104cd85f9b5244079bd3a22825ecba4800800f0397a1912c4f01e6ec2ee3361f8d70c6714fddaf9d0a6f2f1b8ae53d9269cf43125270dd0a171f13a3eebc358ed9167ada468b56fcb73b10364231f84c238c5b29ac4ba50475404bc6b2f41e78ec12d5867251b319fb27c904d8a3eb963a04c0c5c385d19728cacf94bdca9cf9aa59f95b463b8cd6a8a6c9cc0ba63e9cc83c0181d2a6ed8b4717ac2d57a202d203eed754cfc1c37f89151a88b6f59c09ddd71a52fb9f889b84306d2ed7b842ed979a47b2836d7b071686aba6c8ebeb5052e37e13055f8fce9ba784af68fad031eb8838cc485574711fa84bb7cfc13141dc389b7c4d3771754a0b6f25e78f53da78724b2e15bf80d48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h55f123ed02e8b1f7c5dbf27ba53d915e6be7152f20f42bc6e368085f6a692958cf6201876c7a9c13b4da592bd58991efe1f2dfca7458925043884dae38f015be029ab35f7d9760c5e59986a4431fa5c21c327b104dedb6ab9e49a939f63a80e05f43fc545dd888e4522a05aca09e470d354990b06e531308debf00d6b8f822b5b72805866e4af4772bb60792be6cf43681524bb8980f8a4ed216119366a0a211a5d3332344821881f3cbd2e2ed301ceb0b67b0ad9cdf18c7793594e0924a17fc56815d95fedc5ddc2292b018a5a89c387055d82f864be6e370558804ac7add6eec78435c0c3d4025015aae21fd94de9a2180c2bab785653c36c2e4dadd03dfea0d27b91a370c550d9cfc66ea74c470fc90f1475e0c70d011a4ecd3559bfd20a80392fab33a2e339856e3d41cd3faf8dcbb2bacabf62dcf3f42f33a73a03800e73331d9c38ddfe412f59e74536e157e2f005614571b39ba229a6c9524668090b775f436e8ba4667bd77e00655292cd7c6398299e4698552e77701276cd008ed9ff16ba0f9e0b09630660c1e655e01c7e794c1ccb61480ff5987beb763379d21f881a06da69cef0232a31633653a9bc0c5c7dd3e1c42b556c9370c480d07229dd3c259c9eedaf3a6eb82c0cb0de164d256d63d70dcc173a63f4d9c618e7e0e00cd13cc1239a89a1c4dfe54bb9ef80df1c62217467d69b9b1556b0f60019fc4378e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e2ff736a91e720aebc7b0281f7e1a4d434ada706db5da53dbf18404522cebfdf771c8334c17e63cd64f31ba1f4fd1b0eb30cff39ce5ec16a79537e1e9913289c6507af18fc24a7fd38b2f2da360b0a2b147e7919cd1709d2df086de656060f8d3b94138d8b21c40b14ad0bbf113a80608867d4e54090641367bc3ad2adf60c4ef5f84eb37254e99ced309d7a98825841f7a4b1ca864d2a0b723e4ce6a940b86f49e94675b3ebc9c20e0dee6b883c607650e05755d6a044abbe1664e416dfa613ce6901089691003fbaec8165658f0675b14d60574082de32ee0fbc50361ba5d5b0360bc7fb742a7ca2f0c82ec8e50ec8c8a7f9ab37b6109cc016a1edc8d20c75501a357cdefae4b1e1c8895fdcd13f3ebdcd635075d31034f9a8807db9f8d2711889274ac73b7a4ac8e5f923a16dd9694a9be3a12964c19928d3f289bc9a13d3585928bff1fad150de5f3ed9bdfaed734a84a7fe14c22a132493955eb629ed8d4214b16b551c6f1481a1ce8d1a8e6941a4e8069d778a7aedaadf22f5a83e08e4869554d714103747487aa560e0b35986b38955693be896a16ece5046104f8b54d33b0da0c47b56f5a80a841c9ab98d29a36ea57e0626bdf30c71d12d643f212087502eeb6378ab9db736a52f7e08bb091d90975f7ce65edd8f73a79513a1d9fb11ec59d4a22b38199cd4a63aa7c93168451012a16cd71e50a0428c08045e28d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h50ae9a6dd93b47a084d94a1865700c5d3a890303e1d39d9b9f108d1ad4b4a5aa443928372e4b67de1793301d037b4b1d181034259846b25fb9e2ef6dfd7dec31e9344c5c389ff92f316a55de2987b794989cec2e5c2b21cbb18f1af4dd1bd88f88687d19f378ebb6cd259331edcb415907bd2c458613e4f01ac11af435d5395fbecf56355be5a7ffed0904ef132bbc842c8dca940bb563618de266320295265a66d338b4bd8cc8bc1f83089bb72efc5dd3d1d386803f5755db23575c137c794c0cc2a452741bc7bf98ab9b4a0e0b46fc9571028f843b297ae91f57328203734492e18272f0592dec084d396f4e51313c9b26f53a79df3a4a0968ff589819c2ecf5b1b54025df7bc147cf4c3b12c6ebf7268345e496d3280438651ff7ebe4447ca5a0dd46963ed54e1b674d8f3b0f6f0a84188e72fd2e37957f192c8dcac01dd207535030dbb016ecff575968536e04a441be488c7c3870e0c105569e658f432f3bbb8f6f8eaa7d8d663acd8658f0c09f5c4d9b68a21a1d5fe2ef0f3d44f17a19af0f9d8f4d4aaa33e8b73e89c6a71730f7741e4be0e861aead5a204067fd208e6fde6813c56d925f1c54cdffcb6af1faf1afea0e087092df6481bb35ae4773fd20374128c020375cfd31dc9cddd79f159dbfd90349e1e3da6100f8365a1430c1555573700ecf17d39f3c3c04dd8fed5df6f0db1013db0e214ae7bfb9da831bd1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2c10d051cc23caa40d379ae9af98f45c2e3d6a54a2efb176de5ab999fc1aa49c5b1a5da223afc8eb89ee07ef6c8eaad488da0b4debd9597f8d359cd4eb725f4d11bb8455417a2342c31577f47884626230b7d9a45a683f5cdf4f70f2bf3497977eacac7a34db7b128658d6b4ed454b16e0d91dfb8bd1caa6efac823aea042fd0d3bbe50cf3bcd0c1ceaceca968ea2aa9d90c3a8e0d0bdd79c5dbacf56f36dc394840cae3617acb917ca49ba0d039b3627253dee594f78d5fba303a72cda45cd6f34e9ecc09bfb4d658fe140672e17cf7fcc79cf299cb15a2c15df7840cd99e0f1de25f64a43501a8c675151568b17d27eb4b8f12c3769704541598d42172a4536578bd406a188b747986657c20bafbf89a3502ac79104d4cc4f22fe234309f39473c79a8f75b98be6b91b233d314c3f84d037020bc2df55c7ae161cfc48df940b927f8d511cefb11e334c40a4ca6f2fb7b63f69cb3fdd4ed1bba9674ce6c0c8e11fcddf3fb3c80f2828326f3edab5fb170d138f0a18e30223deb55a904da2355e4c3ff1fc42fd2eb3af289b8425786f8fdf2a57f5c5677c757c32362732f7d8dfffc7ee8d0049fa747deee5ea899157d8fe80bc66ee94ab15334d9ba0d21bee63be382926ee116c03ec94a95e4448ee44ea15270f42d4db6b121d0f9ef620d43eb4471e3a87ef80ff58513385a7234cfa0ed19bec5eef6002ac950d15d5aa6dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h99306023837f96fba0d746d33c39bbf6631f951cce285528ab24c268855b106d13aa7af84011f89e7fc5d7f3403d1fa4bf14500e49f14e293b04c9776acbf2ae46c46a3c58053c2c6ef3a108d453556cd419f9591b875af7b7072cb29c3bdcf8f0c192af42d2caaf417e06f84f6f4cd4e9cbac5acc1e6bed80ab2fac952289c84cd37d94b11c946fed4c30093bc61573c29b3fa65a850477e075ad261658eb7fedddf85aa132733e6b6abf5e9bf2b23593207f131a8315cbd1c8a6979a19ae97f3438acbe660ca4066eec776979d9be92d770f296f912bf67a132122cad643048b748ecaa500adae2156ebc18c09e9cec4d5a34a6d00c3d1c474689595bbc531afb669e3a1f04dc23baaa7d7b8cbd9341ebb7f7dcd99e3527cd2b091ddf51f88325a9a17eb333b9eb1efc6397a58661c2921935a7735ce28201259367e8c51d459d6737e063491d2148d11b07f1b5c72bda80b2b0954b3f5446eab3680049b2cfd8d8e7a43144c1fdaee286b7a37c5b8acd26bbed9cb7d9b4c37bf0c0278f2fbb82fd56fabc019a9b97ced20ae0f66d4334985c582c4e822fb821e6b4eee7d6720f9442cfc927b6e9e7389bd1f9f4fe562c2d1382f2e19cb1a15796dfde3030ac06b548c3445916347a1fe1cb117f1651b83dd58b581b7785ef08b61fb533812fe4ace8fafc4fb43154c93fa0023cd0f0fc38926707e98562c423752dfe87372;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h473f2bec28d2158ec71e15ba6f77331f646bbad0b9270965164fd71b3d5f1193083c324316b66ea7daf2d6bbdbd6b3d731b1f66504a23d3772559d8eb0bd0255bb95dd9594edb0cd6927bb133491b25c8cd77ba6df4409c833c9602d31745417fb45b96e55eb5ba2263f7b9bf9efe839155c9366862afa7169a07779c5832848c5495f75f979485b5a2926148e88bd4dc97e9312ca58081dd1125ff4a2700cc5cff589c12d473a49c66c462d8e8ef7f7997194c40bd6b036ec261884f8999a786e954a57716336414ae05a9f62c0029d0e2326cbc1582dcb50d0b9a7603d6af6e5e5af7231060a5bc6462cace94350e9a2fc271d2536aa6076932f3b52d64b47fe120e06fc937a64cd87c6aa8ff927ae7d254c32b1046ee8e32f99475bb2de4f3d080ef8db61ee6402632e66476752626d94ab91b7aa0881f77c0f2774e40fa520616186b6dd8452f385f1468b9f38053c9596b9fa68750b5d4ce8140d0c98523903eea9e6202526e88a44cb3a4dee47cf200f0f9f9a399722e7b226cfbbb908df36e06a62355a9233856eb072923e510eae8ab962ea45fedc24e2b85be1ae37378eee91ab5f3eddabd3b89c890905ad03e2257bba7b1f49aef708cdf6336b103f3f573625d38b5dced330be21d666fabc58c91dcf564091d2084c79c5b7d8dd5fb6fb3f9552daa3063b6e3ea636e49435333800872ef3b7fc3c531772e3ce8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9d3467e78fa44b7a59161678f515cef540ae38fc6b857a757fba194a578ff8e2492e3a919d8d5b6482cc58225a85e78bb29ec7d22d91bbe4d7d6231cb6571bdcc30d2963b7678522118fbcb5546f1d19f5879d6bbdd5b10a3816a207a3c4bd92d582318ee5b1d1ede08ec0c56e9871eab974ddd52f6daaca231f593b528189a5d0bfed29f959ef0ad1f0f8a708362f29c37b12387817a9f32e5edf522ccb80fac53fc2cec629877e80b2e04a4b0463e883808274c4ddc2c1af549fa7138e116eb653745e6b97fb234a3553a0f36bdbf30927a3720bfc29fc6c674b591349cf27e7db74f111d66e8f4cf46864c638a330179c7970b88fcd8d70f500dcfbd276fc1a6e8be31cecefa73d8bebfdffb5718db3f316f4e6da280f2866f0388ff9ad97f82f5ceabab4a62498cde0076e74e57689d65b4cb9110062b4b96a957fc5ba7e8442cbb7a2f0d9cf40873f35a859b00b689e39bb6703abef26596330eae7386955d418c2afde10e91d060f93b6bc1d9cd57567079d522bc959773a38b09d75855bf7a396f2b829c15045cfb21e4d6507954f5bd6f105d2fca4ba307f98d8378c02e8b351b30937c317dda7b433ebf2799555a69122bf53381fb195f074ff72725470d6fdf53a463180501542da3ce1bfe2e6896b6aa0ec745a2247bf568b04f2fb5d5c621175edb82a8a9e3df6ec9dffbcf871441b9089ca0bf5c8e9b83ebc63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h431e80ff4ed83e0bdb3ec1dbc7fa58f5c4fe459f24b36976d87d46848b87066b1bd0d12e16ea57462b1458685fe583b7a14f9f5c4d860cdfe49346d1cb64a862c9fb8c8f0d1b4131a7fdfb09e17b77b0f1bacac58e86db6a70408ea0fac6531cff7581dbcf97709e2c9eb65a672a381e7e182de914e5e9dc18bb307e3bd104d344a9f3f0a3cc802edfdfc3fa0303a0e7af5609e9e72b066cdb280289a2504e758adbd9c433d5c5811755ade5a6cae7486de4ca55873e9a52e07b8e6abd66db692417479d0ff1eea2b0d1b311f7a28aef9ef6863d28ae61a98a97150c6c37b0024990d9fb2c0a32abf5620e3621f26c63f1c2de89e1677d6db2ad823d96817e6167984e7c34d6b36c7373a5dac4ce960342b3563301cbbae29484f38e5c537d102dfe68d6fba1391fef7a9d8e5b3c5a5ffa0aaeef95c087a181959a274c23c604639a513257425fe717dacd449ee33dbfd98cc3c848ce33aa9d029e0a5e8a6d53bfdee1c66ddce51abafa64330c808171e9a55bb9d0eaf8a15c545f1f0feae8fef63fae61accc1ada26af48c08730dc9879572cffb3a57f7d67332b22759d253603bcb450c0da98b943c0f39b656e5c9ce772675df8579c21bb8dc295d0fbc1b89a34f4f3f1ccb38e0e074908f2f915e438521d7d7f0f3ac1f373555cf4455c8dddf922daf396b9f20e5597f1e6d1132e1ce4eddb7dd4d068e480ad2309069fe6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha288964860835596746812f2fd58a0cc04582057df22e36009e6f6b90e2831675bead20975c174deadb8eec89d141563be441f4f0cff9fea609d67ebf74cfda1d8cfe8d124db13d16966d26e38c2cb38e1cd01c5677615d0a860d0f8a7d64f85180d2c9a879e049e76d3c6d568650aca3742e276274f6ba8e73fdd109400bf0ef00b038c4615900c6deb526ed95c4ff1ac556e94f90107e99352de36b86928786e9ff5aeb51531668ec9be2bf17c4803fd90a34d4e919cdd47c77fd1c0257bb4a0f5a50c585c04ecafd1a2c1463107a4698ee782ed7308806f4fa5a296fec2d3f44090531ebbf049d1a2f3b340d7ecd318d1b495ec74f3be1e304f588461b9dc30fd2416abc88225029944b46303fcd85f7cc1a34851bb2311a892aa53af8dfc3ed6bc967a6a71a43f191ab239a0bcb03d10a02b1007f5d531acd4deb17a075cb5e79c7b2fec3ef70336dd2ba0bf28dcec2472f63cdfa7a962fc7faff5293aabfd211847fbdaddd3871ed886669a8139ebb6c25603ed4701f95c0c873087a98c6255abd339202f745b931e74522b98b4f935b4176e94099229cda219105d33d484d5a034b0c14c4cc4af9c1c40d66997f004287b9dbed7ae498b65c1453e214d49a727d92f57b7807fc017be1ddb57ccb3da0e7a54d375428b35258fd9dc308d1938c3371d05c4d040d124cc2f4f924a7f9ff0b5a0118915dc670444b4742789;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4034bf9a48b51d6293ead23f7ff0067e8e0e7141c27b34555e15063bea7e5dbda4209125a4b36d542efb03ec39d01899473c11ee6b5d81b7e80acbf2dfa4587b2ef658ba1a60eefba10b70f5fe49d3cc0cab6ed2a5bb8480ef5523302a362cdc9250e87b845ef81ff5b806de2461e80a4d94df23611184109fd23fde519b1b9d958030d50e0c4482681a7bf776b944077d6fb97c55c6ce8e583bd65445ad0e0c4cf2a82bd3e1e2d4e9c67eba5e458728a3f8b488c8017f84c4cb45370cae9c933f9f086338352d94c3c166da1f3045af8d3bdb32ba3313fe5cfd02d8d67be37f7d392e9878992980826ea9bc4b59538ba0c46abf5adb404bf4de8e90093fd3a6fd64ee37bcca5ea2e64938b67875b85a5d72bb0aa24e57563904618ca04e874bda51e37f83481336b43a8ae02cd77a11840af7f6d2c03a7e53dff2cd078593cdb6125c7f7c0731b2cc8c6ae650eff8a59cf6da8ff7ec2e569ea6961a24764685fb12f0e22e35529a6689e0b9199c754b8769e4f717f481562b26f838115fc280c51ab44c1113daf7d13c16eaafe726bcbce37ab5b9b0be8d05a117ff9ee24068cffa33ca93febfa8e959d741bae59b4a2118e30dff5230fe06a69fbecbb22337873f5b117b4737f3029a72455582e3c54c7948bca72654d28381f864d7445dde75a44615e8f9e4f99a941af666a7572e2d29bf39354c210453492baa4aa16c86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he9ddd6ba9fd2df0e08162da7268a33c41470094369d7032330087dae62db6d0bae3e26b1c8d7cd74cd3cec4ada39cbf0e758f4954b920663a47f5542de6545a6194bd1de9d0cb2bcf51b140a3b138b716b189ecaf15f0d9bfeebb66841bb0e7ffc86751ea2bea8634d71e2b13a3c597949c1be63c8d0f6a1f95e0be80ce4495601e706f6d0b9faf237df949d763201e19e05f9c25a48f15cb7e8d9b095d466c4d5d19ac21ddb12207d7932b42be3fca7a683639aeb161e1168eee3c29ed1058388497d45d6b726c4e8d927c64f06161009177210770a0798b4498bf4c973e0ea6c696a3f47163cd8665256a589218f4af3427c227aa8bc96990a73fe655537901eb3090926ee40637d5ca6013df5ccc7730d90280b433a6fefda74c9623f5e5577e5bff36a1c92d2e50710fb26231dba82d8cb7e3defc7e158c8085ad0ddc7e62b0b7ecf8cc2a9ba2afcebe5c06d3620cee0f19ece36d516fce48a4da5397b22fda11ee6cd2155ef6e6d28b71a86cecd52633cdf1ec65bb49f1b5085038a9c248557ee9c3afeb35e51c1adfc6ebd3d985c1b1c0f4f740270274b3950502e44ef5f3d8613c1e62263e51e3fa03cb8cf4fe7d241503d4595bcab4f5bb0c56bfa513e6bdefc78788cf5783f506994273e39fc5718ee2aac1745aa1480d4db5cc81a007ab31c16aa3e9b2299f5b9e4947621dc8ea93d651efe936b3bce03f35e12b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8cd35c3fb84d46f62171de1277ccee876da48cf38450fceec1e72ec88d1d13cc87a56e5d334ab5812df129fe5b937ac42f46b8d32aecf4a51a26a1354309aea6f0cfe611447d704c4da4920ffe16692de209c1ddde822f0b7cb6b673f36e0125dfeba5bad9236f1a8f8ef9f34ff9da866c3dc289748168d528b0408f8916be26e372d760a20e3b3817441d0f805d7f233f53048327e6b230402fda71a54ad940af7da54843e4838dd6f8725bd546e9afeb5a209eaf39240f69c0b4797c0d936844350496a6fa710bd9dfb04ae13cefa9592877e27624a1cadf8ab3ee972ced9f88f8e3e3083701258f8d0138f5b5c93f83527aea26bcef5c7bed02ba2770e291a7cf9165a24076003278069db0c27b399dee8537a903c5b81bcf1e79766a1d72512321fedac0da06227736e4cb49046394a17ef642d694e928540b9a77c252f48982625256d5840e8438aa1cf53fbdb3400aad602a2f9ff52a67e07e6f78c0841056400de0972a8680009e9dae0cf57b43b21f86ca8c363620a48d1eff4a80de97161ad9ac5975e080da9547d64322889fb99bbdd8091532fec4f6f443f4fb330c827e7d8965eef737be452128ec43efb68597e908f49878cc90236f9a3bcc826b991eb78571c3e6226143cd541928fecae865369e4968e5e22695b901b51aea8aeb978628a0ff82bb9aa24aeaa97bae2ba728a339dd28e463e4b51d407f092f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h67e4ffea0fe0203fdc8ca80eed5bb1c23d47944270f7688f6a84d507d90e6c07c068831b0530210d90d7c10ee5e0ee277d371f933e6756fe8af108b636fa974c191fb6c60c0cf7fb6f698f98a57a0b9e45484bea36ab310e08a5b62223ca08fbb060f5fa0359301389c789ccc910d66f4c5496847529f596805b906e3685f127623183ab170eab5eef6c97eb8c2982d8e2d899df41e66760a6b7ff970cbda567bef716326db252710717252f06cd96e1352c67aac76d30a1ab276f3654ad0d71bc72558c29fc2a328814496b5e55e030478d5c8d4ae9f7d83ad8722ba320aa3f2acd5a7b44bdf710fbc9ceb13df5fd0e466598ed7f73453b09f5512badfb18c2d533f128e85429b33345e4537bd290088ef9ec19dd407aab93268d905a9b0a35695a7939e7c77f60f6b3e051873d01bd41284c89559cf77e4296db9072a33b2dd7947a305cd6d817c793bbfc4f3547e53b6e402768f012d558b40a5ba53152ae0d4d2cd9a4098131e6652289568b4316d14eae7f21aa10750616f5efe5cfd10711dcc3311118456387e85ea2461866e91ca049a24fe0c54f9d90fe454220083d6076b91c42eef8dc622849f3c6e81f5b3aa54bc8180a991433fa4f468b78e2e4894b598041f3c060a73bdfef817a5bf06a30351ac975a67d9f8c2e86736b21e1a006752afcfc80badcb477715e8e484ef745bede745f28fd1f42c4eb43303813;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9e7bdc34ec0799f3b9f1cbca66835691880a415fbb5f84d5804fd102746fd6ee3684983ded6b1892a80b7fede0eecbda57534a708fda4a25c82cd566ac1841738297d486e1cfc2ee277d0df114faeb0c23c04cb5d79eec330cbc964da5b40d8ae5e17341dd44119fe9b418ae78f9ba253fd2052273eecc28fd471fa1f72026fb1160965e9048d0663b8f483fe746d84dbbe6b1dc72bcc0726393a731871256acc88b0b5095eb165ca2837690b803ff02dd44ba502c269735bb30b85732cf9152e7ea7143a6a305567327b34a5d3daa4d9b16e2b940dcd2cd906beb84918bb89dff1be3a5a9f6635a93f9e5f73c2d873e345fc93fa695301da17c1652c2716a487adc1fd1a49f03a1a10694b770f1bfbc57a3c0fc15c32dbf9ec34ff53c35179897e882b9a257cb45fdee25b40c440711af0169bc4219f11a535bec6b5ae1a5bcba5e8b7723b28d2b992bf170578737369592ab2fb7dc80c580878e549054aadc70440aa680289b8d9f3c40d3766a1f128df100173b7865fc850030eedf837d16d46e5088a45a83c599e570ea0fa84e2a9394fd50cd5cfc8c8a8e12a95eeb25817e228d592c2efec13e45fc9b3cd2c4c896742b379b54d4cd8283f4607637d3c9be466ff4999bff023ab1d0f8cb057b37e340ca2b1fba051e7daaeb4fb891461c90d8aafd865f20425a29aad7974e62678c74fba9ec381e4a5301b75af8b2e3f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha5d7893637501f4b5f34c307a537d753a8fd96fcf0e66e5dbe71bd53d481e8f2bb0e47c5dffad195796a5d8ba6d403839658e1bc691db3e375139a63ebb27191e257efcb45308fff2640c3c6e48282c786e90dd7cd0537d2e2804a5bc38b0b7bd4eef62fa1525bab480f8045534316eef707c7435ed2689c12a95526484ba2e323697b57af4ad840fb4cb36ccf8d36871e76a989272da92ce95cf1a4364dcff4cc475fe363a7f80525f74b6a23b6bf1fcd46b6b1992558da61ad0c3ec0e7f98fa6fbee2087ec7422fb32616130905851a2cb7f42b9fcf8063b1ea9d26cfd90f9ecca5cf507811c879f8d39ca111cd12cea492d6b547a370f3e8de2ca4dda657faffb4e786982925a29d5c716f8b0e6df30e600e1a2e447e6d266144605cd9985f90546cc84c35bb91d51efbaf9fb3185c36dd8018ef24059ba4ea340b692eb4e6179eb4c024daaca3b7097b629bcc6a310621f7aab467e160fa817e86cebab96aed5a2459d3c76b25a70c4264aefd0ecc4712d04492ce887854f3f2eecc036166b52b892d43f207de1eedb19ddcba00fee724e5fc213a4c038fe13744efc29e0affa401a882cc4aafa0969d1d97ae3b477d15fea4a462449c1104e685934ffed3ce3ba7566ee831fbe70e9b53bf27610c305c0f735c535d2a03813a841c5201cf5925e68e7d626828865efc82593031d9cdd433031b21b9ef2be7b8ea8de32f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb2ea3736efb7d9ebbff68ef2c9d0832c63395c84ea10f35019d1b07e930006ba4727a550f6f3783ca3bd4877acc772b536ed25eb6680337e4da3e2c6c7484c5d6f4a0e6c27e059fe3fdb72de40d59df1f17ce31bacf5b38c890416847ed895ab8518ca41ac3e14758c1f3b00562594a225b7401f6655e83dc0721933726cef772f254c652ce60812917c6e7c0a2b7757341a942fef96c51970a99f8341ee34b8c8966aa4744a1297776ea0efd8eb4f03506d7fa454ce21a42022c69218af2c820147444ed9944926ddb266bdceb64e4318570c22a0bc1733a74da1900a70b07404cf076cdbd6e5d29685e74a7953c33204a216e10a6c4e0020f75fe360808689d5d611790645c1756870bc2df19f69e742203c931ee0be06cb81da3b221dc5a70f76236a56e63e0a2c0806f89186b8781d3c82ea58c3073d39bb2bbbae9f0194871b3e3eda97606698ac74933f9e96df1d4304270d26c188305976fa76535a3877d59284b487e964cd337064eec372702f5ad7308b63a03139fbeb0a111e5ea7672763d970f0952d36cf5fffbe1fe785e9d8385d5ee229370523f60fac5afb7289c0fd66b7b4293a94de8b9db07c637bdd8142e6d225b9149ba648484d4a585597fc99ee5b85fcee02c00700ce39cbae1f1ff78e0d89d08b23864c0c299c705b6b5069984a6aec0c0a262e21a83b4501908577312594c6908ab9de8676f37262;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heebea45408c830acd2d99ed86fbc2a49dc14e3297cf8d6284429aee7894409e59933519da817d595727f812888c629b725670aadcf642f7b83e19c0af0a63d483aca47d8a09344174f02a02b25caba9f375953d77cf9aaaa7e86989916cf0c24d712f7b5c74d72d8a4354ae3c513f332f5d3ca32bdc092053fc95c5faf53c50d90a9721568d5f75c7093f383f4ef59ceaa48c258e1d6f0d67dcd54f945c770fb77accde29b0e03d634c24bf180aaea1b21972ebf1692361e0eb07409624d234655ce966bb06b3b5b548b9a583ecedb8193e49d3b58ac48b669494576cfd4adea08d52b2c1976a446067a7749ce8e17a583c40df19fa68c1d9fc972df4f4ea134c5a9c93d7b6927c85cb2f8023264ed5973f34f9dfc11c965459d7b4ddde48e08df5c1f84fb59efaccd11bba9054aaf94e651c542b0633fc37f373c082d3cf22d253dc50fef7006f494aa5d8a15bcf5df75171885fc4ea1127f1b018a9772a8844fddbe5b0fe26c4482f8cdec5de13edb9e3080b66315e4d96e5ba0fcd5e2caab847bc8afcb5503107b9ad9b5408eb70fdbeb7fa4d85605f30b68e32727ecdbf92d3eea854c9504ed65e7c37301798c4e47d7a61c9e2d8f767b9bc9ef5f9cfd244a654b191df1bcb56376609ca2149973b3142786076d725ee9ef4230146728ce7d7d39d035667ed4f98d2488bc88150a108e582ee58b4b88b071d3cb2ec5969c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4504e94fe9b43f7d94f0f3c3f3306cf882f030e34cce5dc3244ddc10ef948cbcc78debc89d26f081031b17397f39d9ddeb58c6bde6968aca8498a81d933eb9368a5c85f184637239eeaff317beffcb6870ebfdc9796d93538d14451d4812bb94e8960a1183dfec167de9125f2d6f917ceff670172cdec51e5d278bd532f00d63a933c3a1015be91facd217ff61ba59c212ca88f018cfc5d5bba313587d7694ea054889fc01e7ef4875444ddd2fd58eb150d35f229356618cb8ebfde582aa0d1c3f1b40b035ea0aa1c7be3acfdce11b5df8a071de94731d8f461e43115d6782df2e958e0c017490ed1e106af8056ad8be09e73a7be28e7727ae8096aef517d30fd207ea50bca1658bf9534a1c105d7354554407d4ff31e7f6c151c78431b7f8550c8152a6f7dab79e6d456649c3b75caba603eb772f2af6c325709ce0a6e1ea9b7342c3bea93559fe6897ea59c5e737136734b980946f671cc4ab7fcee89e51487680aeccd9b935c370d4e23e2acfdf9d07b30316060bb43b7062cc686a9f2839c6db602da26e5083962f48e697a21f4f64873f4e747888277ae851eae1c74eeb8d9b875cd194664ef19e3e4206caef6814931c1bc368547585545de6e540eb120ca548056814708f2ceb78f1f0de2ebf4961f8194ad286d24b69905473ae5f8db7cc950ac7771f39c2210da91841f880e0872947a18fb456f911a973fa90f218;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h44b9e84843d3af355588ff8224c34aec107186160c26cfea78d77e2f81b8d80b61aedc50e887f9a8bc2ca33b009df909d58cb5141935d3f6522b2e3c807feb7d75e01234aa4431355d92df149955bd53bb5c3f48d933c115317b39079e534cc2a7efe8b986b5dd83a2598cd26c525a18e1af94a32276454c3986d3b36d51315179f2635775270ff2790b464bcb16d6b6c3b14f59e172ef431bfb482bc6388ae76686fe54e9dc9a206326b86e5b6bf7c5915927dc302999f69ae922a841e84fdf1a5ccb3938f55d1577c94780889a49622a44a3b9e00cebf03f53ed082eb53cb6aa78e1eff24695249339a88b6758774fd00a70d43fa79bf2bb51e68d93a222716b041690c142246439caa883c6c6e574e49b74ecc94c24ee8ae4e8c083585ceb82c3f87f1c260e29fe01debf7f59847c17d21ce571d976f05f643d4d73de57ebecd02fdc163a5daaf834d2b237e271e5425b212541243f4a29b7b67a79aeca875b48f217f8df8bf2938991c7f9a23ac42d5246e7760d3b617292057396c9f713606cc48432bc3849f7e8de09af7ff7ef08e593dd3df64aac0a4672f25b9bdf8613b2478e6d930747a3b73459edb4e8766cb36bf836f0a1199139b43dd34f924d7ee3ded8aac0c60db1730f0efe84c44c758f6d9b62361d7e2e80145033c6521bc877ff82935e1f15f2c23c5dfa95d2862f8789eddb465902a4e95c7756b40633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h662b0e54a8f296b7c81b31df9f5f8d82617c6662b38a41473d407f4463f058c88645bbe8d692194f7957da1332f20a21b9ecd02f3a80e29d50679ed1f47a34bc9fdc4936ef515348d3b98ee808307cd5d6c6b71508a43b34fe704a520784db76c50267327209fca4f520e1b47f65db7bc64cd151bdc85198465451a8a500625d213ef4af8f3dc1cc727f13a5259bf88a48cb4f23286a696b10096c7b68b7926bb80419564d7ea5484a10557cddb6afc51674d6af521a5a5d3e61f922dc559149bc588f2ffc7c77f331aff97aa0232f5d083b3c4f4c1de84320436e1d7f384f2e35d47a8ca117ec0c6c356031b666596e68c096e5e3b2d26d1fe6cd6c2674c262fdf62414826ac043b8a56ae58784b6fe34e7a1fca59d305a3957600fcef18a4f421c7b2b8201e332815dd5fbe661abe6bbf7e3657c643dbb04510b77f27cbbae9f4263644c9aee08729a0889ed5ed199b21d894bde9b5d3c10296fcb7a060fc0fa05f6fc16d8c362119736a7564616318178ac65932eccd2cddecd583003d4b18fb2b9e08e70c001a0fdab5ac53f683e1b749d1821b8f65bc1331ae4f1e8ca2fbf7ca908fb5dc63bf928f282211f075c3a3153efe67d41c6018a307e2bcdd43c538fa097a30ae428ad70631cd98eb32cdf57f1bfc71c923971ae0d455a0d998e0ea3ca1efdeb4cbc6a85ccfb80c3902dce941e04ee7a352d2a8f5f961ee80f71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h89c937b3e9a182465d266252f964f2f54774979dbe3ee005c21ca395a247ec1101f7e5f1be1a30b4fd2ee4d28098b8b8858c694cb525b3bac818fd49ef0001fa86c967f3c004647d4b2737f9677ec933c8e1684801fdf1eb5945990ea3eb390d7373959e97afdcd135e7c598616a3cd85954772bbc996ba01c1917dd416f0c54a7b4b3793c66152059fd10d3f16622635f47b7512a77d7f77602a8a315fd6923954e721aef08536803ad07bad6ab37a2a51be5437e94953e0213e1831b5fa07fc4937ba4b955b51c4976dae380fb40c22772ccaffbb6e676bfe44fc2cfb2a7e047ccb331ef49d253511e56c6c8b7207cb1d3002b2d10786eceddf00f4e0908b13192a5a8ce0b213f7798678b515d6a2438d941b9c19e767a969779269e9ff9f998dd0a4138078d4a3521bb0e922cdf2335a325d57f1cf2075892875b9e438f813a5b5f48ac1939c59b0616d8b413702a90ac24e76af4e622b21e61c2903652d4b5f585df8ea92541a1e06ed07120487552510c0f4030a78c2906b719b215fd6f142a637122c2cbd055292a83dd21002d30ab0d1a6814f2c9c195f9fa39d1ad6fe6940aad50cb185489e90832d7df8fbe5b9bf2ce6ab4abbddd1de26b3d08c46e8b4d50e963790f52ae035c39cb7f330bb04f4d635e53413d812d8f42bde16c1ecf5fd07b7b22f69edd1989daedd7e3c34ef23d81d009ff2143434b226ea41a1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hed00dc8d15426a16e4d86714d663fce4a0ef176b9687eb432be342ee04291d0c2d27d0fe9723ceb497649fc802c2c258a3833f70eae4529a1887cc332f26d03a892b8b221815c7d76b1a189f2926970664950f2ad442ebbc8831696ea8f484e376a300c2c652cc3856df066552571187f005edb283cddbe0cb749ae4f8a7e75a949a4f925d7c0606520e2d6a4c519817d7b0701437ceba122928950460f443942642ec25c962c4fc02cc7f5e3270744cee16f0948ff099fccbb42e5506a9915b1a21548f696291c4febec94a3b9c165eb3a8feb972fae916cb1190acdd9a30b92282e6235ecb57d1e9eaa879b7ea554b5fa79bdb5c285f2cdd60c4dbb3f49e8c63b6f3a8662b505b2a2d1b6cabe42104f15d36406ea3088ab67a8aaa718aa951f0bc12e18dec1eb88c81e1f395a36ed3086f9542b70b703bfd1f138ffbf6fa9cf9fcc864b20e19297a1285501bdf7e744ba923e0b1ad788a2432778d96692abb20b1b308c15b800ba17281e07bb1a7ed771e78ae5d892beb3cc2d8c5dab970f319de1c2277322bea5c587cb29bd894f7d4380bedc84fd518dba3b92c7df281c9a0f70eb107f1baac6f5d3d86b20161db979a993605d54761a81dad8006bf8d8d410d67e1fb935c954de49103089c31779281ef4b45041306d0001c05e0acc85a2c4c02317d32ec545c4b6b0c4a78b879c74caa62a1d949943d2a09660daf4dfb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6df318ed38941ce7b588f52b111a806f26ff7856be3ec8366f9406d353bbb9a8742f3dd464b2c8c79f2d1ec822ff26640cb25890a57912efa10792a0331e2535648b1b47ab89d9691c93fd70ff5d5d979ba5b7685a02d5207fc78a7bf51536c73852d8f23bc76e6248b865f5387defb71027ba89e502c769115a1571912b2018b0e05bc188c1366a6484d8cadba0b334ad46de46ad93495e0b4aa0bca796689b7fa9fbd43e7476301c400a9662e0b019e04579e20e6275d2d985434e67f5d00f99e7c70a208b97d403b26866764310135f8e6834861fc4c4d4f81b8db0c3a1c3ba87b943b175d94111a071788084d33ecdbcd9add37026217b137594227eff6963466279da5b48a9abad9d1c4d1f303cdd8bddc21c5dbc0570fa38157bb767a1db2de7fcaec84017ca301b4fc41c62cb6b8635b8382ebe31bda6cef553746577bfa72d526ecf2099e8c85fd46c2ef47d6a7e81761997f51f42e9b6f4b77624c4bb7611dd77bd9349410e1306fc7e4f91fdbf8e9b9e12bd7d1b3d2f8279439f032f1561754f91f4f95b5e69f61c116751e8ca4bd4ae72eb421cfe459fac4e29cb3dd016adcc04f71217af2a6bd6b70a6e7302fc7105b1356df6929a0192a097fb5735904cef1fdba974c12e400457e6550c564ccd1fd4d63f357218385457f49f99ec0fc72e9b80a9843c3dfcd81881a00dbb747c7eee55ac51c999c2731c966;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h246cf271987480ba27dfc03a58c1d8b7698607381f4a6546b310955d8b41a195d504645773e5eebc85501adbf03edf45d54f6198e0b6bc7994e3d4c38d86271bd1792aeb42883e5aaef0f42ef676f7d70bd45bbf058930a8b3a079aa7da0cac683bacbab92db10519ae4cce2cbfe3dc55120e62458f80a7b17f290ec45ebfabf9c4c74d59b1b6405ebd0d49c33009c8070ddca6143a9f0212ce79acd505a821c986b12ce074b30276ad5a00ae98e7616c20ee85f031afaaa3f64daff773d407a4a27c2cfbd33fe38ff9ba9234fa3844ca68728c5a77b1048a944109915ec309de94d8f47af58f014eaf3ef2787b30bfc805aa388533a9136ded238d372444525ae37b47d5d01170afb6beed715b89cdb2aa5f357262c88cacf611b93ae7851e29e0b3b9945d7320e63a9a500b2ae255fbd46927366bb83c5b43efb650b2a47f0d59a814ef262f8e25c0b6cf0f32c777fd505bb1f6322b21ca6f285de919ee07c95fb30000832fa5b56f8bdad1b0211b28242b612d787876d0a0aa12b89ef39c1e30238f50878fc979033b1bef89a895d82289b8359058fdb4cbf7fe17b9325a94eef539fe750b6e6edc9b4e1d11beb7e5233ef66b3deeb47311a8622e8930065034887c8921fef096a975bc6869eac553202e8299126b77c709af5f88d0db1743a345a950e01174c087ee1b55228b9cf43caa809eb6a92244ff8a009a6c36324;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb77d6a0064c1c4233d40c71a3e4a140b319d7b710aea3fefdd352f5867591e108a8be099889e9563037f1e9f56cde741eeff20ea8eff55efc46d8b8d72ed6cba0ee80e6a413e9c25528e387b0a329baf36eb672cbeae135f2c6f50ea082d1619a4be41818306179bc3cf0e6153bfbb54899a9c986268904e5e15d856e0b08ec366053d308230b778d62a195e933130b18cc92e422dcbbcce8e06fc8067cc321b2eb0a434a542971b652bfe25aea70edf12fee5f7b8e89273e7949c6f462ebea667db106b9a536f3179c8cd8b94fb7a479657f12cf65b0c8b351c1a535d99653614e94aa4cd8fee5010422b938421a4744a4de4f89ca7d8d7348cb68b948d62dff773d57b2eda06c7b42b2efe603b3ef296ec65ba3d30e3580e1b71c7ad49724447ff28e156e230bcb1549d121560f4145bcd97ecc67803f4469039c9cc4c68cd3685f99d4faccb6de1e745a51edbd09aa5c664cd07165a056cc772cfdc3765890b60821c2caa7aa12f20924bf1abeeb2f34d7e852fdc2b5d9e98bee24b047f9615289e5d074e06744a0d439e7b366b1d426cef9f04dd5136aead176f370da05fa81ee1d433efeecba83d2b102af2ec499c63785545903207d78a293e6bd1674ab55520f3564ba69c8276f59c7b72b7feb7e14ec039dc5043b4673a34b3955b19059d0c31d71d12f6cf773e572fed0705d74de92acb0d72e0e0606752a1f96649;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1280520af569b606c85ec3fa772fde7705af577592bff2564e153ed5c11ca42cea0899a72a3a9c0c1b8aa02100f4f875143eb2dfe65feaedc635c2735524d02978479f644fa31d32f919ea27f48bf6f29e282d3b3f9e448612042b717c675e0b7a493489e86b8f5ab5b43a3c0e8c9c713646f350583102f1d52adef661dd9eeaf16736ff7d368ff40723f5ce6c29cfcb7f68498e70ca41dbd1e1eec00cdd1301f16b2e3a7a301a647aba826ad172f388256ba5767959580be08a3f24704cc039061bd2178a88ee70a920441b1ecb12f807929d3b751dd87c3c4ac2e6d710a26d76e9b8a033299699779d996853d83063da98e18d16b2f528d0c83524207c098b2d462f24d959051f76ad8c23e807b157354dcfc4b3b76921f594f6e570dadd657b854d265caa78c0d4a9f1ff40f3da34a5b21a34ac44a8181131fb31298242d75d3eaffab9d088a91a018ef4a357d16b0d04d69f238a5752949c14234d7983abc52f3bba962ea8aed1dd6be5d7c3777f883d6c247074f06a5d6968094ca3c2f95115e1a6abdbc6af6f333d952301d6cb0f1124e13d3a7d751ce22289836b9bdd81493bc332b40dc63a3adf7f6ea814b8c5874143748ff1d048ce16d2a28271e630d324d98ae9e58882bcf4a69974e34e39494775ac3cc44a79713764a2ab2f4721aa79a6c724e09a58e3d3b2cc8d36e483c5249ff77cdc6c112dadb751d49de8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcbf990e6d57c71f0c2f07eafbf391482b55039d4076602b4be55d9fd8785a03285b1c929116bd4f9f12885940a8668cf7cbb3da50f9efa2d9b3fd70fa9fcb50e838a226fa754d7a84ceab225750db4ccbfff695a416ac470524b79a821dcafef24ddb0b547243ee044a8013b13fafec7a6ae3c99d9d5881130893747c51c82ef491017681145dcdf6574f412cdaa6f3049474ba773643ea6718a6689a972bcafc036d8bedf789cadfd2a5e7924234d76437a958b82ae730d79a38fc56134eb5c35911b759c73af964bc3b954c1b184f441e47d876f377affe6be4309062b5c632fb7b3bf8caddf6ac8ed3f973fa3be985aad11ef6d98940d601f2bbd88be394e88e3cadb27140a72426d6eb703bd13dbd3a42e290fbdbc20ee110d800775c7b11c67f420f25bdf736a3c07bc28ca38ccd67b303006e1d3fdf328649dadb5d5d1e81e595f5d4c548c0dd6e5947dde4e3fb6ed635b607a23a992fb5143c4207431960c2270ed08de8b292e5f5295ea0894f4190cb2b896d1153ac14f815ad9585308dc741ad90193414c7046cf4369fcf35fbcd99d461085f36794f1566c2a60b8a4d3fa0719fd436dea833e24481ecad869713781481b4990b4ec2e71d52395a78e570e34de5aed802973933aac63a3101f658b2615eadf2268f03c80281baa4e721d8ccf7b26d31d7e0aa4fc2b1c96d5a8d717f9b4e08e6b8228c3ab86f28d9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8a4e8baf5cdc06f1d117efdb2c90e86c525794fc8b4f84a53077a26f19d2d8ff73d2070e8c40dd004e94e26ea75cf8f3eb6c9dcb6ab75473e4eed0efbdddc4d502a0f1ff716d208510ed31bfda488448f2670dc4fda822d34a820611fa22648a76d5c3fa90b42ab747527c734483e318d436135ba9c4e762881205c0f4ab21ba4e791490c1b0125b782ddfe6141c71f3f8ae6c706bf7d625c21b0caf3c9e548f0958d5cc22eb208c282bbc351ff6788636aa9f98b84fee93f619c67379804304aa0d7e5f75f2870afcb4f98288caf3a94178dcaadc374970a10bf6408cc2deae5a44c23bfaacd49a18cc1769a4714a9a59b4bc1c593d7df8d9b6c1bc95afcf7a7183bb8cf340c77503b483a13ceec0a3e1e058048ad63ecb88eb19418c3499575caebfb1b110421bc5b2fbf47107c2009993bb71272b9bf39dbb973ba773c62471f4577014956cc2250a6bc63ea3ee5d4d89e21217b51a81811d52d4360b5c34f97cbf936c9653eb4ecf9301954024bb3750877ff49e1af4de0dd4c1c65496030555f5c8a6aeb283b0e872a2f5b606693502307141b0dabacffa71c1fd155f1b08e3edae7ec74694bc92d7fc66105ff2e1aeb3aca70671e5ef138909c3b27c667953438b4d598079ec82e5bd342fdd59571f30505c3ede5a09f2e574bdd83fa0a392bf086ec4816dc6e433ccc9dfc35760d46cd43c18273d395b893b0549da43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb184c60bb4da7f99360e58ee9847ec10ae347e6652266d3fa4c9addad347772996ed3e4ab00540bd60dd5025e52b557c5cb9bb2945fad833ea96b692f691f4d0964f775b8be65a95ee1f80a0b2a5c10e853435cf1835f12535048281207483dd597cf5768a419a2187f80ca74dcb5ac1d887cae496c0cbd0a55c72a0915a705ca3edaea86b2f750b4c05f56fa6534bf7acb3263de2d32ab0a8cf7a1971555282260d38049920d97758fb36ad8861587255e0aff0de74867782fa1ec9c9801f5f197eff90e87a085fcb4dbcdf3b69dd376fdf5b55e4947063095d71ca8238ee6bfb12f67cb2e9f9153174a501e788f40d70561697c402b6e44c486a810366af817522a8c74ee69f6445f6e688eb1d060e51bea9910b978283225cf54b333902fcf3bc227348c68a6e8a8f3b1a2fc23da9c1be79c7e6e7bd216edfe49c1cedc5b7aa5f09f2d0d3f5f7d10d32d8544030c3ca04fa15a68971bf0d0ec036cc8ab47cc67ea265ef4b8652482fd71f6bba130a3676ada5793e573a3ff55d70a30e015ea81021399f67d2e56a28d499f37f4e208be0e4f9d2b57d4780f25f55bf917185b1aaa5f9e519b91341636ca64809772c4e863ae47da9b823591562b71fb04b480fe85980d9ed649b17a12c38cb68e94485cac499579ae0996343124d9ca942ef557301a269d2b490f16db044f5e98f892e520c93ea85318221baaeb4e47cbfd2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hff6f5d2ea1e09929cc0a3d48481cdf81bdaa99b4521894771d70e644c84b2774c7f08906cafc8c2ecacd62da44ec882ccab88678ae9ebf2758fc5faffc90b8b2fad688a5c22fd1baadc6ebf350392de83fd15afa5a21c67557a48a3ad5ee038cb39e635c7b420af836396dfc59df0f3800a2f84d98972bc302255ad6594be322852da4a8fd092174de4ff4e5fce33e976a95c9836c67ece4c2ef949d4af2f529afea4fd9933d7c83d715642143f3065e081c18663cfdc81fe2b1cc428d69a0e5e8d38e1b6a0b8fc72ee9af96d2b575fad42f9a2a2f43c0f43a3e3361e40bc4072fc0fe7f74edabc1a3925b2ac66e57821c871c3018e5b02d70303a29ea837f2874eac63cf6ab594ee3eae65aa11af7fcb1302171d1969720b1edbd38517726674928332f3874eda248da3f6d340a18925ccaebfcc151074008b1f4d56c1519f84f5a080e3dfc297f50b8d75bfeaf4328c0d79deca9813f7e2829553b958f7861276f110c665a9e3bab297a47377b35904180c69b14dbc0d1160fa30bc66dfd82ed36e648f1815022e61fd8be6408f19fa4317fa5984cc9287004fe5c252cfdd92a386747714ccfae7886d9a71c7b932790be2e18b1124938881027e0196e8883940b506ac22901de51b8be34285e888b6109eccb93aa3c1bc3d6fdbc507b09f7fc0903b94e7d74ad05d3d14afa26e9fa34cf062b7dce9d4adb275005b324f91d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdfd4197c4c6da4b5c067309e355c256ad1c227786980a1b40b5ccc6b833416e8ee591b483cf478da39491d98afbeed1d0d0eb96dc6e6cc6b96719d61bcef7e8e8158fa06974b78e0e868040e95b86cb804446becb489be1897ef5b11799ed3fcd79edce279415b5098f842dd9c59f59d6554f3936b34b58b2716e4362c4e6973652707c27c0639e12c621293955590a202d9c02be7cce7afde4a6d59d7ae496fccfa295c4ef1351d2aa526be0310e3c4ba2fbb54fa0c7f75d364e232fa92a8bc660718d334ca9a6c32c7c7f0e4fb4aa975e3e7d593a5b25fa4cfa791cf60dcf4eb214de21de3f4139ce015536e484c06a435dea47563bca52296d85ab4a3cf73797691582b50c764d38828f54f01f79f1212132efe67de9cd943f0b18a932bec678c7b2818d4ec1c004f95fb3b95bfcbe98cbb50320b62f8a3a54720b241f4a5d966800faa6f516695119e8c9b1c184f9a426265f58c2c7d4dc5976963bc46e26c97c93e387e951bbe1207c9ccc43e124f8afed13aeb6b84363907205f26f3f6639e007a9d7aadb71de434b8473db248e9119acc4cbe794c35179cc1ff6b9104f913f0d9d8a77fcf4957f07c7b8eb825da38968d255d299a19ad0022280017399283c2cd226184ab688b2860dd53192f7feeb8b7d9e4226679ddb09396a696cd216abb99baaf57ef09432164d29c79aa9f6c7de84f2e8ce007288ebc3ad9f0a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc345dd6e210c79a1c9b0aabbf19ba649f567c93107be05504f5d68bd0f35ce2d7a784ebab3e3dc4c730119e2385cff973e99096ee18e14426d3a27b5c48c1ce6e62788f76d87c5de32b52b5ce2166770d287f8c6410f10de8ba08bf58198e9a8af614d8cd60bc8378ddb04b4ef02cff5d8a7fbc891627a4f65f381edf0a449a8e3031f1aaaf9d63b7cca8dada98a8663cf471d84b9d613cb99649a3d0e756ad2bfdf18d1a226de30a998d2da6f0b54d26fed2849c3f45bf2fc41d0f193e629f45e03e60b43c306ca80422cb4b2f4b933acdc20e261611543c648663812caba65430c3cb17bf76640d86a44825b6d8feaad358ad186652fa9b37b546fcb3d442bc43a13558d6399029b41a6574308ae86ad4ae3b0c52432d47a3691de6bd16e3d3e33277282250cbc01b55cbd4e352ac0d0e812bb18ca4f1ba8bc5279dc25d1a6387d046fd97cea524a2e88d4da23c7661f3b7e63ceb9aa81d0eef7146a4a338345037032eca30a1e12c738fb13d006f610ed1da72a769ab6cab96c4e638e7eb081745ac901a6a7ff4b306c3db0283063792b1873736c46047d17baa81ceda3b934322e964975ec7d7c782c9c9c09693ed319996427275d482f194a58355564dcfecaed495e6721f670805515d2691e15de8c00b0d142a74da38c792c3b9aaf15cb4ae043ba9ea2ad1fe4a9ce125527b22a5bfe8f557c9471d29f637559baef04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd4510b688252210386c5ecbfcfed71abf84197abb2c92d1aa53d00c541dff64e67b7c9978d9c75b9486f4bc9a088bba333dbf0cf1ce455436805fbcfae45a8922b2a0de4a017c9019fe40816be4884b932dbadd84cbd12b666e09f9d4c66f88dca980c0554948b27fc38c9d22ce68d886c5a43afc4d54422fbccbfc8c520a94c7d75b5ee5e1c640dfc0481ba381af4cdcfbd6e9a83c7e96dedd4e9ddbc5af358735de1b4171efec0b7254c6b848f96dd90b688761e737e5752a686932ef3b9802c82f532029ca61057a472c1bfbd3616cb34eed134a7d006d18e75197e83bdeb1343c05f0675e4dcfccf13c52904af6698310cd927c261843e8a58a9828b60ba5676626f12fdcdf5455c710bc46a1f2972a7bb158f4d622accb0fa6c20dda1c56456ec95b6019523707d72b8171514b58812152e50286c5bb5e7f83ecae6e577d781c228ed55775b463a483065f894e9000191017432f60895ce4fe707c27d62cfaed55e8807f59a213978f9f15d7dac332c829a0dd9bc2ec38edca9ce999d6202ee4b11b3de9b0c2d2de713d561d55ea99e88da5f9e0ed6000fdd0addb3590a4cc594ee2a148ad5e260290570e7ba72087299f665e5a2eb983cfcdf281bfeb115d7e7d68e8049b25970421ba538af570dbc95f5001485d2691473cb1650dd1548016f098cf12d77c0022c213ab42c16ead3c06845e57aad68b5608e30c478bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb9ac7599cc9276aac78ec73163c767edf61182513dcc7e2ab61495ca9e992e576288778bc726406d30ddb812e387b84872cec6d162f930614284cae90c3360cd8735324c905f769ecdd982b912704e394488772ae6fca04475647d82d99657d5051b094567ea74daf3d1044501835c9ecc7ab6c5230d1d00ec9a23a247c8b711e6095ae2f3920c83c975eddd9190beb3485f401141fe6bf3891adbaab08108d3a709de3310a87bd922beddabf54cda2c9e2b45b2c6b99192fa8f7621aa2b2df26544baa3db700d2f6bdd12fc8145f8ef20317fbd758af2b06b08ecef400e40300321da08e1fbab0a9cd33639eace5847dc33b27d8ea37d30f7f21e7763e3f3bfa035f60f9666eed3cdaf8205d86da4d7b9454572667a56712388d74088c010abec55ee2c22cd4cb91de93aa4f664e1985bb87bf60c6e682236d00e48c21bb25bc3fcda106211d5dd9390852905957a5e444083a32b9a3a52c2e718eca45320b1842b910007b38a04c15ae826cda9e035094ea6be77a2952075be58317d747a110784af4f97cde516a0c33cb50a6378aec5c92317891e86b2cb6607d14940f9f4eff4f9d62f7eedd5c7380368eb3ed1c9ca31f18d6dd5b0004639ee8dbd88704866bfee83a3563d76e06f0f3d6d92a4accf591d4ef15a0f829d9976998b6f6fe9b23547bd0d28c7267c022e97135f34847633c243b51a0ed2f360046d5b9fc31c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5f463cb2905991a49936d24e4c527bb98b24f6cdf3adf2192863b11db20a41b8a75340e4d69a89094c58899c9554dcecb79c6fe3296fa4c683f7398b9e4519270014a291ce97db5fc9e369a68018d9895b12d24d110ae3ebd4f54909414f6668e3475d8c6879c65a57cd56f170c5174f9b5681776d8329807763954d45cd9875f38ec411e0497fac3816cd8bd16342c3fbf6fe6b746004414e4d8c82cdcc0110e2a7747defdc334e739da7580cfb7a1a3a660e5f8b8b34683f2199094d0523a686843f5d7e0f0ca0a23e120e5db56569057fffb60bc878aed38085b859bcd6f5e44feb146f48bf7c82089674908306b7f70a75709cb8b95778979390eab2de468111e00545b49e565fc872166741cc9708b26d4c553188e8a09520426c4a2d17d8488dbc413258aca2e56b51b4aeb2e2b6516ec7db2d9a67663b58a7c79b4e8119b4812f96ad0c4945b7bb006a9f9e4cab39825ee6a46877481443c58d7a3840ece6f5b3f2bd02ff6b6a09e10aa3b9bfeb647cd4a9de7c91773d7c72afa9d405384275ae30f7fd766d47cc7247e3c8b0453a625a2c20d65b23143ad580d6350b8a9b37e124c958d1b816d50614997f031e716c88553ace4f92deebfdbb1dd58d32c765d92c95e983b9dbb9b8cc3e88587b5d59041827e60b5f35b7184d91a8e55b4a5da03de6efcd66527d6281b9a3ce9a54e5464273cb70ce10aa07405e86ce;
        #1
        $finish();
    end
endmodule
