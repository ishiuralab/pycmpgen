module testbench();
    reg [14:0] src0;
    reg [14:0] src1;
    reg [14:0] src2;
    reg [14:0] src3;
    reg [14:0] src4;
    reg [14:0] src5;
    reg [14:0] src6;
    reg [14:0] src7;
    reg [14:0] src8;
    reg [14:0] src9;
    reg [14:0] src10;
    reg [14:0] src11;
    reg [14:0] src12;
    reg [14:0] src13;
    reg [14:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h926c56f06b00ac8e881ebb155587086c9dcc799a857993057435c514;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a100eb09f9c13086ba3e7963ad4365c0ba391821a971070d5b01ccc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cdd42a10bc20857e976250bb93a3b99e7c3c2b53611e1b5960667e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2d507bbfab93e7a05d6a8eef4aed3eaa6c5ece621b5b4148fc2574a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11429a77828bac5ecd6fe5e796eddbc719ebabc0c3d07899ccf4e6438;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he48574515b17953851743ae99a55a4427b770c1e87868c9ffa47a60d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h902e54eb7024ec1367d97008b1772656141e58626a7ce4e9c636864c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h219e6b702dc2d0ee7d0f614bed73ed35d93c7dc76904c77a9b9a5974;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f0b391e4074a311a87d390e308ac245f17d5cd4652194495d4d4abf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h146fc1aa5119a23eb40f7d236ec5f6dad7aad5d2727190acef1a53f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7357f0f177de8c7e141c05409a64a8f41dbfc3b3881f1fc6b779a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0d56cd493b6048f9ff17d18ebe8d0cd0e9e2dd8a1e9507e459b6a13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4b482fcc1fc9e54677aeaf85e64179d9512852316d19fc05c3689d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb535acccbcafbe4451ae57a1399456cfa82ef564aa03adce17a684c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c42c5a12015bda97500e83694fe34501858c01fe5603a7b4cd940ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3455b52ea33bd6dec1dc36cb138f1660b346bd25b82ef3a47585da01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148604881229a775d84d289e8aa12872f90a382d34e8f1c8f42037516;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37fb907292b182c1f3e68f986cb629cd3f2fc2e2c6f26ecf56b54349;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h46637cbdf68311bb58d37833645bd9a15b892f29414c1db62bb86c38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2c48c2cea2d0a94d1d839bea9ebef0bc4ded967ea4ca41fba9d960a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15476b6db8e90dc4899d0360048c9de321d909ffdc2634503d9eadedf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6e2224fcb72a142871107010859ac9c1a2b766e837c6ed8db3436a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190dfc664c5711779d1ee48da74331774f4fc269aa99ee82199276977;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec82158b6793bb437af823cbbc828e315721af71bd63c082bfc1cc1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h750983deb7d940ff8639249cef23facfdcaffe121a896f9b3e296ad1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf1d6f383497a5fb9b9684d293ebf1250aacae00cad84d93a14b5116;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae6bf1faeb89b1f0eb27f8f22f653ed3a8547de07f27f33b51c5c88e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h54c7b4e06a2c8effd3bdcb88331bf3fdd4be63859fa363129b64d72a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d1bd60a012d551a718ec5f58804c5223e4b2465790718b17bdc3e45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f51a2a6973ddbeaf9d262a69988956ca1abf563cb28ff5800652610a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19494f53f537e4df200f9e385a90d063d9e613bcaeb5e95317dd3d233;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a561b0345f302f3c071b3d32e865fd0edcf5a91762b25d6fa0f00f24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc39132652255ec4b6b1d951ffb605e6c2cf4ae61ac4bd8a2a3b5ed8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db1a4027f5a55adbb564ff28d9784c43960c2ac1b8dada1beea909d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf33e694f0cf807bc8c40688e8ea15060f13e53970b70c860dd2de9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8dd875208a839385bb8dabe0e6e8fc0f61d1d836206433a06bf5d65b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b1fee46e831bf660130c8b7bc69f76edc4dc806fe02138db4895163;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13b269d2110ff26869d2cbff57e9582d58028e0802ce2c7818ba0ba58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6128179c35aaafa3d9c286887a85efa4b8ebb29a6c6c734841971373;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17b41e287a1284516250c59de88544797cf1c680ba2df4d5c8c44158a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h97e52b5f9c2c1a39c8266cbc77fe9b80a0aa39cee1d9397b335d6ac1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110fe6a6d5ef3bdd1e250de7ff50cfadf855f9f475a8a7286d6da6a29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190f2b2173fb28d226015398c01598a5349d70c33de3365db09551c39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b146f225fe3a3953fcbae812fefe1752187baef039b5c0dac9103a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a038aeb09ce0817f6deea608225c7befec8d494c8c7c44914e5bd85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171d0fc42e1c2a04c442cc41a0f100c0a1c77594bd1afcfdc1b347838;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19b540cec19d3c361a4b2411fde61c744626f3e79bcc347381d0e8796;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1992832bb35499e36fd441ab14ddd2462658d771666157dd38e4dc557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c60668ada74f4668745c29dcda29031c7040620a4b62854922bb8e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123dd3c6210f911454402563490e1f4a8c0bbe10b5c16ca7fa88c754a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2e671a4bf85b1df646301faecd0531a3bc8360dc264230b0d6fb023;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a34f85319183efe7d34751c5a1b9ebbb08a148d3f768f4080276f7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c766a687570808a7e1873c31da8ddb0ef2274594063305b8385e5992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hab5bbdbfcf38a2aa2be06fcb0ffde1c5a7ca987f9230b6651f487c78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he33a2a99e5397dcb61f17d81e56c4d0169b96d70b18cbe60d00008b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe6124362f5ab3584a8e078aa5417e7e221131fb62ccbb623ae17e28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103ff89741a3ba85576c340b55f33ae7eca21b5e2d5eda0a1cd22303f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19767a04f904208694954c8904233d3d3247c43f93fca022e2d39c324;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12774b21b777776670fcca19ae4af0a94286b91f37d8d557213717ac6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14368f0292e6f458d855643f5a2370e3a639f79a7be79f4b86c9c8fcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4561910a7dbea5813de6c721b627f7f84316f9a986987178f4c322e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb317d6f4b72721e76b573ec77db6799119d23709437cb9892f2070c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd440265d78621169e3eb0e0b75ab3a4e385b5b0477e58b6ac0db208;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d83689820d092a1d83e9dbb7056c8fbe7c7570377364543be8b7249;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d6a2b4ec200063d76feb2c8fdcba979df0bfc2d05d2b8701e9af0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18420722168ec466236e26ccabe86c94165c5a2377fefc14e358fc983;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb1b797eaa1d45a4c4cb069197007e75eb4bc55f85883b977cfb15175;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc956405985103c649bf9c8594a65f78f98117099abb666cf04b9a83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d29a39a5f2f63c96d33dad87014072b1046202783fac508e8ca0547c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2de9ac9d12e8eb5b8e9ece64b41e2e097eeac961c5b632c53b1ed852;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3846d87801da8e173599bed2e86fd1521414ca01d2882eb8c25800d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h130caa26f725e0771b86a8b37c8e860e1e08a47e48203121e30b2e22a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ee5d9036d3d0631e5fc38c3156fe112b96f64f1a82c85dd9505e58c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110336d6468898e0408a2e4f0ab9898c0cde436b0485e805f15d8b8d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd1ea0ebe1c1b458b693425ab9b817319494e9182e43d24dc5eba960;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d097ae5e42cd6791a07d8ce458bbeee2fcf1767a53a1c09cab9a51d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7d6017459cb62935be72bd3e6d8e9790a2b4d086dcfb73dfac376438;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f6a6283dfa8b1f60a49abe5d552b72b118a7d2082604c557e0a30cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc37662946d6483b678baf9a4ed6841464faccc0c1e002a8333449785;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha777b00a37986cb243136df0c4547eca2ad248db6f0abdbab63f602c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147c6bc32f2ef3d03394afdf4b9d63f87ca95b2eb05278dec7fb1ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12df7542e5cd97e6ae2d9c809e5815ab7b358c882ce4198dbd91080e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h971ac3e8cf7b0e3f025306590f2e58a619269c248c895eba97211fad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb9918ae703a75f098115161a928aebcd6558d26a3a40b828f0d071d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7e3dac6e29c6ef35b910b287dc1fb06e82574b039f960952d8592c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd578ad5e87ff94e5674cfd26eb3c436df5a20f90010e876b946757b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1733c1590669a738b36884bcd7285868b71713abd71defb4673896217;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3cf0cad863e0831aab2de1f737100453b56504d23b6a48444cbb6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a6d9f0f7a92c965719bdfc4aace303b4cf7791a1662cb4d63f5b941;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141e429bd3369f5a26da9b6a0160cf31a2f219a4321e070fa98886895;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127991607a30c840580380cc4e46cc84a3b1db21c729d33e9fb1e86ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88ea232c5bd54fe213141849f63fdc8a265355c8e19de3f7c4144acd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf116bff0ef46eb9a0110f5ede8e0fdfca858cdffc60ac7258d739058;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd217aba4707489b3fc47b4a7da10d6fb34672d0ba88ab30cf96365bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h187d80bce163abeaa2ba342abca3b6040c4d05f0cc34185b6e3f18dbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf0c7aff8362bd92d38113f90de9bee20a1a19e86be6850e9808a611;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1139f1ed3924e911ace2c96a0166903d80f5a46763e804723585732c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd41bf4678452a613586c68e5aea7552eaf2478511334eb30ac7540f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c9cf77991654408ad0596ee3f65a3f02b873bcb0b375f15b2507178;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5054f1a754820742aa988072d904d2346f0b604193590a49114ebbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc299b319b22278bf444bcf15606280f95808295bf614d2dee4dce27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24c83feb6e6654c010fd0e23b8c0c7b55fbffd269736fb7ac28c91fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f5c7f6a8f21e83b124fc488b2ee07e8e885e6f9a03ac8683f8cd73ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h249a84e72b8fcbdfdeb1987b6cf690320d3e8113142179938fec3962;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20879f986e71cd32337ae8f7dc38697e01314be3d0449d2acecc321;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1228a55b470b7d82ff56e242f22687231e02fa2d6e6db1f377c885303;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd7f6b79f29a14e07772fdb77a241fd302e12b85c56584be18091d60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4882ac44cc2982180277ad79d77bdcdb224fb081428620bcb6364ea1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18448a677c249f20775aa4794e531cfbfc39d2f33c8cd41e6cd56e353;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafd9f1384e4f1beaa8e2b78bd9d2cadb018d798587618f70a8319a31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1724e62923eea215f394db4535667e5ab733999b267a9452c280be342;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1154bf28ed392601492d50186ddacc30e3055ed42e0ae079ae63f7612;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5d1acd2c9b6aa719efa2d3042c309a362f35de4b6b96629f6676543;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18ce4d48a04b9ffd9ee796030669b2994bff50e980709f0387120bb10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he0e837c703f993225f88a7eb18f128b01810ebd79540d4e63750bc9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a5279942ed2011e43a2bda282df9f02329ff71b259f317021e7f7a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d6226c1d37fd57698424b5f6c8a3c5daa9a6854361c53a1cf8c7a5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188485df24b8cff6af82fc3ef25ef097263e082bef94df3ec9084a491;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135360d6a4e2a79dc93f5246064288d2224aa202f63122c6dfe8cd9b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85afc1b673df27f7a5c53502290b80625c6d2e4315a377cef25beb77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hca8668d167d90fdd7a08d25b93c2b1d0d5f1acfea62fc4f5d3995515;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7a3435929da382f7e94fff5f10be12c38d294c9a35bf64c8f80caa6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fddec67ad2cad053e0a21e83073ea2f0ce0ba02df2300227b896955;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa04e278ffcf60ebfa66181c69f9cce8b72be44c6eb842e6a0a42bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86d5a33cfca17a6c05e8bf3115c5a0c2663735f38bf3899aedded45c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6b4cd83185ae0371f1befd6dc8468bac5e5827ad4e152042430dc432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a3126f21feef864cd2495fe13f207c6f34d7474f2a48de1b6dd672d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed7c9590fec6bdb00af5032671c4ac0a67209a9a8e48bfc9103161a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150ed35add1fb67de1571da42db0f2c2fe2cb1062f684428ad2d98ba5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1680beda057745c765036cdac1b1b5b4e74f947bec3b8bb5a4a2486c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1479d8885cb9fa16a1c54df7a91e3fe667ba086b6c0a641142c0f0d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e9c842c1fbe250204c76c32100222d53f1cbdc08dba86f2667231bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1353daeddb27c8c9e22808ab1f1f686524501a7907c177f012f1ef520;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1296646d058adf060b269804312b0a6cdc11f23f39d5f13e9dcfd7509;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94927942cd56af65db97f3ad1dd7282f50afa434f65584dd491a239b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1674bdf390813829abc0e03a6df8ac2f016be07b72bd9d1371c896a58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h855a5215640cf70f601d6220d1c516d25dc6a83af2de6e432646460;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf63a9048a2e62d54607831d1c7c264c2fa6bdfb129b82329c693c6fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48c0e06b6db635e42c4d992b4010f8d9c7d6536a7f5cf7a3667564de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141a3a38d3bd0022be620647feac631006b6177e0011a4be0ae39dd31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h373f51a4f26231150f494c8f6a6676976bb4bb8483dcfd59f4deaa1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a371c22d112f36e16f06299c798d07ea03c6eb3b0582e513f69b8df0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14fb06dee64e7287f597093fea149f753a4a448f1eac113768f1d07eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f5f4a02647693d11efa6dd1252f953375b25003aa7f9dc4aab76cb71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e80831f7a7a9b08320ca2e182cacc800b133cd3f1adf730fad021724;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he89068c6e19f61cbab717348569e470b6b8faa9400f44d428e8a4d80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f73aacbbbf812805a19cfa00f8b1e338977c21e6f770f76a4650ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87a59452b4aae27697ba8232cc5b8e888a131d21293a0cfe611328bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8d9ad09a38e2355adff9d8b2f3e64ace8f00eb0763784983a63b8b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2be51298550bfdb2adef6b3edcb83c86639f4e3c86ca6f82e71fe6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8709fa3b65113a3b32f307342748e817d35422c3c29b7d7a8267ae4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h841a1eb8b679ac346a31460f88e66b4984247b02ea35d943debcae4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c5e319224667ac780ff46812d3fc4e405a97f7e4b9729421f35e3e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cdc5ca75d249d7445ce89fad9e072f677d969315f6c13babcb9643c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a300d05ad74c842eea6e03048132669e9398adf0e44f899a294bc05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119b7d8e7ac62a21c92a9f2f0ff0b652089a2d84c16ba0708bbcb0b71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5d84897ec795e3301a0b310b21864808e08cd74fa7cf4aac28415bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fa88ec7807901a05bd6a78ec23f499da8bcd8f49bc5b913f31f6b481;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffe0e7fc06fc71719208b897526fe82abf76588c7912ad582bca40ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2edde54975653fac707621566d8e7e88e1f31d277b972d1d0cbddb08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f914417811514547d0fb05fc4f738ff5222fa7768de3b2388ee35c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c28c047760cd9e2200809cb604ee9211654c93abc26f6965c8c8c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c53ddcbfa97364187a1585f54eac0314a5ff267adc07591a35659263;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4cf764d1876c5aff35cd59644043fa148836f1b326d75a401f50e791;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c243a79cedf872b067f80f1e55eeca613f2a3124ea1a44af3e5ff6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a91d14adf82f1685530eb747fe87031944bbaedc7b1de0e77b36e2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb37b4c661ae09e38894b93eca660c93d0aba61811d6b1f97b603037;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ebca1eb8bf3efeccc5a07a7040e2a70887aa8b4b1db1e910d36c627;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48aaeb75d7d9c2e9e973ef72ed6829e93fab366a02ca794f312e3903;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h759cc31e4f23a637b3e3b9b118f1e68da9bddd9eefd0449e818acb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7596feab8cb50caee05b4142bd4952501b21daeb36957a1c74a3acbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3584c70458f7755428965bd59f30d961b20496a87b58a2ed22b1e00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192c9045e4dd2490c4b81215e27fa303281b1521c13723136f95d6135;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7983edf77f6d34899d1a61eae962f60e06104c2c5e99c134e4d16853;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bcbf8a90adb0567a70082f2bc86f73493b457b98f4b1ac59e97abad2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150ef74a1ace8a8198a11f1972f36134b06e90345957cfa69cdc61157;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1374f8c29f92fd07aa9ffbf634d80904b4cb4d364f262cd99fac8f3d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3c1918a369b5ab6e917f8a9f8b1bfe2e8e73738e4fa4f4c1b228eea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a661fab406e5583b8e4a2f4ac2906bbceab57f73fcdaf2e180f8c2b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70e517865aaaac3a10c41949c767b02f90a58b6a5ec472b93cae8243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ebe771e4cd321bfd11d8984c5864e65c37f9c77aa59762aae3038df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbee3a623b431cef1248dcabb4541dda04642f55fcc8d60b396608ed0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4ba4f0830680694c5e16d11d87a742a6020cf9c18355ffe6bf53d4e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h154f895cf65e44d0d309469fb461169ef43fc7b5816039e9465113d05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he395f35eeceabd725dc425d93cc57f8c1d22a896c95fbcbb773d6c2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19522fe0bc597d07daee1646044e9f25e82df76b67d347cc9bf11ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h186ad6190c926c89d1707b0d257050cf8d42d80960a12a2eff49d46b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h464172770cc7aa6f3e15dc9e1cee3f1d6944ce98debd4b8b4fd699c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e389e5766308b9659183e7b0b7ac4f529fec2c7890805434ad28267a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f55f0e1afd13429fcc906e25fcf556eef67ef6408a674fb6e19411c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c175eb4d1f58e1156f25750da824e4706b6e6f4d24730c7fbbc673;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf0a82a41c5cecfa77847cdc69406c9e34d23f1b488eeaf52e59ef43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6260ccc503d31b483eef3d1551ddcde7865dbd3b89ace813720c787;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa88bf5e42f031a94647e682864daf0060c36310f300ffb14da61a06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4223fb7f1c6a7cc25d4008685b98cd7b2fd7a367095160562d845fac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123b08ba51554640c5b707c55b839e409320ebab9bc4020d97af6b440;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3bd92758998047ac245711c2b8da8516a04d32036d9c9fd075b4aaac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad6c95305dba4d237f5c84208111a61af47cd4c5b30f89a18fb6b544;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd8e2482f98f64409c03fb51d045de0672d7a2495e7e626d249b75a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f6cb3f3e782c404ab7ba142c9297645efd5be0e7299035a6156fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h365a7c7f026cd736a81328de44523ba41bdafa038df3a9957e97c062;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdeb618e58bcf3f6c531329fe9361bb58306cc39b5e9505b55ac1d1ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2b854b94022e69191fcd4b8afe83d379a9ce508067b1b00d804d56c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a35fc3bac7b67145c9ad5bfffc21bf6a201dc2c884a0fe771a2b7097;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171ce36b056e30b498ec84cd5f62efd8275f24e9f9864d7b975eb06df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106f09e6d8379860968b65ba97b8deb9cab88151446524cf94d3d8de3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f3c4af076e90c51401a82c5021cae87de20f73d5406234c3b0bc170;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a3922548724c64f490d0983053ee97bdbff406ffcf34d90cfb5b366;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf886beaf51b1633a8237ebac977f1a11b453a28c303e3e7fb57ed854;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4ff771a38da154929fc1e50d1f20addb026fa8c016e970611aa4c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16de12b3990dccb554c6669051f34ad2f8772f62d7d334eb496a33e11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h104396037cdeacafba1d6fbf904f5f884a99d07e7e89d1a25c047e78c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e512457e4ab3b423d6e8cad81e2b0a8cd38626e4c603859c800fa05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3cf130ceb4152e8ebff9947356c8a9c3de10490fc7af0782c414fa2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195d5ff841d7b2469b9ed75551fd9ea4995f24ba7ddd8a1009094f028;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1726bd44b6c3e327cbc7119b6da44730d98ada0952886a620f5253c49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5006ab84255c0a21b72575d525be9bca27fa3df1716b9ecaa8b2fcc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a48c218eda3a4a36d59f46f6094080e8d8ef2ad72bcb76f85bf11ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b89a3adefd8fcd6d96f562cfda7e98973c3bf3a8b4fe600f928bb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h559cf3c7086699753955021673296e3866d30eb060d7a062efb27c17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f060f52ef96a4b62f65c5174f64251d605a98255c6772f28908fe89a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39df4d6c264da5ccfd6a5d6f65652ece83946c1c0529b31a1eb351c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13eeee800c66bc53c7a59fdfdc4145c3803e14d8223e7772f31c3fb57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h968b7d22422b24e58e7715038618d827a34e1b66191e97adaaeae80b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ed6f8b418f37d5e611bc4f683eee335965a2ca038fc912412fa2e15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1663fac816675d8d13bf8342fbcdcef089af256a6d049ac19d43a26d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3a54dd77501f68be778be68b2c5c069048ce3345425ebd9a496604e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1446339202674ef9556adfb0c21d055c698890b354344345f27d74e2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92c38216f222385023e9a0260a0eec4442b849a72c467d6e4e145399;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h179abaf9623f46eb14a7a99344c8ccfb19f6fda291101c72b7da32492;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc19a64425c8a7d5422db2c44331c08a0bacf0420f61a87526892c69e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18cbd46960dea336c96b27ba74bdfb97b0523cddb2644f3be1a84c280;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1989cf1aa8ea0a26792f93e744155e096203d85cc52e07b0f98f85428;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed2798c2f80afbcdc743837476b5aad840aca424d5a30c0b228b83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8d4be4de34367e007eaf7454eaaf1c9aaef9e997e91ec0cdd39aa74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b760e4f00a799f49f6d86cb9d18e0ee4372f12f28b1fb05438497ce3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5041211b400135ed1d6fabfdcb686cb4409ff599f1208c35bab617a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3f76ceee0e561c3ee6235124ff1ec381e21f6947df12ae5124b472c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h522c348e3e0b39199f87d259f45c10b0bd9c533cd4310bacb9be600c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135812c4979a6b72f4d31bc75a543735d93ea734a620ef51d9f847a26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4f62ec0cbed91e80a8b9cfc9c0d0a95bbbc3f30bc215440ef74442;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106d27983d604c9b4d927b6e2b6fa29c3240cab169e81eb21119338d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haad2d4db1cb2ae88d89269ecc06f395a4a31f2884096fb484bc46a53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4e843fbb48a927ffe345ba2462b753e97706d1731b5f25dfc6fe0188;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h165cf383cf3e3bb025300f7443b63b4e3bd26a15f15f6ff0b56d16e29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d4124f94009a70aab837989e5eba6f24ac5546333d4f97b7b3cac00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1871acb80003267029356ccb46848085fa5cc812494bd6bf37b68bdd5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d5035d1c6a4f4aff92bf8e578eed2dceac1b8c93364cb2f3cd0f827;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a70daa42b0704c75ceaf5d2b1442f1612085be412abbb204ea38bc21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8fd5cc3a824465d817a7862ef98258cd930b6529681f80a21f7464f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha54dc6c1d7667257416ebfb74508002451db58d4ad2cbb3bb144fc7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdec0f293692b364e9254c6487b2b2f0aca3781efcaf8ab17023c1cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a59a15cd5d8fe32cb281ee25b48c3f2ffca9cc7355764f55d0c3015;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8cc4e0c3a8a0f96ad3076acc503c12b97df8d38b0dd22aa1cf85493;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f8c5ae6918393f0834597030dac314f08d9f9b3addb54a218c4ba83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1878314516f32d27425a38ed30919986cb1bf0ac44339ea06418e2fad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7336b71b36d72592d44c920c54249dd55dbf22ae880431976e7ffb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192a823a8cc427d81f94663892cea0250be0c3015a118c541f6eab11c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7d47872542677cdc4ad65cbed8c18f881216bf371b26014d03c559e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd1b88ad91550bb2bb860535e5e4171862ce6c6a76dcb2d762e06aa2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h408e5fd56a5f583c26c73e0fb8997db9343bec8851a5f5cd86b9b4a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ab667197938a4b2b9c6a7141146899644fd265b03af156e5d67f307f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec98556959e77b63ec7b43644f58ac8383b631119b22e61440b16a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1302c43165dfb6f27d7ba83d23d5daaf6762492916e0337d61a17c782;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb13d126cbe7d8a08f573da6b732c124c5370aa862ca5c76c4eaeb948;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0bc8c4c0cea65e9dfe1b08a59229ad011fb9a8751dbeadd4b70381c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dad37167025a5b98fc47e07a4ecd8ed98c029b711fd84033a352a194;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a005794e9fb322950b890f50b0ed9a6194c95751733b2566d0a35ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad04a999847dee6c152c428471e0da859397454190c3305600a98144;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb85fc1161838dfbae37cb27bd467248cc9103ca6ea30c20b7b9f621f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1605f94bf36d608e0dd497718cdbc2baecffa529f128201e384c84509;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a9316e88f53008bc0f23f2c97826c25e34880d4399b93b5baf19b6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26a4123f2fdce497398d067d992a53af0de1822b10be68a17354f282;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfbc40083392d635f14422b90f5d3cca43972e228c68a1c6eda6d4f01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d10d40f0d88fe8bc872f450a9e915fc390a9e136184e26fec386f42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c4a3850707bdfa5e9a94def142dea724d52030d4d3a19a55899deb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e3497ba60f7ede013d825cd8321cbe1bd37f0b0ef4ca57c95b30f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h107aa7113ac799973bfa04a68155566d2de73d2d20b34df32ec3e5311;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147aa88b0c7f5631c2671827147365a6ba969222f501b2b4938d9099d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf38c288dbae496d108a6b8cdfb3311a4aca623b91d17c6597b1c8c2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fd8db787826527085cad7b068c2f4255d8cb51a918049f3b2483198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1696f6fb7227b12ee452c7a5dcc13f687b00f75e5defb2d85e100c2a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a5f81e76f6b9141100c291b7ed751bddf4691b659c8a4b960382327c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb9c960162cf000172b5652a3dff308bcbfbb3b5deb44f6e5034ad02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he63952db3f136fc66502cd07545d0946866b05bb645a4c408c76636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha91f22fdf4b873cfd90affcf8e8e2d00085a68c3b3762f31ff3ac2be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a118a95d6f39862da45cd4a0b4556ee5b88f5f8183242d5258b1083;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1588f2aa9c5c1cea85e74e136cb20ffd56d83d219a8a90695526afa40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb971fa6ed9ff7067829d6f2a8a102644d83b80ff82c7c1816ba427cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1320795292cedb6324bade08dab228636350d52192eaef6e936a29469;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98a1d728a54a7975377faed81b0ae75186332b369e5e7d78eb363ac8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2df8239cd21015126223d4c79ed6905678dcef58e88228fb90ed980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6eaa4f46acbf555c7ef83643a32218da180b3a82eb07b809aebb863;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he3352b5384bbd117086d5bad6a23e3ffe7c9bc020900369727594fb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a039ce29f6383563d42f4b28e9dfb6eb8376b377716723d127fbca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf37c48ceea7ea908b96905ac59496eff45fa08ff864b461bb4a2c59c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h50173803e39604000fdecce7b6e9906b4f1660d215a9c1b0ecfe8033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76260f6d23595bf9d2cd3058562a3e31041d72d01780bb063333becb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0b4679daa2d10cee23022f98ce4cc587ac37c43b8b4e240b9fd0870;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf1fb03446c5d7725b45bdcf74dd94ebb71655b464f9a25e4cb72a8fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he9ebaf693691ac704ad60b4907f34e03de919a87d3455a6d2ffad0fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h22ccab71d5691ccc9c9e9c33d4d0dc17ab4b7a100f451e48b06de7b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153e17f657077e221fb87247bd0cd50eb83688d06c6f88fcf44879c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc07788851f213c63c6b03e0e9ba1f559ca1834ddf6c40f8ba5dedf29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h502af7f118b9f73a1c062140a38cf84e7a43f143393e53f101e4d4c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33a54cfd2ac4acf921a50df00d1cf84b06225b0ef149025dab73bc0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde5741d3fc2daf00441028c0ad5edf289fb814971b9fec75cb439233;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d35398c1edcfdcd9eb577d89641355289bb200797b261f866199c65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131990e948102c84923f4b048268c6f45b256d67f1d5d326a03c17442;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131d70d7f19fb68e895ef2d5256809ae7d495eeac1193a484915070e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11402e77f66e8c65a14c70678351380b2a6271186e248cb49254128ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cba358c38f376b077376d5d1ac58fcfdadcb73b71362602efc90a4e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb8b58f898641c8d934da23c3f467fb220503fd597b775f3f8ac0fdf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136acae3a3b4c98a519928b396a2557d59c3f023528fd5e3f79ab15be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83af9a780d8f9b5ed7a1ec1b0461b8e5e09b3720ed4a8f2329849bcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddb87e4ba03ca6e15504fb25a77a451cbc460af6c5450d6367b711f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h107314eaacb5cf028b3e5b1505e9491f1a6de8322f543e9fbd7f7e031;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdfbdc6dd40b52e7405b4d4ab6d19c0f367b94dc508521253bf8dd001;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c1bfb3c4a6bae35808f4134fa6ef40f320d6fc338e193f539ba3c45b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cbb9d28ad6227ad1905a3fd17941540e5a3e105e2565ace5cf5a7c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1acda71da31edfc06bae06608ce7abef6859d15628154ad4d8f6fd789;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4be7808db0888b89a95f3d578ee62cdd353df112ed4210ee1d1e928;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c278ae819042d1d6cba65f51af7b9e82830fbadd10670eac6793bab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd34cc71ee66fc10648e3f1b64d081ed571ebfa262de161f29d304b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1031f1336ffa1e811cae9ce54d50e13901584b652d89d6d84584f6b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c46640ab3940b50aaf120757851a3cce24515ae069eb978f22766583;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha271b75c96f3923abd269aebcdca129b9c4ae1629dd378f0c65f8727;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hecbdb53585306a13aab8b54be6ab0ec605024db3b1e56ab1c58daa0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda4ffb096dd5a39748e2e5936ab605ec92a16d051d0be06c7cfe2d4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110137c3599e957faee7ab110571c8a14fee1ee08483ed1d5e023ef0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10391a6ef695c0c88c0d52de1b113c29bd01a4bcad5e795f8248eed33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha18eb95459a685fad02de1b59d39e69007dd917220bf9436d89c1beb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9be80549e1a06fe30b6c007241280b9ac8c41f4f0ea0bbe8e9721bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16da0b3645674dc9bd42e04c27cb9b248d64daa3a1a0e88ce158c8c20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b751b50b99e133194bb8722c764ced867e0d9c8dd989850e1e33743;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e35c6770752c8731cc87202ee6120faa71413f43a77798fcea30b7aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf69da86354dfa91c3d89270e0646bcb9510911bd71623d46f9264508;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86a3847a532a66531937c5dd6e9de04edb34e85210c7ba20821fa932;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b264c7fbd8671fb584cf7dc0f00df41e6ad2daa81576796d9f575467;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h182c66578c8acd69bd3b1971c9db31268828b857b07147c188e22f3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b5d853fbae709ad9c86d27a7e5e1064c4c733c9e3c7124de0c4a508;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1efa18a365297af189e0508252db945710b0ba5976206c45515b72e05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h161a0b4fe81e97271e0618e1a5f9e2c2908193367911c9c020f95207;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c251647e7c0ef4ec7e3de0e6762c5d06b0df49597e742d22a3969b57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb435a578e8c553ad275d194abd740c8a30e4fd0b261c37ca62d3b4ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc7f50687cb1adec06cf03f44a8660010419654d431554aea4c07a7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5340809073c060da4330c8f664ad89ab67537253ce024d2c5dcc01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ce79b418a6f393eeaafc70f725c7168287cfa45f4ccaf54c0b4b54f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf3313b916f1f729395a281a7e27662d311709547e2d6f11d46bce884;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f644d6000629156528f373285af2031097cf18d75ad609ad43cddae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e7b18803f7fbb933613d0adab4cbf923c064a146bc83c75e8a1ec8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101648950349c41edcc104712a11146976126df424815c1e95c92021f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h170e63d2418f35bd9d7e90e297de335c564484d3e62f60d930b28c437;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4c2d2da5d5881c89ded7b59d548b78aeae62df8fcba7034ab7223c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb99e0a8b701868afe94dd5d4d874d48555dddd5d2ad1a0ddad9f8100;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8004096584c6d26fd3c8386bc75fc45aa5c63dc5ca4f5399d3ce3137;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1b7e845a37772e4445958ac094bc6f5fe55ed840a39e343e7bac9a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18e8d2c3e7409bdde502bf8791690727fd6a3e70adf7dcff7ba7e614b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10780b725893437b7229509aa7a50106669768d4a2be5af5a78b28379;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1a70e102d86b63455de50fe8b665b5be8563db4e73c8185b1d1a7a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1905ba4e5b28362b4ff10a48ddb6e03fd445cde5fb47ff737a68d608e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5ac8a74cbab682e832693df9ec3173c533465d485af03c9ace6f4ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f4d22c3e664dc3161dd2a058745aebcfaad6de73aa454aba22ff06d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a53b27c99ef38badc358b2745479a82fadd4fc9206252bc520c905e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6d22e1743055e40daab34c675e3c95b94c435930dd43e57b58f07a85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15afa1851502f4d1a9b6063c02eeca838d6956b116de00e0e67b08a80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea9b7ecb38e4fd483ad37fbae0b7d4e3dafa71d57d6ca6c21ee761e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75295e0eebe2c1e6960cae43e4f196f63f5304bcf07124ff31c4f6fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd058ee60b236daac3e2131dfe39d6945728242dc9b3eec748c87c1c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b0495b22e49284d818699b697b933e9ddc3fe9500cd877d8c78c365;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d8516721ef5bf38e9d1f7f1fb3c1ea7bd600a6972790d280ff6313d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b5c384741a1e20f16324db61b597c2da83874f05979a32a76446c92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157230355d77714b8d461d48b8ed9455a74694b2f22b23ee95c761be1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb444088dbacc61718d526baeb93b7b002f4ae2ab7f6dffb6f0d30f8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h166159dd3e2b881eb0473252b82b7f6546babf0e90383d5f57ec41a1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b38e21bde1840ffca8dfa15d0d76ee5be406b3db6fae0acf9605083d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a4f90259261d9060620a56a728b6c81526c3bb3eec25f53b01325e55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a4234cfba8efa75f53b905440f11edd9c2777571820eba36d8b2c20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffb24004d5f878aa5cedf3ac31e906118d5f2f6d8dfbd9489e2f50ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1872efbec0f11815d6b280f57cd7cfd07123f08ef706cc9f929767e06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7b5878a95e011335b4d92460f6f3505686f63e34ca8a203fa6d498b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8c2071ccdca403f6229faae921674d47552f125e6306c37b97f6da1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6c652d754d860c0b79ab623e10ac2aeb29e446bd35290bb5836c39f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9be3cd271224bad8837fcbbb850ad310c0b7cd274a956b9278b3f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbcb3ce030831392ab1b0b7a938996a93ce7aa4de274ebbd30ad3d09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e8d8e3930f1ed3f90a16c6797a750f533d67bf10c2eb3665b35039e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c2b18ad3e979297d2407f381eb88950fdac58c7e352c475424e382d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135b3cccde1a10a49a1bc01ef5d94d10267c6f2464e5db6ee5502012f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101328ebe275f2b39972b229193b2c5701ad3d21423bf4294e5467616;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7c0bc548840c1537b287ebf5d4e929d55bf07d9b59e022b00aad41a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaacb0b55a658a721ea1f4505a68428db78145602ea8df71cde7e5eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75e941792ab29d0834f4d98e3a6c3be452d970bf99f9934171053099;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76cbce0909b24fd78d0b7c2759fe45a7e5b2a7b5f7d16d0d3f0471ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3aa89e15be0b6863c1519d0566a33dd3b8e82b79e7eae3d301e99318;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc94a7b4a479862f83406d7aa90b94027e26af44e1e7b4e67eebdb218;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3605b722d2c535c9d41b8b203fce88e470762ae31fdbd6822ca8085;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14696d7a1d0f3b5b42e64bc336cc6dcd4142aee62b8aad7da4688a8fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfaad990f4be7eb6a260438d9c46935faed700b11f50b05ca3b6c83b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7d22327e1bb4fd8cfb4604d9b68bc8223e9858caab9850ef41365d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd5b88d786c610690801aa9f4e941b78351d752211732703b44cb603;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137dd9bf7822c722e50754b960f9dd82337dfbceae30c44f0d832d1b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1793ce50289c27cbe7b0a416785bb575ae4d49a5306f68ad892ff974f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f9af3b42c6c67afc1f6ce5ad25b572ef5d30f129601c622f25ddab9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7038374bd2152e497d394a3f9a6838367a6c1e7a607c5bf00eeb86b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbea8f72ed570da38e042adeba3dbff1a4764f5f5d29387c1f2760abd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eaf72b151a1c07f2ac8d1492753285e45f42100847c62f0859dc2cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177f31596d246d0b1f5a59e23cc2fcfd4bb7f0c5d1e1f025b583808ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he543266d2716429b7f7b4c5a12d8eb54a7a1c6daf56c50f924f24bb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf01aa864f669b19c8ecef6e8c9d6801afda8a56484937efb919ee20f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39fcb9634a6fd9aa2a8c80dc022d399154906c41ba330e860e20dc90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3959d31f91bd00b362c119288d0cb81e45b3dd68a20f6d9e3392123b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127207b984b694fe94e2be6cf518b36e83178c7e5bfd3d7553a30a99d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d51530ce354eaf651bccdca893e01dc7dcae5575232fe967766f6163;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c7e25904c1fa9f3f016853bd66e2044a8fd662a27a250ce06b8bc8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1afc990ade753463fc0409236ff4b5134d2fd31bab8385ca4d7658026;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha06f9ba3cf642cfb139d6980581428e670969ad069e1561a33c031cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h84bbab05b48bb7fd35b5cf9bb18631477e8184e71338606e406ff845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1223a3c2657493bc1403a38a0ef5074ed4e6d3851b4cbcfbb0de51495;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4924bd246b055b22549213fe8f0f0cc54d66a2b69948f1fa9cd3de4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f49195b73b6fd39bdd0d6b9dc0698bc208e190de455ab888f6bb126;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15bffe374e5e0c7091302d8d568f2662fc906d85c26fc8656a102209d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f41c255f082432a81df01cd8897a0bc293e8d50f093fc17003c174b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e4de9dcbe61bffee2dac602526a32be7a24947b449eb5d908ec0c62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113528a1bfe90e5bad86b35ac4330d1c9aaa18691f16ef32c98885a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d29dba319364da626d14230dc10e805ea5d011f3ffdeb3504ec2a2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94174f96f72c62a7f1763922a2983c03a37f75cf8fe34e11ebf04679;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb5805f64e68f1c0e02432d755cb6c8ed7bedb341bfb449e996fd1e18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1802d10592cc0803b92ba9ff4ecc98dc29fa4fe54f33d2e719d532698;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e545c2a0fd248d15bcf7cab83d058ad704bc0a9998f09033710dc705;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b988a2cd9fd0547ffd461f187559c08a538a65e0cb8dc83a9937c9d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120f74f41578d120af40d813add67ecc5cd1733edf90ea2e77de2fe63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95151282bfe9c5fc3bfcf3b0231fdd7eab58a775147802a10a2edee6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0db82875de86c791d85ef9e18aa584a5f77f7316c8a0751315da74a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14539a128f0f816b4e036eb81248500f5f752813f00227d5a0e5206c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a3a2ab4567d9c2fe63529db05c6aa83e7a99f6b308b141520bc24b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3de03db3780f979dfd33a2e78a552f18656767f4b6869b02caf4555;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff84323e7caa2d5034bd1f7c3d6a0ae55537ead5447681f7d9802467;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4dfd28843b9bf3d787c2ebffd8c87a4f86478f6c6d6308d7a27878b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12fbc0b3381a4ad14589f66ea7af074ca54eb38926af5f276658818f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9568d9ed4bc3d4f81c7d3f412883e65d76e1877271349091a10718a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aafa1c2c79a4aaacd070758404273a095eb72def8216203cfe014c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ed92c94ad5bab3436f1ce69bb22e7e533aedf18d9a89eda4ba87c73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ed0d9b7bfdee2c1a32d32c0f7bbb69590d49e73407cdec642840239;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h166c260ffb357b0df72d718183643456490ce7ec48e64ffde3bc3b6c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd79d3749ab2ed46e6ea527c8ea157e9d8201fa251f00e669e91d9a7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49661c163ae7beb464bfafd3eaf38c33bc3622bbcb4f51181abf9417;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117c3cfddf3052da08605f7a57633b288d40942614ef0d7309917598a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1722a84f30238c86932c675c8250888731bbdeab214bbf46d24a52de7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee204299560958970a471edf77cda6076eb5ee5253311a9e37585431;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b50422e46f96d3ea56b52021569ccf6212426821b29443a36cc9325e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3d0755e86cfbcee4e38f1033c514c158a32a45fbacaafa6c8b063e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78dbf8949a9a8f279e211147d00fb2107818fa138001b50d415db147;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17da16b345ef271b98889b8ceb3d4c9a2bbb6c958400019b0a48ec695;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19be0563f83716d4179df733aab8f241ee0b880d524258acfc41306d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h857c947fecaac0780425f31fb29c93de24b365bf9108810c7219e24b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c2d5beb8a23d1f062702b950145683ce5eeb4b8b0c183a7cd565121;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17eb6c5f2f01b049fb470cf8f9d57147df86ab3b34ce071761c3b081f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7cf9dbcef6ffba765b0e96cc45d20448ee9ff16a40b70dec523d1d25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ede6b056cc1cfb3c7c1388bb58b01200aadd5d57f0ff60cfccd6056c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf55c097426d6d630648588bb852eed75f4c29e1c4ad594c072d8a687;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ca30f5582182b1d47efe9b86b09733762e6b67b12a91848e233b742;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h435b3e47df6075d47e69e45207e3c1fe514abd3432e3be828c519415;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1badfd61b7c319c6c9cfd045950872849269cf61535469bf42fc629bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db0e0bdae2ae597821519ea32c0eb3d2dad6febc3b6d757dafe3c1a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb234d6eb5993e44e47e16ce68b43dcc82308897c44f5bbc056797526;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177994cf6e79381441bfaaf000c6ed5639679df3c36e2e8604dc4788f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde1109fdf98fce046a310ea331ec5e12b3b4cc5dd9d3507323d632b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9ee019c312a37d193943f1f5cc02f66c2a26d27f15454dfced5a244;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e96330193817c18a332ec436fe39efcbdc9796df18a90173c2ef1a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81de5bc1f15a8c5327530b0d8a65407d48c2160e2081f6efc90c8cc1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2b40e9d470282dbb6e7b471bdbe52aeb1ca0a54972cf0865a556268;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a9f41a6f79d7c785950c037ddef1d617bd8ecc9d19e2f2fd831620b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5102dc6039eb41a23072d67d89cd85b63be254847a9ea8b4c259dc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f30ae5fa40430429a9ae94e996e77434a4103be1cfe32d4056e0110;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169ffb1f7ddd1cd3c416c422e94f697dd70a2adce3390ed14a2b902ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea546ce572e29f5cee34f8a4271187d488061c6113aa97819e0c0ad3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f52582f5d77c35311030ed4e5437c6896156f6b44706ff00e1e24564;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1211f1e8862a8adf0e90b73c92b2cdec58f09cca6c7986fc7b49e638c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b87ba4a691c1fe4562465bb85f9c673da9531ce550dc566ef387c623;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h60ba59c6be9fccf993473bc60450e270bdb11e1b5f83bb8e6bfb2cb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18ec6402c7da2767e61167936d86c247e672d04f6d888d1013b44708f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a04a9ca851697b90a6553184cca4fdbbe09abe0aa87d99e468a9d76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92eae6c3cd06cdf19b8fe9f6e30088d8aed819d6a2b6cd8d1232358a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1621f5dd1f1353512a1dec40c112b611f4c8418ab9ff0a147724ce6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b85472a0e84346d48d7bc33ba6512aca61f4ded2b5294ce0f370be03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb9148b71cfc20246e7e6e544582029a4f2194e1e14fcc49dcdb5fbd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1823e2f1a34b5fbd50cf6d0e60fc375147fb70b04c6cfc32957ed557b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haaa91a5da707a44151aa22cfc17d4e53ed560a4061231840f4041697;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1381dae9c1fba7d6d494855725984c3e67197be62c27e3b042633e751;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db043697731df6d21fa2064529423209249dcc78dda1e1a14499210a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191cfa2213a6934bd56d281bb459cbd98b2ff2d18a5678c99be242305;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16602bb12c31699a88662e7b58b0225d61801fb40dd231c402fbb7f07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1148893704e7f36a6a9fc404f0824dfff2117bba94c465dde05b9559a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h69e3e6f2a76d8c7266c1c2854069459b34c64ff5297f5467809f05b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125f03c58cbaac6f4185f5dd2c6f028ddce480649563fb57c79802a5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131914d21da2dd5f9a4a2f198c057c9c098fa34057988aa9f99bfede6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4413bb3dccb3935b67e73b3022832cba5316aeada3b9848a7de113c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca191f97c9c187e6a879688a7ccc65ead475a6887ac0276de59963fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf530f47c9a866481528268495157bc91c959c1ae3dadbc2e12331145;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec4f4845c221ad38c59daaebfe62af74dc6ccb85007311a4a75f4606;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1374fb826134fb7392bd64ec1cfc7713795c11555a37de0aacbaa4f8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h128dcd2714f87c5e3f3ddf9acdc91e861ee7a0ad9797e2051612b6b14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d8c135a29bbcee9a6316b0b662817c67984a8c1b0db9b449facccbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7da0f6c35ef896e0b0acf1407cac1a10229e328bd95559187b4949c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6eec18b3e31db96985af9105e80be84fd3dc8dfa482a029d1410b9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd316e4c1d64b4aa1c7ed060001949882c3e0e44290b74752bd6eb61;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11703c9ee861a0f7ecf387073224a86ae29b60399c6d636ea973d01ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13332eae144b2e8fae7ae299df3a629bf4c0d9b33c5312b8acf0eb0d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1448bd58e34e4dce0b592fd16283a84404e48d28dfcf62a9840ea34a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1415bad0f339d726f4876b8339f15e788a1c5402d1a7b25ebcd48618e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126dda83748babec3e2aa8ba5e2078f3bba698d99438120eb8ab7ccc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff7eaae69bf22e6ce87439daa24886fa23d44dbe75d349cabee2bc63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b5ae97aad616e7781806ba9431e7bfd08e89ee8031175f148d0cf04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd0841c2187b5356b8a6401317c78d9bd94bbbb45e29581483599fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h54c45055ebf7b9645ab91157a6deab8187efa076517ece9a4ac91331;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfedc4515d6b4e1b66c7ae41c6bbf24c7fb18d08725ea25f06364622d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157d4a1ed01f4b7ec32efc7d9fcaa573f8229bf4dd785c3999f7497dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h504d2fe17ed01e088e0319be99d42470df985587fd3c325dd73e3f5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3bc0feece9a7aa7ace05864d595977e455fccb024bd619ce8a35a680;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1800bc9ec9f98e9bc316a692184973ce19d8cae80ab0e7330c9d1c6be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4838dbe4e5f113eba889db7f8bcce098a0a78ff295213cb865d481d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba7c954f81677685de37301d44daddc8ca52e056269deb779534ba62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d7f92878d1edc4aaef8ad65156071cf36a573d5e36768b6e60f69030;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c572f81ac61dbeda04a3084f537eb09ac36eeaebb359acc08f54088;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63ae1a219dbbadfc77a96e349a4ca5cfb185088d7ad7fce2e297b1bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64cfdf24dc78a8036bda8cf5f5c5f6de4fa4c20019bd29bc2a97c51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f12acaf6c044fa74f558e20666bae43199a931a136763c8ecf50700;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f4a2f410a124ff857e11b4f522322f00ac313b83497a7e86ac3783;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11460fa56ae98160a067837f66f8b7322fab105576e30928f8c254146;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h144b6e459a11d5670985b3ff1cfcd5b13c812469e9456d7de4a8e752b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had5721fe271eff904ed4ca2a89f80e65ec765c1886020259d668676c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3b648911aae4fb5f95f633661a9f0207caa33d68e41134b1427b037;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf71febdd6263ac9032013fa112fd1e9f0750fd80754cbc60e22e3f70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he74f76f49ed93dec6b2b5c2efa9d24e3542bb8cbbc0d6db5723374c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h227d9bbfaf0b020734a35a4201e5b72f5ac44b8021cb70ac8fc73c4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ed9b21733bb070e8b8af74f33da5334854109b262caecac3ce86743;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h73d2a7f094e03e7c07edc741a468d15a8af337df05e78753ad961d57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h144e71d468815b7c6a65481d8d34300e41ae51a58c8b48523fc744a8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9a72f339695d080047fe40b7d2307f95782fcf40639200092a732bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a74b26d7dda9236c2431708b75d96188a3f96ea7d804ce4b9bb8a27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f979c9f21f5c2d371594e210212be1a90925e4988a289a02f6a9fc1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142fb85be5ecf5d404998473b67a7a9d82cd496f9bbc257a704ea36d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e08a61e7a96c3cb03d240070a5cc0bdb5761b8ff4db9133ec6bf4308;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he681be1c6afcb07c48e134aa2d3b01f5f92b8678865261bed1e5e6ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19cb4d52ddbbf23da1d20e7e3b2f58ffc48b892a327f8df368be00bd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4e9dbf01cde50abab856df55e9310d7379bf204929a8c1219f802f0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8ed195ff003653ba41bbd868b0bb3075464b4797898a6c816f69886;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109b2f6c71342f5163bd366f29d27f366c2032626569a3383d4864c19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87c70489c5418761fd63494d71683521bb565722852d4d09dba6307f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14625d10141f823c1b53f5e64ca5281cce9ea2297606400692817108b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7e3b1c100ddc5a3b42c67ec87e134242f09fa22c592bafffdc7d8a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19502b6d9ba33040733c0e62904c2b7cb5289acc59faa7828b90f544f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4495aec08c7cf20377300bbf11b6af74856042d35a7ba95037f7e8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da48ba11c72ac2221e0fbfaef99e9ad0d9f6c90dd056bc4aa0e59d57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h751db70d332f6314f918c9365658886bbffb67648f7b8a4fae38c23b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1edd34f4dd684c2e1129c527aeb9dafd5145ebc09ca242c2c0bfcf798;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1104ee2998d4968c599c8876c9ebd9b39369914d9b192c03d3a842b1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h581a3a3008d13a6e7f8a224fcb99bb3880677195cc25bc5ecf80473d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59cf0d8493f5b29c6610eb4fb0045a45dc6d28e24ac764894e17691b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ca7e335868a7505a73e0830362d09fbe155514bc686547f4a038e33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147b0fcfc6733d0144b5c6abae75e8b36725beaba5186f8950810da77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h145ab4a4515d358b5a08e0ea334cea289e43654db5a8dc1919eca1e03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76a1fb1092005c2528201c5e3dcb8ac801fa355db9d5bc6fe4e6599c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a128059f1d995dd9f08d6ed270a6f9397fb34e30eae34ce6f5d8b0a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6a8dce021253304b8534f728ad2cf5e0c9bf1a53062883f1c04fa42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75fc1eecc4bcad3b4e631e6c9a25461b9f9dd7f9ab1b1db0a5dfb579;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e92752a0d1015bab9efec956accab7d9262e3ef1d23bf64e566f4e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf98c7666abadfa135863f52bc0defb9fdc0e3d996a537a6bce308c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63e76085eafb1f5669bbd1c2e2c37ce78b014ebffb3ff5cc610ab652;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed1f7156ec773591ccb5b6d55971c3f42d165206ce3225773b3501ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1322a2276ee9bfccd2dbe3afa5a612c8bad606e18fc6466488c2cfa27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51588e5f22679a693de0016d5d22967a4d5f61a2a29c606e88e70fc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1157af36274a459d80fd65189a9feccfc247b92670a02e0aec87bfb35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea9d87a124f5d73fe4875853c435a64d3a7b22e7b22fb1a351c6002e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7e1bb249a77c98f38fba11720e56bddb2ff4a6344fbdc211fe8403c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb13c0f2c0109d5d0d037cad16dae0290512bad42ac4ba3174edbac18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd65c2082873df8e81b7f715fe78653988ccdde3a300111b58233eb3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e32b4f515263ce216ddf17becf7f9c66425bcca83a1ac5981bd18e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0cb894196ff05dc8be59238b723678a6a27576fbf36bb8e09a22337;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101d27028bbb70f30df2a93d1daef96a23fa9f43d79b2267e1e97aa13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fdf218f16748b4cec0dc5d8904d63eb183ed2419d0b20d56e007468d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h71fd5506d6806d1b72a385a47026fa2c33e21bfa67d01d15a8e0c020;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h626a01d17c412e8bc200a3bb76ce53d45023fa8b5caeac881d92ab41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f517b5bf113424feed1b31966f763e48e7303b0758203bcbf6ab5677;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdf16695eafbb6a39928298522215edcaba3fc5ea8faed5bf4ef066d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h676777958e28caaafda0a28ebada8d1c898b4724981110a90a767f1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7c078069fc648156abbf5923e5293b017440696ccd06113e8ac1cd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6260d5fbdb1fe0c33adc75f0ea5a926a0f2192011a86ea9fcf31293;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d4b6782925f64fc2f0d0d63ab2aea549857780232c18d93f1d05fc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11021e4a75e8eb120f1238758034e2d9c21773fa9c41ea1c89ae823e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4962a0f810d4a7354c73d8fdb34f6119a682bd312e57851fed51598;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha444d8d3d4003866b49ad4f468c16f053f3ca503001a78a27cfc023e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f723f3727f4daa8568befe359801a711cc90f9b8f9dcf161374becb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6cf1c6b50d962370bad4ade86fb9e6da1a27b80561cf0092de9288c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131ce4613611110c65468e2fef4e2672b7985c5df51d7d3e3f40a09c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d8e4110288c881d22e927f5e04de51e85f5ebe7401a0cb76d010392;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3ba4333e61558da1bfa769645f4c9162f310574c7a38422d6bd5503;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39c6ecc7ef82dcf8fe7b8c57854627a06f75d2630c3611e0672865aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha928255a4c8e475974337e4a3fcf32b484eefe3548acbb7672a3df42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cd9bd0139577bfea74a3249493e17d7786f5577e5ab25f65365f56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13359f7f3f3f64e32de1aecb553b39cc1ad78760728147f55203e15f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0504693d94bc0c9387111080399768a8171f00cef16038161b2e62e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ad31adb6c3d23e0905180674774143e7b57db56ab010a214f809cef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd39d8299ceb808b4b887fd834408f9a0de8a0a3076a0bb2d5bf993ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h35b83eda66fbf66e0e43bd1ec075d985b69169fab44786604eb3e5ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188df303bbe677892c832018908cff097360eed88b59e3eb903ad4b17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a5ed08730ec5870410a15159b4eb10e8e44746231e7a89a7a16e91af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1426ef40c36c4ad059682406ec0093c1e9389fdee1f5ac7dc82dc61ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141743142d09605fca340ff937fd6c011a3410753b75c4f70152d894d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdcd133f64da5870aa1db977ccd0e6134bfadc9be127c533741a259ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1991fc91b35ed56039327ce37c149f13b1d3f86b1a6b898e0f91e4cf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf1ec266f2de1e7b9d4d231645fdbeaf37749e95e40acb744723fb0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cfc57c8f9f995ccb619baf8237701813e539d755acd336c8f32c760e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee6c66a05808a05647f193b698c05885fe010121513213fa82f07e25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a8da39c1caf96c2d6e76d183514273371854e2ffdd6c29bb7161e189;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h99213ba9e7a6cd41d5760fef6d9d8705ae147fbcadb217de4c41850d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1879775556bb21b0307d8660cbd1621260278dc79e265507e65414f89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2497c9f303fcef702aeb9695c55c4fb5bda9cca4a38913686d603a36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2d906ce0ba6b18a548d89ceae6d237942f0586094aa1f725ab19b1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c88bf4a71f46357675b841521884a2f39824335247a48afbc09f397;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30b944b233c7c5abad6284d1e6e20520d930b66f736605a89c9ce5dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17991b20c0ff0205279ba6ed4b905e7876488ffdd92864ecf1f19b170;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101972c8e21b9396699a0444a517bfe8a194ab8cc3a3a5f827a945d89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he0b5fda9ce3180f81793cab9f98b09bf640ddb69330f725e7f868669;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd89a2bdb231263b3bde6d2fb6bd4df4948f9e067a8db5d11d8103c4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd7adc13f6259d858875f2867eb81f6c5f8115ca4886c6b621464cf74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc67c765da764ef4563ff74096b61bd94c06d99d19548d1439152d70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf220a3ba7683e1dc51bafe2a65eb2cf446c5818118f51acff179df2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ba2de60ffba92e048d463982a272cda8299270946af43a7541964f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h477f63d1db630018aae6a7753b73582c59715df9c7481aca903f4a70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3dd6ed89bf548b4d9f29dfef24f3fdbec9e97e2ae42ae825a74fa0f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha97467e2880fbe708d9deabb015470153d885aa753f7e7208c4f78dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h54c6748c47062e86a5bd3c224d515f4a06281c44ff1451de6a214eab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a92ded7f72d8165ce81b7b6e6ca10d131bdde17593d0fa4403b28722;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a64d2adf08fa39403d3efc5b64a563beb319036795823658c452b126;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he03953ab84bec8815894dcf409e12bf47566400bc354ae192d320574;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19b7438f49c10cfcb5b0d164d893eee5c01ff0a219a8eb01e9040e85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18246e73c386032582595120c0fd236316454d6bb8dd71f233e372965;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e18b6438829fbd0bc9695042954f576bca5c1d73d6e699548e0f7d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4cf04a434b348b9cc3681b706e09940ddcf864b43f9178d05cd88b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19ea2fe305791db8464001eb1707eb2bc466e7052d31770ba8ca7d368;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32b6a29c5341e497c0c54929bc14b25cb6eefbb9de87811c8d30a8c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h144575f97bc8790342ff407fbcd424ed3d321f3537bfd165931081d9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f6ebb0d6d48d0e919c1b7dccc10babff9fa9395feb5a35ce3f204f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c966589c6a440672b108d87cd258563cd754d96c7b520aaee60f466;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1695a82bad552ca512fafa70964775b68b126e9703bbc2d22aae667bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d193f983fe54068ed8aa4dcc0863829ea32dabdef94eb5937c123a3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b310435800240cb2ced9007e0bf986e91bca0c11a96db2ee1c0df199;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hca5337e428f6f31ff0aecc2f75981e287e2de6f03d9c15ddb0d7b7aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3ffbabed7a552e8c0e944cb2aeaa6f2819ab5f0ca4464f0052092e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1174929902c16ed0b0b0f1a769e80da51afcbb249efd280c9bff15bad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc7da8b24deffa2e973d0c0d2bbb490c13c5ed527d087051805502cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d2c58837497e77a30c28c2222724e245b53ae568f3454d1c1255e60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1718a719749c6a0a5a7126dce0ec0090824365e35fcd10f388bbb4d71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h567a641314c5ef3362b5e833f6810a39faf201f98f24e1d08d9aa269;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h68b0df0cbe55f5998d5d4e1a6ba6ee1df13a39541379d6f488eebdee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c8212aa3b9331e20a7bf585962d1f3664db611586648cf8c0ed6742;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62a72dee2739437ed9a57dc96a29f7051343ee00f1efe6ceb7a969fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa86958ee2144b7c72a112b6997bcf89be525d6e546b818adbeb7efd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111761e85fc48d670e2d81793b42ed09ff914a4c0e69c996315ad728d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41d03de6dfd25a3101ca9342f03e00c39edb2acef67bbacfd0b7eb53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11cd39beef967f7726e65288c418c0778578d01e81a38ef39ca34c7fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177580558777c8af2291f614f8617ea40da1ba60f500234353b7c980c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h100208365ee9f28c26bae5c3d4fec8c6ad97d287c4d06ac89bdae6f3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce389346ece2aa219f8fc07a738e6e3ecd8c0bfcbada34f19ad62ffe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h167667b9d2025f4ee399aa3fdc9c057d177d39ed25b3bc28957f14578;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1509695eac7200804f929f97bff1e466acdc4b429f0fa03fd2dbdcada;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153c5fa7590879d936f6a91b8533c5ec848e8cba1d052ad96795fd616;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14fb4c42e0f70ce20cc0a6fb6931a602cbd408ba09acd1b27c56a56ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190476fe9a53db7936521fe19beae66f92dd5921e965371bc5e6336b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49c577c73aee2082d9356885b2e0fd5d86de9af2ff96f72c9ed614b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2076ea067133404dbec2c0812e2111c94ca058ca8b4732d0510db8bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109a36b3fce2928b9827cb227f0496228276cbe136046dc91276c6a6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd97e97dec9b7aa4e8eefd847924280ec372c5955f38e2a1fe716db3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a67604a5e767fa2f8e2bc7b9dcc0a8b0d7ef4a5f115479c44ce3daf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff140e796af25774bad03b24bcb342b8f52c264629c7dbc9ed5b8557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93cfd682152349e3bff22afe7e1f58508d8724a221954bf6421e4ff2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h180f6aa3b264680147328b44d901bed70b0fd3bbab71b6612a16482e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h128e76ab54ffc01bc4dc3e4126ef66bade40f7967a20095ad1656aaed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c4049c60eb90dcfaa86091ff0da64deae003774763eb1d42aaa1f7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b10ffce6b201f1d04e9b66202dc0e2ab0b23e1724b1126b2a339e752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a86d5502308415de337b52eb9320b4ac373f9a98ec900e37b8ecad22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e981ddb84715bf06fea6be6af8f011ad543a977b02d8d0a872ae704;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec8cc519f76be857d207e908f4e3a8bd82d1bc81f7b684c932478a34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15174ca7e4f506c0f1d8e56d3ad625aca6537395f146ad6e56485e6bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36644ebdbee490271b0c4d90d9f0915af9f8051736813cd44018a71d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1802dd35c0a6c1e05918e58b310761c7810fda7739895cb11de500954;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha5f73b58e862832840e33fc180475de1601919cc9f9371c4750c1cc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ec9aef3881cceace01870aad5de92892a73875a348b3c8f496f0bdb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a84ea36ec51fb1a8c3c7ff7b8089b97db5b4c14e2c4d285ca6624a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb38ca477bc33fac274089a724dce00ea0e7fc1d3519199d3aea3407;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b7ad843da8dfa6c73b2f422b395c9d352165285020e1f77d5ce9854;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9bb7ca68339bd90b982f77c1e6b9a1f4d7dcf63ec7b26046fbd1b84a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac7c9d6e022fb4e392de505aab1cac107029d9c4257059fbe8456632;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be253e8befe6efd5368e41ddcf474010b4d5dd1aa2dcdd133bb16857;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf31f023ca282357b599b82c015452173ccd5207dcb41b07b795fa8ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e35ed7a1c3eb25c1c92af7c8a6030491af0188c3a02a967322ecd56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0cd2e11e33db631f606ccbcb0e4876572b6938e46a8dd1b43a19d2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14cdf83a3713f8cc24f0c83d7bf0459f8003578aed07df726d1d2f65c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87bdc8863a75734998605056990c4923b2381ac0393cf75609f3574;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85bfbf9c1d0c4df60b87e77befedc47dbf775eaa2a3f9f3a4fe545f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he2c96c8a618689149deb02681cadbd66d82101b7d9ffc2a65907a69f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h400dc60ffc8d37ae147b1ddb859eb285bff0199bd3c816e96f627226;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb05d1192dae11fe590ea8f10ffdc0b8193046ee1501d06a90d0a059;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85b7f01d7587a1a127b596f45fe4167e773787a15653fba3abe4f6c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he41cd4c734139e33fbcf5e1cee9567260295ac8337c421c9d6734ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4db6571abef621c3ee269acc13dca175f2676ad30d4fa574df333fd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heab3f924b9bcde1ffc32a3e370351f1c262c4750a336d499a7c60b6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82a942c0a69c2012271523a190f5b27d47b1c498bc55affbcce216d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13798b5415ae6fb7a5ec31797e328c4e810e0a827584ee799bb1da771;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11093a8dfd7550b931010e4be409253b3b2c811fb1e13e4aa9864ec71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e462090e6c8f864201bd3166908d3cb9f7794d79792e5c3dbcdef70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e657815d3ce9dc621fba8592437dfb56c929af214dab57f51aadae00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h144757fab03f40519f393e7250e6b6f480885408038d491a4c2256e06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5fd7bc6f3725b85eb0ef8d5b0ff2a4341179e8b95c83bc14a1c550c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c01401f8a5de0f20fe2c6c5bcb07d65b49fc662c3e90bda2d7cc6ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eda1153decebdd658525c0ce5a886bf273f159e46366f5911ce1d54e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1092da82f9f323ec9f21a9dada576b31353999d970f2538b65feac3e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf14e1fc89c183a688ff3bee175def3cdda4ee6a1cbbc5fcfc090956;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1d064be611cf314b093c445eb40007dfcadbb2c04d1e7e421b259a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88d7f40d31a242fd8a9fb9a46aba22ef503a363937e390fa79e810fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a205d43d228766938b4bb9f8577a33c7261951e33a20072b0f7f4da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f24a5aa46d772a3047ba1bc8599d1770917dd43b0a67afaac6a0855;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15852182ae51dd2cc95b852873c00c8d897a9830a379327d1d8ef2280;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h609ab73f89e630a4479685874f3b1384cdb908617358f19ed00cb713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1495e147f5a2a073d184c7d79cbb26fa33b03ce144687ae1dfd9f489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dea1422b2f3f21654c36b1b30c40840b5fd33a5ed8303eb440c45793;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13db5659d90d15376205f067d7242c0a2135643f7d5df56aac88026f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1ac7ccbd520dbbfdd2b2eb7614f661e2bb2ab567c510409ce566440;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a5d20d5abf3e3f2a769f91ad418917e03aa7b9b56cd3a6ba2515f74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d1845fb46cd80685f841519235347dda6485bfc237aa2dc7fcf65075;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7887a95036dfcca5709d9448740324709cfca4a89e3768e71f4478d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78a53571827a33d7d6a55d904df65d8f0046d0b9aea5c46d37dc16e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75e501555f9f049ae5a5905f7bb5123a6db2e6ce24594ba3b4f045e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1233519d1379d81da405ee903c83509973272533d80f0f31602d2758f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd26b48c029b58b62ad1da4916381f8485acbf3e3faaf0680684f42c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126ba8ce8d5859fc2fc7690a03c2e0405b48f8b631826219715cb107;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd4ff3f12cd026d4bb71418ac00f5b342062b78cc58a1a104fde631e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha506251ce07dfc93a4974f070f90980780e0230a49e5e91c80fe1879;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3251abb09d0d52a9d6bd13f8bce3a83b71c8d75177efcb6eb77cb19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f281c2899d00f5c3a70597dfd6a2d4fa0c9663097467cfe7df5e20a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c675d7d6a4eae3b3ff8b3c74f6c8a5d1c7420d2776c0f1beff080ea8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4e7c2892c0adc06f70c5153b54314a3a3abd26efc4e21d7824dc5ed4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb095a79b693d89881af2ca8dd2628a7394f95ada0cabc7cbab29c81e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbbb24489942d83606b3da244242c7f1c1ac54699e5b66e1cf91420de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1652ea2ea766fd897cf263b427302507c472a915f76609e409b28b0fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3e478b43394211406c16102ca89cec5ca14dffa9ed86e90c658ad5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0893e604fe7aa12999892376a2ddad027717a709d35ab912ffc8bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac887f354b259c964586974bb60dcb2a0f9374ed5cfb30fde316641;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81b5a14ce80a964c44e81180885bc62036138f0b8fb08d4548ea05da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h844a65aaf5469abcc3e70a708f44ccb44373622bb8a491b1ef883077;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h140a14fac4d0a44f797c916f7958584b6e065ad1aae3bd33fe69a01d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf029d1a909042229cad7edfd16cf5da4b8eb5589099ea8bc709ac0ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9cea12a69863f6daf3b51c7d5b5c7826ea49c377e103e3ceea521ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9620f311a09f22e5b445055af3baf004e1dad74cd823dc9e55bdc45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16bdc0faf1ed7417c877c8ddb6f59a53c37a0c59b6078b25cbbdee06a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b9474c5d354e99c5e962c90f5c511d9f20424ad678b4196f5ccb49c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11dc2334337c6b8f76d9d8f44898b8505d3f8a52dfa0b817ccae5529b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2b851bc37b8b8befa43a0b2f934434e772dfcfde35383e980f8103c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101b29449db2b92481a0c23b3121df091422e386da35055f8c28b85a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb9840bbdb0b7f3b45d75e12aed6ce67f6ac9b79df1e84eaab9b384;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda49a57787c9b30bc16af0876b8467f98f7fe58920a3864219235ae1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126761b1b2b86c5583a78839d09632c3cf5e2782673146762cadef3ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3c5cc808a5b924cea41637a695fa0f6a381f8a1cd01a09b4be9c73d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13082751c13a3ee8c935f8efbe04e6c44a6496ea480272085d356cca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0e85946dc2867560a0e386884c93c90b1a967e29b55ffbfe0488195;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a6dd9aa17585185f3856e8275ef41af00516b457eae0e4f169a036a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h183bbc3f597f9698e3f4f601a14e8aebc6872f995860b8748317562ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9da8f94461a1dbade6767785117436170977fdd1ef1b2fd959741d02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdfda2952745013f22ab7157de348bd315c861849b2ff59762d444fcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d3150bad53bafc8932fa6a9dc5564a167ce355354b546c985d260fc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81f06371c6298a10a143d5a9d9d1a2d8c0d29d77540b688995e6a2dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8252fb42a4bb71e1bab3be02755bdd76beec200b2c295fbecc823992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b680d6d4363b88b8c6aef7b178b1e6523718e6d1634bda1947fc4ef8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba3f7b754a57967e480ea9e0c4b421d442030db642d932d40940ce05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb69ec75d49cb48515a18bc9afea9b743c1fffebf2211410a4bd02daf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1993d2588f3d54a0178085eab8d9f6ebcc03e0e34eff6751e48d877c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0a49aa5d9340c090f1c03aa326999eb305145aaae5138ecc1a79a78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34bda997d07c30d31f85e81fc5bb0b3ce976e827cb9ef90bdd5abbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed0ec92397e52085c2fa7e48a4ab0d77cdefe62bbe3a6b0a98e530c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9aa9e264310460278d9de2874393e78112ad98f99785a38fc55319c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5f8d72a7e9dfc88ab367a50067a6fc8215a3b26ecd5b1e351c08a72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h121a09d40fb80f249f043265def39773f1d29e27bd9807b811cd16653;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heec438f087e763ccd66cea1b1b4b968af7e35986aac34e92cd6233cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f89031708a5dd587dbe02567279fdce8ae295a0fe76360ecaff8f9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f6687a8077517d3218ce25bb248f4d7d77ed3270dcdd6220f96ad33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a8cfa10e03ec047e2086579cfa41f0598d53cae0e2808a9ef6c28d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f5eadd03d50da6b7806c159f1f4c2b881990660dfe3037a7ec2bf3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8cdda4440b08bd6c2502114e383f185232c3f36b6b2012a6ea666921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf056ab86beab04a5520dc596b8bfe3abadc997967fb1887e1b158e90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a6d9e0b421ce9c1a8f495ff03fd9c7fa65a02273615a1b3fdd80585;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9401ebc2d788d3f4d97ff196bf0beafdb50b56d3658be53b4ea3fb93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h978f26d27184193fad66dc6f0f29d95cc9729af4807894ba6af2902d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb5376213ce86a7a2a9acfe92475ce700a0f14f22d5adc2a0e003dee1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c77c5fc565106935f400d2c8ba0d4a3f7258d426a4442b073f13cd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134e4adda82a04cba08e4dc6cccbfa63f7031c1721808425b1748f7d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11457bc24d37eafe040b6054ec5cf89f05ecaef0cc86ad9f12f977124;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13003593a8354bf17c69ebff575d492783cf87e3949b3fccf9273ce0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17db886c107a68c814ac93223a300c3efc2593facc048b51ecdda15fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e00624734732d4f37bffaf1f015c64ded3d2c4c9a25e3692c65134b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9568a60c575462eb0313b56e7f13f157782f325f1b5eeb7a6f770543;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd75a387a03167f59fe1e12212e527f7e3b2d63a7b64140814aa7a6d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c4cf9792dc8d62ffa7f64b64fb40e9b69ce346d86761eaa36f2ca63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h741a5bff4c345acd62fa3758c86c3f3b28e19cbb2b3e7ce86c727288;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a5b59d79a1c02d14fb918ba63cbd415e068bb37bcc9fa37e0862c96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h705441aeda52c56b6a605781e75c33f17932c2e17cbd336ed65c971;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1185492cd57fa6352db2c91bbf8ed5e9f957e952ebd0f910d45ee860;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ba79ee177995ce855043aec274df44688e8c473a57eeab4cc44482a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2b68a11708430a4e16bb9a3b6e32166c4318c8aaa0fa292dbefff9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1236d58de5511275364cbc02a82db0b862dba06abebc14738c815075f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c8f55a14c4c4a53d803688ce4bb33045b70eb107d765febd87829a30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd767e33342e2ff331dbd5f404a6f88e03695f21b30643ee0ed59ce33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd656624986c9ea1888873f1c38aad87b486191cb94e378bb2a5c0c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h650148a4158edeb2c2dda336464e28e81ac1baf0ae69359d2b67613d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdbfa690cbdd4445fba523b4f4e1d8ae724fa5a920f02ec9abf52c1a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51451861f6a48edc76d86a5c48555d52fdb3a35c36462ce233d54876;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h523cb110152579027457a1190ceb54cfec542fb79c3eab2470af06a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe7e3f3ea9c5b2ee8bb9c0e4fd0cecbf6589aa74b383bffd87be723d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19aa07e8562aa3580930a14091ea0100f5e9d413b6b03013e08a5214d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15fbe38591fa99271a572bc3a71ed84c74f0b26362909070a5b5e5a9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb22e75ef7a352d017b38b182dd72b2f7838ad4abd49452136c894333;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176cdfd8d57b89e6fe366c7b3db98c3a7f70dfa032792884e41b2593a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5472d1f5d50eae7367b0a4c9caefb702871f5a4f9103e1c23a50827;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1303fcae10928536f68b34800043522852f0d7738d9b22248d046453e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1732cf61157f7b63ae35acc8608ca1b0110c8c561346429b68f5cae43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f967f3790572d1eb2d1153d8d8c3ef3ca0226d2262ab5545289b931a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83a0ebe88a51eb4eaac18754187eb9ee0d8fb837ccd3d62403571c0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h628010a516886a35369fea0b3237b158048bdbccb043d7471b07f24b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16e7c739b08742e7ea27f7e1602247f675b234c2fc36c6bb6d90df49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a8c958782dbe86fb5538a3e8882eeb001ca61cc43e8ece5d6004516;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b86b338fc739c1e836cfe5b64470118a42fb10a72b8cc984f0875d31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b311c24e95ee34e889e88c8826884d7816cdfba97122d4683c0fed8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec7023ca3e957ce73af081d109e57fdb4188d7afbcf2882177e86671;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca741da34b2cdc296db86302d41b77061adf2f5ae9dcfb596fb13c9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h57c7a590ab2a535780e9c3ae4012c948b075bc91c6f56884c43fa742;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ee2f6507e7426d2a00728279c8a6402cfbab738f7010573166142cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h186aba7f1b9c16a1a8f3d60c49397b6986b250a5c95fb902d53759a3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h520a7e4c28cc93edbc7db63bee9608f825d9c61cb58dc8cbc3a6cae9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hce84f0d40c807080ffa9da221199bc1751689973f393bfe708cdf3c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61c89af61b02103063a0c62bd1a1cdbbd530f6c9d2fc21aaf2810d24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1332c64ad0784fb0bda594b320fc89eaf07e84dccfa384ddad91a998a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f627f6a8604c17c3784a3215b639ed7a0838bb6d06e1554f1e0c3de8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec6b58d2ef05eb8d40d23d68a6b6cdc895cda8487a1970cac310be36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he33e53e428958d052771a3022521f7f462d001c6d62729674d592f04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h959e65d3d62aa0fe74459b033f4cd7aed1b42e2daeffb7c99406e003;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1beab3f014bcc2983b4d71c2f81c747fb32bf35cd5f238fb6be510428;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123fbde50843bb23f901a877e2e64b0e71b53ede83684547483224281;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h608d60b44bb408febac8dda1c677300da76328e2bb8e46cac3cab29d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17756c1fbbf5a577a590f436d98da7540230679698e47570c6ea0d12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d5b75e00cd864042e98d1c7367048991e9bb361f040a9007438faf0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h628eae15f06fc08a2e67a416163d2ad04a4f09aa3ad9c801ec0ad20f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6458a86af8e313f92df7f18537c703505ed21db8d0285096143ce19e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8bb03240cd5ee5f37b3f965ad762892dc8698c6a1653a84253adb2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1781ddf3d40d79aad1c288c509cc7875d6a4423ba89989e714d09dc50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha430bd04e4c34793066fbed604c6a174253d0987f8ffa9fa63a666d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3698ddd11725c99c5e6faa1e928c89102c2bb7bdc6e1e2d69cab807;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda9d9cdca5458ace9cc09bbb98f1c067cfd69375b4f373b55eb8933d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b775dc4cfaa77e31e3fc4daf1e280c5610177c4f1c1046e1c1c2495;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10127d6ee0db76af285ee446a1c26432475a0da0a7aa1cbb5a6ea49e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137ea89875ff51ad84eac07ac878eb4d6880ab36aa0047d08a1606cde;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14dfb69cbdf5b01b3e321a8925d8684ad9055569aa7ddd73f2224b15b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h544ba3e7df002516260af4b33b01d308f6f629be4e6d91e92236c62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba6cf523fc68e3476202c54d400f15e5890fd76e398ff88cece2cea9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8866b2afdaf66b612391d025e5543c6a177d1d027e0ef831ea50779;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a477cfa6744d8aa82363041d9fae61b7c72c506d07ea593befd2c2ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha34e28ad6f40ebd1bd0efda26b421e5485d6fe80cadb1ff542d9ecb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81dea9063699932f80c2ae44a493c4ce9bff6ee5acbe6bd0239a2b67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61af0d8c96fd633f9153094f8b54a588d4fa8d7bfc6cb51e4ac0d88e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17bdd93dac0c13763e29a99486b77d7c274429771fbe9e6e1c4b9c1cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181d7258a606a08bd6d255714dfdfe91b7568e36ed7a9c75cfd1fb300;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3bf651f3aa60d35ecd3613a3ea4dcab36f58b4f0efae7bfa873754d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dbf9b29c31cf229032f9ea57f1cbe51cbadebce6ddbb26d6800c853;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12c019f29244fe663080e8a44b4988336caf49553def832aa89b3b229;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff341e802d70dc3d460a9e21a9344dff2c76c0a623020aaf8de1e919;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17926888a505f3cd6b8a7ddd1bd849466c8d5695154c551a2d33f2ca2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h31d299d9a33c77e28faab3b238cf6cb8e4f7d53fa0885e248cc94241;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2bbcfed77c7b9f022c72eaffaf681714e02c116c82d709bb2ae19dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113e53bc422bde3677dd865faec5112d1e58f0682fab102339eefd310;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83446c0a65b37179cddd7474340f7ffe09ad1d27fdadfa50cb8ed4db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138c4d82a328e591afd0a962538d324aeb138371c408bf326a2fc4fbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86435e205e78d8c48963f3289e10892284170040d21673e07a416696;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139e838dbcaffa5e146987457bad543058f79417a245ba7dc8b836c35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb6e6a61ad731e6ac79021bf8fd0ef44938c52a86ed79c608695d6ab1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0f2705592628cb1aee51d7456a84ce1b2b3348e9eaf603c8ee5a204;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56d20c7315e01e347ad1da7bb203f2d4cdcf7f4997e3b5d7fbe1138f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a9d21e60cd40b231f5d5d7d3437ef2b6c3cc93efdd23cd7f4b708cda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2148f0ceaf8dd285c9d323ee2b84cf28242c74b1d76332595a421009;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95204da87015e58f91a30d3f3214282aa471ae4f0335347cec8f1fc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd7d8abcb5af3ae433390436c770478a23ba864974cb763bc99fe24c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ddb3fcb660f9178c04a1951338ff1f6e9c967c77f86ea6c3983a8613;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f7bcd84ef100e63f3fa918ed1f3654c23b3aff75d9c233bc1675d24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ba2a5344ded73499ad3d91497163d77287bdc4fb608b2af336864fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d24c6f960ea01264d83e24636c8242c77f1d03af800af5d9c04448;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6398e36cbfba71f8de6ca2d819dc4ffb04182f8ee7cc86d4f141faf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3314d4a60c1812db63039c00bab24fb91a9a8dbc3315fe11ff792026;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h44e750158c3a808c8606519a2a0d2472dce293ecbb8f5a7526cd2455;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a60425f151e233c6e17a59aa410df3fd718bcca8344f557463b091f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h73012e48ad3687b7e6872862b68e1c1e9ecfc580b6dcc78e69048c58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70a051c791c4eda03ec8b2efd314eb6cfb08a32d335de9bb6f2c87c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f40a83584f3a5fa931506724b3c2408b850f9eb0b54a9b690b343787;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1075a97edb45a2c1b17c73d27a24d35d6ea77972abe2a9f12cd7f738c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a1d291696c27bdcfd9187bcf64401218aa49fe90c842a20e3ffbe78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f9b4ac781401a88723c06e15f0958fe1b18dfc55c8eab2bb2683a0a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ebf7d428ece656cafcf9138864838f9e1ee44426e213ad7e3d1d243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a220e4b380c1a5c490ae06c8db9b9b43dc318f301018719dd8f13c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1715ffafdb8b30943ba636234cf6142576f6eac48a833380d24932f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a4d96676b4b83b488bb78faf6a18dd198e3e1434def2e417651691e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haf00b2c3dd5791ff4ced96e0f5ddfc8dee6df086cf9507c6e92467bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbddc5d9718a28d7f6a4bc88dc129b45b653d775ca796a432875bdf8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6104caed9db07e9420fabaeeec9e685245ca1bae4e5d721e8d3166ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdaf168a25778b97b8b77fdb6e559f506dda293cbc3519abb6d59953b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2b63b49b145bf98cb1eede92839520baf6ca75cb9fc91e8f7565ac6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15547765bbd9496f75c59790f6d4cddff8186a805e61195f1529f411c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e4e7e2ea92fd85deb589b095ba29cad412939f62065e4896195a0c8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4fbe1d99bcff640fd1c897c8235dc8f2e50d0b24c4d0434bff4576a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd55f79ff82deba60bad88253fbaf7163066e9ea6221811da61bf4ca4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127d6f58059bbdd1014b80ef32a584b79ea9636828040a3b462b8fbc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e4991b50e2de2dd7f426b0c5c8f88f964fbd749fd1c2d4f6a85c85c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b43d4627f79e0b8d73e74e58e93779524cf4d81a615c4c08a9e5edc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc2afab7c09f3370439daa93b3ff3ebd31aa20475e0f3de15d7ee3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55799b05c9540732efd0cc8696f024e707e2dc68085204d359fde119;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136cb16476c42716d106d89df227bd5c3ec89ce435b6bfa8171029510;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e25a9c9e41b90b414f91ee19afb13464bb8d465ce9cabd98c7bd1cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15bf10bbe3512a575ecfcec87dc068aad02ef832c97dc0998deff865d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ad570c23d76a3b12ef2b34685b5026f156b55b8bf088415849344df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d26692cf3757efaba89ba2708a95e0be904785c4684a9e40772eca4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be0145ee3c0751c9a9e030f75773df06c4608748d2881f9c66e91f3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1151cc3af6914cb48d0b54edaa88ea876e83cbc82059663b6be356de8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38721a9362f99564f6ef5ed251fce055a1b0a2215cfc2b033da0b4ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc25eb1816a8559776b3b55ee08dc790243a772ef3aa96d3efca6c4ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2080e8f222dec1836fd4ca4e0dee0728576fbee1cfb2afa1609fd80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90124a49038166bc312888dfc0e20eda5c65047040d0497bb712ea44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbad2219196280d65cfbe2ac8e4430d57bcb7aea00ea05b499bc479ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ddf9b18c20ab9e3f57b66370e7bd3d140462977c8fe4f20da19c390;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d82e8a782cae870ada73d860ff67062eb10d9265dc17ff2fb959dec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d86f801834b5c143861dcfd8bf3a0acce7e1ab717640dbbc0695e7cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1401936df9c50705bbd706fbdeaea82dea51985a411f94d659771d76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14963d438d4e4ee29dda2f8ec1be40c999bcb8390a425d6f15b62bbf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he9762a3dccf70e260a1b82e3836b34a1f544166182d0f885d892d34b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147865ffa7157764772ab81bb68c51eb32b7cfbc8097be36e61e923f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12523b0f74aaa1509abbd89c7dcfafd2a559f69755b5f5faa48f7713c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hccfd9631f11c599784a09e0f39f5b99e7c480b097ead83bc5d3ac7e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc610da29f2ab28382e5e038a0925307d37191ca8c2f2376f7b302fac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5abeb382df0bd53894bbd394a906769bdd5ff9bcacb67061b641788;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c769bfb13c0165eac236db5756991d5d5e89a83f76b14c4408442f2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37837eb9db0d800650d4ea505a28b6e77ce362aff97d4de370f53f85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14645b93e20f413dabd590337846b6c43879f76866efd11dfab8f7704;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11888817f07dda643af94a243e0a3d23832dab07f5f49f4051ce03ab3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f02420f582cd5822ed8ed8e2b032071c415aa6e64ee8c729e3f1ee4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha860243524f23eb143d8ab4cd676cc90a2146194b28e11dd47711b32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32ec438de3fe8bdf198560123cf2e7be874108327bc0a96180d0b845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac261448e05a5b6330e63876081b28fa2492c1f0ed2c731656c2f3a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18672d9c6c6428cdeaf0fe50061845bbb5388522b39a1c4fd80ce6219;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a831197f2f8a9c7af08413da64c10fd6c23de03448cb2e6753f1ef23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf7ed0ec6ee0a7962ad8dde023463c0f112f48bb3289d11eafa45e9c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7d780972f4c7298cb06c14a10f9cd1a2ee4019ac86d7390313e80bfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c0584f58f829682172c099e1fbbbf41b541f5077f7fd8e221fbb8bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h130a004a13bc0bb00b5c0edb5746722c75f2079bee21897b31bfb5e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heea650eaacf348d9c786ca8efdb0d7d6b7425b72db7169b0197001d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d1b735e2841e472a002f9c02af4e26ed7bc1cd6ad6e3e0b9754ab32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h199b14307b5a1486793cbc3b68257a3573ed8ce4d0f65849752485f20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf8e889f3641d7179ed5d88e0f8062144886e1ce663d79d0abc46ba36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he294dcabebf37164ee91e0c8877bcf8d1e71543b45bd97884c5b5e2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8c75e740a60f68a433bcd0e845712ec21bbe07522716db74f21adf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff009d8443e94b54b4e4d33d13a74096f7cd37b5e289160db0afada0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150ccefa4937a21e6b350668be77bd274f5e76badc2fc8e7894afa727;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a707f987c037b77711eea22ea66780e60df0cd534cbde0e4fb9e3f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e68dae629e526b2bd6bb413afcf0a8d2ee0928bb96011fc92a2a158;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fbe1ce32864ac13bd890c2d304623780481c5f7599ba3697c2d9f51f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c2327f2c7d2e465c6792c310f0eabb622dc2aad6038bbc6ee35974a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e30504763b132185f1bb31f09bf2640c73d4e06947d5317f865342d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a50dfea8f6473f3f9e361502e353e0e169815b37c7953e3d50f6f6e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75b8bacfaa40c4ef87c6d7d1356c8f40334c440f00d9fac3a0450fc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cab270e9c1f0705919c6d54d8e8b7553bc891b6b02ab97ce9865d62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12be0b02ff1b75301e9c7b5664b101f2a145eb3add8225d55c54e6f55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7eca66633509d5767ae671bddbd3f7fa5b42bb054ecfaaf25364c89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103ae8de66d76e01ec461fa8d73d06e8271a92e4aadabbc0864f85e7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12838e3e3ad47a996e79c85f8c6502a1edacea872d61cae7b50f756dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b94bdab9423f5f1a27eb1dd37ef559bedbe9f3cce06f085f4ac7746;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a228de2c4663ae93d3c2f1b7ec804d2b1b84dc1aeb664975019d53e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a64853c43a23ed3e95c4308bc7b70c9e40a68e092670ef986b2e34e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ac4850da670b2d143a43945e0722b5595502a48524f69cccf4efb8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a9a097a9c5c31c43b41a6bef830c3eb5f974178f23f6901c724d73a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a989d215b799756c046c874e6ab20e05e5af0bc72e12c513bd5e30f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b616d5e9e7eee14ae64d76e3cb38455bf5a54d478b3c40ee25776f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f579469e01874b14f25ddc9213233f8d218962d0477f4df6b5912cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdd11e82a01e68d0c3397719c53b1edec868a5c0ea91599e6c49f386;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17442e61d3ba6e4b151d9c95a35869ac6b0eadb8ec92360c52eba3336;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a44a3b42ed6642935b8c2b8f402a1de79d866b035dfd1d2c462b32b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd672a9d8fd2d0ad2a93db6a9dcb1c21b061584bdf4cca8a9ae481a37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9b8f27c61e5d61a2bdfa3e31af22441063c3581d209de28662cd819;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1480212ba9f9fecb9c726dbb59d58620b186fd578277c557fc53442;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc24d8fbeb1235ddcf0dac722e027aca102001476339c93f9bf6a3a49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1885ba9a07b6f48609e42a7540c027f0af8b0b0f83bb4dcb912cb13a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd27887fedff106a21f349c511c1cce2eb04d79e4988010d7908cd28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148e4813176c54efb2ac8e0aabb02b891f65d27dec0c1255b4fa5ca60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h46595df4fea78ca679384ce470ed955f3be67e62f2a88ae1522dfcb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e1ecd9c420710ca9e8d28483a14515fb007309842b11aa1dce32d5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c59b941e4a014b8b31ce45e289562619fe786eea1b34a77c05c7d26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef553dfa76f6ef7b32409ce44742109fa3273a5c0875420d19984d6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c26aa0fb1f3503a5bb99fda4a255bc071a020b38fdd7be3ad6f2a3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9de1b2b367e84b24a044e0cd4f8dff86025086ee4fbcdb1737a27944;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb34186b15d956cea4f3fd274571272b186afdc76f9bbe9d7e9959f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a9c04dd4ef1e151119a97a21be5cd989a55a41176e6234f970f4130;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1b0bb5774c3cc208e2b1d1d978f0a3f0088aa1483f121862ecf4444;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5d72b600b14dfbd41bc4ae1b7f513d3ebd20bd47dda22e0b4e55ad0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48c76af771f2f16c337ce3ea3883e3edc27b4b52c9da0270f97ac748;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fc842b22f2ed6b7bf54a1fec195689eb62e05ed1177153d2ce2e0cf5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf68fc41fdc1dc512e8bd679fb5551e03c397fea1e318692c2976ec5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h77a139a8452139caf0d26af5caecd7da2637f86ec3a5e9864484cf9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc77b851e8b0e63fd3b606ae957f5777628313a8818fa5532feeae8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc93cf662dbfa9e041d04a50814ea343e503ee8cb46b9fff6639b073;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7b2560b52c28d979ce1979ba0a8323882573b59964861896425f600;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he61ae02b1c3b59fb81337b3d4696049c3f588480c296bb16672d5457;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2ab6c63356c5f0f71fcbcc0bdd0880833760f08554bd75aa78d3b1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h71b02d5685571904c88838c1b02c449c735daaf4605bd7ac2d426d3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6466ad036406467c2ab7dfa3ff20b972bfc56f35072f41681cfc57a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ece5ba9bf8319b4e1828e0d40220c4f1e0a67f84dde884cc2deccbf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c218c42a71fd948f5dd5a91867640b0f614b1e77af79628418e8c429;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66ca0ee4b5e5e237f6b1372744e527f003569f91c6238ed490669ac4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdf96e5921ba2b9b7a79d984628321385e350f00d55211825e90d7c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1547f541a030e47d218cc74a12e30429281da59cedf4be91d2d309b64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf82fced134cac0a60f72ea5cc560103edafb07d007121bb97bd23f6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8a80de91e735bee020a3c845936132445cc8635cd4c13c97cbed5c0;
        #1
        $finish();
    end
endmodule
