module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [8:0] src10;
    reg [7:0] src11;
    reg [6:0] src12;
    reg [5:0] src13;
    reg [4:0] src14;
    reg [3:0] src15;
    reg [2:0] src16;
    reg [1:0] src17;
    reg [0:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3])<<15) + ((src16[0] + src16[1] + src16[2])<<16) + ((src17[0] + src17[1])<<17) + ((src18[0])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h330181be40cf4dab6bb46b216;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ad0229493b9e5e0b32bce8ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8573b7f0803da0766feec695;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb43067c93d0ed104752425a03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48eae6dff68de329571c8f004;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99af47eb6b779509574aa8de6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9cd3198995f3d0768429c0a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haecd5ef1b9c92de73d4c669dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cc07656c7883531f8852a620;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a3d4b5105120d4591adc0747;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d4de9c07598bbbbc3755a2c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h299d10301b3f6ef69c00d843;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81cbbaa3d03ebdcd335b4b43b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd852e2e445c9699a3352e4ca1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16064281ae1a81ad42768bada;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6ffe33033ed4698e2c8a46ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha547a57d7765e39e6373b53e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a5e88d13e77c85a2f420fb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h461d851a5667d4b84d88d327d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfce2a77076bd15250e4739ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cedba260871d55548465cc1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14f37a6878d216fbd1c6f26fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h809af28d0256ecc947ea3897d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he86890b5463dbe4154d9ff078;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ff48fb42091cc23594d75095;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5131884ce48ec39018b7ec131;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc82c063a56fee4c65ea8dc3f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70d883d974b89f20b1e5a917;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b9378ceb979a15f8355b373e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7c49e5b6d7c82868e6c1bf64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h709d3a3f97f41ea45d23ab893;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6d9460e8353dad75aa4a6731;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fecd9499a7d81f0c77b050ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b11d2375c6e5fe72b8a83c6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fff0d157bff79a39627f781;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c9034082dd09a5c90788ff8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2292443b5d2c36ce0287ce7e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2142075eaeb89917a9aaf576;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc45dec9e34cc3249f1fb3dff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h378a5146a9143506834f791f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5757d333333adc5297182ba6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc56cf5199749d8aedf0706061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h613b418895e40800837410365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eec3b6b5facd3b70dd32d31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3c86907ccd2645f67a4f970f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e470e4e3cfbf66f8c22ec7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71d151a32fb5b725b1340ddca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2af4ff43d5f2d96c4c5ccd71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2274761fe8efe2a08e48c437f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bba61063f114159a2b5981eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae4a858228bc43065ef3a913e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca4887b6024bf0d15664e61b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5632c51d54d96a3aaff9f87ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fd8e5c4e08b472eca850881e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c9c6b4de0ca3fcce3c81a81d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7255d266400c923be75f65953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb155fc886f8d5351caebd1493;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbef939c159f07a89be4d7123e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h256c15ae63831e00b19eaf7e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1825971395a5e17ac3c642988;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h723f047a2525c109d65b00d19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7069538e4644d2bc87baee3f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7b65414f23c45699f4adffb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8525c5661c5fdcffc8f889eff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4151ed5bab41d4069a26a32a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h560bef6e1c99031964018dab8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5a8f52db6b35f105d663c51a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h898a60e7af16dc93eb8f5386d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf9c76b1a7c379f342c0ea58a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd84ec8a508487aaa4fae85edf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5173488e2492538ababd5165;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfccdbd8a117839b0480f0ce99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h145ac2e39938b9a3588b3d313;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4353616aa2bb1b2593cd2bc5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h594a3253d933a2287fe885c90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31680719383c339f31103f501;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccb30bba1b4148f10ecec6f27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d6ca97429628ef0d98e5cbd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c257645ee2cfdd96f6a7e4dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8638dd8407e8842f5db4a432f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59b4c947c2b3ba8d991c79ea2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd51cd4d2a6ed1a35b147dd1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e2d0d52d9427aec7a5d63663;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd9c9946d50834f82970e891e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a13031fb443355a3c6809fd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5ad4dab7477f69ac94c0d0fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4813c94f301031cb5dbb05fe1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15a8c0adc01f2ad39b6c511e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he569e0d1ddc84e472d0b2cc01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fe033f03ac63b3605e253bae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3746470085d078976d0b968a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6a36e9273f2141e44cfbc8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h154a00b848c8e8ebb4d700dba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had1350921adca3da586b486b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66be8619ad9aedf4b5f38f8c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68a33e1937f613c4c3c375a71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3761bace67d0ecf93e174ede8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3627c49c55516675fdf5d9b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h382ede3f8e4b8b01e94821013;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a7574df933b51cc688f461ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ddad9b08bc6cadb0593e7ff1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had3400a965d07f8ff87d96fd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7d1a1d124a3299e40af2290e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bc7372e800af622f3afe573b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc9238b5f535b4423d6aaf947;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48b3692867f8266b162cfe019;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha280419bcd71c9e0679743ec1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d702e02b27264c6f21fd394;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7fb510e5a85605327cfa3523;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4b6ae1ce51f4a7f7a9294cf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7422bb40260dc68bbc2b79c9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd85419a219df8a3b0166145aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cae833924de0027a5328faf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79e17522105d72fe357cb9d91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7c97d99924bd064e6fd9c7fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdec072728a4f7daa6fcb2dd9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cd20f74fdcb695e346db8f15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc1c9bfac45807010b007efb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heef5e3db8ee73c48ba7f610e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h381f423566272379815622071;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88f0a23527437add35d9be295;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a812560e18bc7f702b57c419;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb33c7ee794df391871df07aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d0b60ada6d8a7f3558f75f31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec0fa15482eceb4dc8095d74b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he39a868ecb69d957769ec916a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a40640769c57dff631ced743;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1c1557e3bb5aca2b5df4dccd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7af1e44c170582be04f4c9b7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dfd0318130c3f958149b93ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf31badde0add4339ece808a4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d2f0edefbb1e5387feed6e5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fcb6a754751a1dd76ad83d1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h687533d9e05f27da2820899e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77853b5374f17148b192fbed7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77bb9b9d067633ebd6234fa15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43d527d686909c85545def511;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe31216a221ecc7f2e1c6049b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd62671b6ffcae3bf9993bb4b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3816e325ddb14e2fbf50ccee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha38a8398f538ea1d084aac361;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f607c502ff28aa9f73581dd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he513381dbfd6982a488d5e77f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7f3fe1333eb48d4d3e95055b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30d3fe2ac4f44bce65e17f507;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h481a8b4e5c7159400cc5d3961;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda7f3d1f60299f80afc68de0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha033b9adcf35643381badd82d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bd2cd5fd67da2a5c4e166e0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha567e7756aeb98b39c91749f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e77e46768ffb357bca076c7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52c8941c9c710c3812d84ffb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef56d80a16f621547a329157c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h890a8cc0f18f00cf67bcd7fda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22cc7325357cf785f4e28f621;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eb91c8c7850f723c44f1dae5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0668d6f5cb987fe71ef6d16a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf620db8ee4696c98e55dc4585;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7302edcf31aaa3cc410a342ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8dba38b63494c3a8faff68d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79c0ca46786a9d5e26a20ffd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77522a4b99065ef950a163764;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19d724a71dea95372cfdb9ca6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4783b9150b284265d7a81ef57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1e87e1c4e541e64e123cac27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfa0139d544f50fb29cb14e9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69ff78fc578e7ec05b4a1f82d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2755e7e9e8cb796ec01fcecf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fe3c9b872fbe82b554886bb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf84f892c0613a27211c18a9ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac31ee9556e044971ed2bcb52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24a4d906680076e0890ee68f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb14684d9091a248829f198f55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h106cda6fe92be826bbc6b47f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58ffb093751aa82b6dc35d7c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7975de8c8fbffdd03ac7839a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a78eb2cf919b346b9e5d39ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc809262194afd3caca1ce1bc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h869c2b3458b24cc5592f6dfea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67a6a05461fdb5dd9b2d541c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15899f40b9778ba24f6bd39db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda040247dbed49f8707ee87c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18f7f8dd8d175c31ac95f88fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fb7c63eb77271beacfe764f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc3fd59c7958c53d34e332f14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ee31b5bfc96991848e351d6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h271931efce3fd6e76064f2b0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4543265580e8d7c8ddcf5e695;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8896eb7d4443194f3f02aafc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h847aad1bd2addc86b32e3f5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e3829d67572326395f39718b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbf7c96da35ff19d9fb525c1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72b1fedb868634964e070c93e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80af73b72f06f2d526ab6944f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bf20a8a1a2cc70964968be1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc6752a2806e1473336ae5f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha61356a0a10e2cf90f2ea821b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa90ef287f191b800610e1f0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d77fe8f9a7e1584a130694;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h337a278b28e569d77ecfa4037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h941fb66aa68e65b7ca5433ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9df36eccb033cb79316849e78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha361b6f5744e3c7c40c59e2d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d6c08db3b84ea6ff2f2edbc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f95f008d54155616d73418ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h302eb3fe0bdd369bfb9ac2e9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9982f6bb6e1e1a6d40cf12add;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cf67a9fdcbda513c6e0f6eb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58946270f3db59899944c5c28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h108d0e07fd241f39917d55ce8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb06825d46f448fd22ec33f734;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33fc746193c653c342f835fab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0a945f27c1b461a52c3d3b66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6218e59b665a1f28a6ddd546d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8808823d0c046432cf235b13a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b21a8bf058bc66514f911869;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2674a8fac8bfd3a10f6908a76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ab26918e0414a33e75e00aa9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48e5352d11cd5308ed8b54c0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b588c3700c8288a879965d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbed16d5af4483705b887670c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c823ff61ba06206b96f536a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfd1840b8b1af73e3c3fb5343;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93706aca5ed303e9fed21afab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44e27f4178b0f897a6509078;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3be398a8012d506dbbb0092ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h163fabbdd68296c3a84304c3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bae30d8657effbab029a7f02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ec290713eb9afb9e366011d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4268e3e849a4e5635162595b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65d923883be8069161c15f281;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf323cdb6c7b58296c91efb2fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4b13ca2a5827c07020af9b3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87ba32bcf79ce532066540468;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h786a5a8124fac0453e18b0645;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10993a92e2eeebcc1404b3b48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5169cc9d693fcf0586e50f35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae08a6548500e2c7e0063e441;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45c6a9ca4f7f6a2f0da7ca934;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7befb58ffc230afe3319f4ccc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3219bad311d2d64fb3d5853ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h250ccf793ea7904fd49c31b6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb167be300dfb8cf1486da48f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddfb948ca45d92602dd2297c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f2b52ee88f390d77870081be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0fa49f376bf016a90e7ec4bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d1ef64a43e9a4e3fe94136af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecafbb4d22552f305bc130a9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0c61c8d077ea423412130b5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce7f46a5e501c20b3f4e66a64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62c5322b2ef52324a77ac1109;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6960ebd441e0cb2f5d72d6b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bbe33eeb5a4e06781d132d20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d3ded552026e8ff3b41835a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dbd39148d6e57f5395cc7e7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd23ca78eb565faa6cac395787;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1c3d9520d05b4c03e93619e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5c642929db980d53a84baa41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb03335d1dc3533ad1782b0874;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8759da648203114a2117cca83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h980bd3ec3c5618f715a6fcdd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5d058446996ddb2c51eebdd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha625dd17075e8df118cac8e76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h776d3ca1cfda8582f017060dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h319eb0d17e25e568698f54a99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd677c2e811a2a5ed7f72a5ff9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb488424b2b4f20fa0c25b500e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dc8785e2ba41d581e1a84eb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfabc145fe384038e164c6b42e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1064d307065b7d79a59be2dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h104bb6d523199fca17146f553;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf77e7926675352e171dd1208c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h259d88a9e13cc37861f671a12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h789dff228550f694d2d16628a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26413b57430149e74e5ae543c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc564924f99e8e438b9eddd755;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d21c05ca859ba1103e9db3c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc511e81e39fe8c57116dc6ac5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29e567331f7cd7c4b265e28d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7ea5e65f85f411ba694d64bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4edcd4edcdcd55fe2d027e372;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2917b666fee36e4e524e87bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fa4ca1cd0505af4074cea70f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48e99476604e23f60e63a0bd8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee9c171ae34992f127b2361f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeb3b34bfcf63e904e335ac3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40d143b8573925a9794b9e006;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b1c556a8398d8536251668e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h474ae9487aca7dbb1bbb0247d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1053573728dd23385d3f05c3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd903a856cc00219852ea0ac81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbff436e7562d979099cd89d90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6699d060482dcde0b04bb5b27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d7bd14df40878c636ba28d32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h351ed8eee0d5179558f19be9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h963352ccbae614619d3fefa9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h291531f6f7289d69516627575;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h517519115f73f46b5f978880b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h798ae12991507abc60fb2186b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cecc9200483d95cc854fad7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fcb7b6c97f405b9a5882a123;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcec10f30fe842532ec990ffaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68fe31ed1ee4bb0b590ff7cab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa953fef636974a2103843276;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ad57775420cb06c0a1e6d06e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb973655128f8aa14f6b227d21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef1b8effd04744193aa0b2f5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb5cc6ad1f476a49790b34ead;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d8a9875d1b5189c6ee331d27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28a93a37c6350c7e115cf034;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb68b798c7931043a3f92fb68d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5131886a97ebe3049f3961c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda7edfc104f929c589e92c35f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h914c2aae6837b93b564033eda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8df6a6c2f0cfc9fe402434e09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haec68f59817a06d446a968ea2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6a8cc9d30022877271ea2d0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba8c833a0da95e5e55b2737dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2f0c6f4433ca463e36c4f42d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h732e16397da4a9bae65fccc68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95d51e42c56f6c86c37feb4bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dd86392db32de10ba7add13c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc25ef9f2050ae4ae9f414d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8567e80fee40fb97f48c25d0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2de23b7779d78d52d37a01365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e58705cb13f960ff29c57e68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39cf06dcb551938b056fcc5e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he85962425ab9bfa797f54644f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b1befa5ca934d717c8240b58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4290cc7090da56e19c37e63f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda64e373de28e14daa8b830b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h841aeb71e1f91a515a0bc50f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa3f27cd6f36df3c5e562f9c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37cfb97ab88bad8e89a984ab2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc10741b5d2b67f276eda19c51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd1dc5f1f64270d6ed9ec8e2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57748106c401cd4046537a09e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h638f5e152c3433eda38671da6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f348d2230403d1a206622bc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h181f8aa8ee0d45e6046923499;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62314cc705375fa55fa26f958;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b1edd64abc07dc1b30b0a389;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1121773a61b30f4ad3d369ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7888ea68213ddac75fbed3238;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96fc453b52ad5e795c09c5036;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8d8d56635fdd7ca36d077be0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12ea40f4b0e1ff4c98cea5323;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5e7d223b0e2f8e7d39cabc7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h336502602b08d3b302ee53fd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd808d4df4c7409ed405ae5e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc96544d7dfa31b13969c26359;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd03aff11cf4cc1aaa3b0a5f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef22952a04992ae489746d43b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h446d635f806dd4ba6be27379e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3b4beb12c500aafbe530fe76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h193bc80364f761f19bc39ab10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h246c21daddbd608aa6e2c293e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd871793b2e38dcac4c37d1a96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec27696111d3bffc605bf66eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfb0ec98ecbdfe1cc892e2af5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8d8d199c27ca6ea6e7dae734;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6067e1d51cc73d2af991f2b4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7cebe81148ce64dfb83bd8c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6df2b573940499d43c2313a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4092412afa6b92b29d92f366;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h458d22c36038678021cc08223;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb384a76a97976a92dfe1d2dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36fce53abfc505b66bacb60dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h758a2577494f362119e0bfed6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1ae350e832909ac07ce2efc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h595fbe9f54a6f8fa430e671b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h470aa4389a455d601040991c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bb72406ef03e1022a2cfde19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h284ef4ba6b240806b89e789de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ad52f05affddd3f2d7aecf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb46f8b5c79682ff4657be1a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h823bdf8504ad717cbe201434d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ef4240f690c58aa0a27e4a28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bee04eced2aadfb5a3551c94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44757df501073a4b1f3b51035;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4eccbeb1663a9647dbf0a11e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83934dd4b06404b64dd937c3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h368f32d480c2617b105d62807;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca8b263636d049cb602ef892d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57d3ca0a530e8ce1c0edd5f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83378a9ce278752aec8dc568d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40a020334f10da1cfaddd568d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h482ccaee182e96dbe45ea1c96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd44b1088d563a3059b56e015;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9d203860aa99534cf3b2c927;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaeacbe59fe405ad91833c507;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf897fac3bcb118ddbb47c3935;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9006ee3fa167655b16fe6735;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3d17214400f7feb0bfa4d9db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc798f2f007bc95d3f17b28c4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37ffba99e493268ab015151d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fc485c3afec5d561f72ce502;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16e0423ec775e90915b47371c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ea1087cc33eee33fed82ecd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h886ae48b451e71d3564615309;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb41fca4508306edf2bb2e2ebb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a4dc0c8d4c6d84c425095d7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ad522eacc4b3b9dc856a157a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3300450003cb8b2277ca7db0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85cf79335e7eabcdd935e8770;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aab60dce7720dbcb703127f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf51e22369ed1762fe1a9abcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a284333575bf5a2efd2674b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7cb739a9a2b63e3f9598ed4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h650117de65de1c0cf88facd73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7bef3c7a2a0ece748c7a2583;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc11d3422820002f75552873b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57773fc79d3c995b4f64c2384;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74573f08d3690560c64168130;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h809ae6c29f05174f141ed9257;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heaa6ce434f935853db9b9ddfa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c62a8c6ee8cd161a60a24f7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb32915d2b8bafd1be5793887;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc746f5a6d54f6d7e43ccd4d25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ed1bbcc1e2c1f0bb09f5dc79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc1821021703967083c0292db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74067df7c8337ec3c8c808a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d6e6798d58dbb48289bf045;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdab607fce6ce7d6e16027952;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56c7b4533fa12ccf8b0ece703;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d02025677dd6a48a4813aca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d095b4ad7aa19808779dfd26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78dcdfd550653bf89e182e00d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heca8cf92cf18ca157696f10f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e8dc62550caa0ba6fbce5b9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd498b9794e4bffd1d32961389;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a719e5c0f8478042a4441d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8210e25ecf4e96945f2dc7892;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47d9723f93c89928a2c11cea4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac8496fef190ffe8f32234fd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he361dac2a365df0a932b1ae82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdce10a2088bb26c8eb850dab6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc06163c078bb804e8553ad44a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h787a5908b418cead4af2ffe0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haea3a6d66de4e1da2331f516c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5761aa356465db46c0bf516fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90d47ff0528590d3637ad5212;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99af332f78ac595263985b4c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b709fd4cc0d0cc1028675aa7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf211bba339a4929e6f871898b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeb12724f6e511408a27e690a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h210655fd78d97d91a73eb1a9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc136e0d18f9a0856910c57597;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h683c43a1651fa0f691cb1323b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3205ad2b05e2ed1e45251540a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36c488ddfb89f1d97403542ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8466475147b728a84e90a6ea8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h529cd71ecabde638ecbeae050;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e30efbd20b29a354e24d205;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73c86a2dfbbd153f2f4a3540d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34c20090a615ebf4e3c5742d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5974ef4acb392126f8ade0c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3016e11440c3f9c5075d81054;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd512f7df638314edb9cebe6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf5471d67cd5f8549e54f4df6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d6b74d4c7e0f51d923121093;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb60a52267ceec1f2cc0cc294f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2270408bf209589b9a31a4f71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d55b9e2805fc2e10d6b15b11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h418ed6a5fa4d321ae52c8f245;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f6f0ee489ebca9c1ff6f1c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h657562de04fa5763a038e16fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0d71fcc62321582946d24905;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2354e6397f7a9da6e0d04f6ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a2a814af8b079344b54a54f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82c5c828988ab30e4da86f997;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08fa5e6592642de3893deb72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd6d7b9052b12e7bde43a7b77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9173d3d295ac848b6705503fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc734040e1a225004211717d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f30e8475e562dbe796e7eca9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h642d28f560871f7411e30ee11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe1c06f3c3ed829fd00634b29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0ebd15ad89a94303e0f1ffdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd269004dad8653d285da331b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd54fb047f5e8efc439d772b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35f2686665b45f32ca04c9cb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac9f20e4d74a68a089ea87087;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22cdc50e0479bc2e4041e8479;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce66ef09b792d7f6da49feb45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67b1a6cbdb4690317221e5a18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb4c16f4a043ca535b4391c9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5ba7f44c3db783db355813a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he858df7a0f445902df8c8a907;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda969436b241370d1b3f7b50b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b7adb7ad369e8b4a011102ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he583191cdbe2dc3cc6b6ddf97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb349c93f3134fbbd918976baa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d01e6a119d972114eb2c9751;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h972071290baa996865c909aa7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8584e526cfc393c26869cb3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cd7ac5132cb33cd191709e2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6fc3e9e86ce14fd6aeb71a14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h936c295cc041c9d5bf20f821e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf228af88b2dea78d752b6bc4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f494f2be5da4d9ff2b24bf3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe14a9dd8a4640ec7c13ba336;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7e24d6d32b26b26c9f858cac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39083601752baf689cb398b46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65405bd551e3832adc8afbdbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7830a139d07f5bfb8a7e459;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2559d7237ba6720c04d3b6a57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hceacc149c7ef97d98a7f31a57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf884a0018fc7379a7d3313a25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdca41c383877bc723de68196;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc798ea537ed6f9d5c48fcabb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2debe857a0f1291fa9bec2ead;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc97cc13291d247f350e9e983;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5783c55b34b824c1a70a4452b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb64a86643d6581cc21bbc1bca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bad27eb6d578be8546afed20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b60ed84ff5957e3b0a14f45c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7384100ed866ff2c1c3f8fd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4f9e73913579198e6b94b41e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c92b755c43e785470487920c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb01d36638a5b9556190ab10c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99509e0630a54e692fd03ab2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4092edd22fe8b3852e82b739f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h318af01d5f3e502810e215cc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h635395ada562d9d273587595c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4df796ea954deae5955e39d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57097c8eec33880206b3fc631;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c30e9614dca1871fbf0d5a5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc75fa9dd25b9605cedddf2251;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3f5060498e8b3123406fb751;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77dc926f392059a86969c406b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2388e9aff7de2de14158cfb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fc58c0469a0b929f6f6ac2a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c65c8dd095b70256015c15e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29338dd6c197bdb1d46b7ed8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6eaa9afbb84c2d4a313a66466;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0823f332a03ec44e91159219;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb40197eb65d5b873300b5e90a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e69001d45b03f4caf8c0298d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61202265a3f332abc58af87e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38e8ae0b7171e50da8f0585b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e22ce1fc74f18b9fc7560396;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf31ed59e9f358b7429a25d3b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ec0ae1c1f1d3559a63f11c97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96476920d6bce9e23155c775c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf01a53d89cc51725e22c91f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h142704e954bf73c8facd18fd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb20e7b6c257c94b1d3a2a38eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4490fc88c362be6e6dad44780;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha73b57dce2de07bf42d669b4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64cc2f7b50edad890f57e8225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab251664ebf31ab4e927f5dd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12da85b62b09a3cc0e84a6842;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1716e22fe26d4e551526a692;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3fefe31415f3e27ffc33d5b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30ec93d7120f30294f8811590;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4182b2846c32953931d1db09a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f8323974510d2f298b27a9b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd701b20f7691a231e4c6ed273;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda6bb99df68fb7a3189dad1a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b206ad8700d2c056910f2d92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heaccfd23d5a0e324ac1a2534a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a445791e633da8f78dae2ac0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h389653d4ff5d6c3b42cf5065f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b876b7b3854a2ce8aa5ca797;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36bf0e085eca408d382150a2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24196dab370d05bafb3dc8f14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1e420d1452a7d01f5b614984;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa0c62c7c7b9a925827863161;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h839a6ad7326f7752dac7916b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75c9314ff310b1b2571f58fbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55b5e3cbce4c1a6d6c48c1cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he51e713302f148b983d0869b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h943c4ad1193e3e4c6b17dfcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12820e844da153641ee78c175;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0d2c2735bffbef780863b15f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1a56ddd9113013defa6c34f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fbdcf662dc97b96ae4c9dc79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ab28825d43522be2c6b6f3ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b9f5cb1504485b7d6946519f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc51eaee07c5ae519b20be3888;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1c0062f3139450e5d2fc071e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb84df41e5216f7020798277e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h645b4c68dd53df4766fe8338f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69469f40cd2059580780757ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h300c2db576b271d52c31cd8be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h927f8ed4c3b4e460f259a30ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb37fed02fa6b05bdafebb2c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c0c3f723008e48defd5501ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d79a46aef08765574d5a7330;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7ee85d9ed1e535943e02736;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb64df7b8cc665d68c5f563eb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ea90d5bc7679b48c9442c72e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a82c5ef1451ad2f6ada765e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7371566df580dca3ba00f7945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf3b7d0e435662413ac9161a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9efda62228d1fa159efd57b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f74db17726cdf0b262abc799;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf24f4c075c1d9b1045518a25b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa5b496db78f5c0372d20dfab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab7fd47efd0c4e1622e696de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce422011d027b2ab80d35d470;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f9b88a298d9df0813da157f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c7acfe8c833bca94c5dde79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd043ac8687ff3750e523e544;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ea554c8622a51e68a477ed50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc628c78c4cb53198500b52d94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28c03378873df1274c27719fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5879d6f28fdf5414be3f78443;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbea5b5fc3234e556ba6c89742;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a5e1c35684898cd67ea1e1d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6612d620881105c4689d3b51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8cbf9810cc545e7e05bec9d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h832d4f9405c6fcd94c3e0834e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h549a66b75117170d4133b4616;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f43ae2d6302450a9d2216360;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f7b3c1d7dd8165e36ece3b2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a50b26ae6f4db548c743bc28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1c22dbbe90271d6db2a0064f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd39dfdcd8b9fd68e3a536121c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdebf570525ad565f4d056b27c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfdd21d13dc28ae0246d75e6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c96285e2704e245e9e06574;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b978e1ebeee64da35e55e080;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a9a0be7f18c2103c7e1faa18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5b1696d5022e3f04097d3e0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17166117e842f91fe0510ee85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5623c4bd157ff8827f8aca105;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1526c8b5e948bb6af2e048255;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haea1761a69dbd9d0b6885f5b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h799c34b9ed485d7303e479a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5374b7af98ed2c100d8b9c97f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h748dbdf08a82e85a1dea311c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a088b070be7cb3dc35b63a31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6bda1faf37460595d85328b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d633224ec28f9ec9ea469adf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40253d1beb713be5aeabbc806;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had222d24b9876b9e7d286f825;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4ee2efc3796f2c7f0fd2c3a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e7dbcb3a19afc3231c072767;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d08a23a60de8af7dfe5a1e7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95347e186f2cbe119df5a8f66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0f7296e5f49dd70ddd7b4027;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac10129563e818650af96dceb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h154fa337c20515e0b899eaadb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36716881439d69a0148a128d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h636e3fec4057cd26597701b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde54ef6f8cac0738059f4e073;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce84c11584b583121995572b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3059e9f0d7b313d8e35437985;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e0402ae17e6338f787b30cdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f4c9e10fb9941024ab3df1e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h244df45ed7b6cf5641560090f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd3fa2734f8d357143367c0a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h721f0f733cdc746c5da7b504f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22edca1d0bbf0585dff16da66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55dc86ea430ac83320c0f8fa1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h274dff3ec6ffca912875f9d1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fcad8a9a3db3fc08d08794ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebe7b82f08ce783baaaebd08b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc886dea069c47e6544890886d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10f5510eeed94a9fe14d799de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25a2e63c456d026454e8cff73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h697964c50123d29d33b31a6db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13e50982a9c3f21d51773945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf4e160512a12c76d94c1e753;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8000091204d27c9c9ae5a13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc67c36da4e8e0f6a6a51a2ae9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecb86a38528b2d251318d4611;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha01ff68857ba7242bdf4a5c63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha87b57f0db09613e5e4398bdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57adb5bf8c2545f53774dd45d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c2d8233c8d0c96d62444b585;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he16e87eb0dbd2a184d3b66b4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heab6ac82b973f081c132beb32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2f77468bd95aa5e02ff7e307;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf569a574233d02751203b698e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h835cdc50a8384bebecfe6567e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10bd2e207459e42f911925ecb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20669332ddfef4f28b59e9fbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h559681af575cf327e008e70c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf64d33ad0e25baf68c982d9de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec68b31200dbc56be86ef7b2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74b6a079740b4b45c3eea6571;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8f6acb2dbcefa7e38efe9856;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h836981bdff499f9806b0bb314;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac55ab74c58dff2edcbcfc370;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19dbdf7b06bcc93c0c2329436;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22512934ef0036bd4d6356fe8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a1e50d5f95cdeaf20534a777;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfaba59a870f8eb1460c46a775;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17e286a8aafb465286843f46e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46b7e73930253c929d6116a6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5479b15b8d4c38b9a2aafe696;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34861d815e100550ffcbd93a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3d9300912eb14815000a71fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9abbc1c0304828f22eba6a94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e0cf8d268829092bada00151;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8ce2f3559c6281f35ff65c0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haab27fab480c9f9a61d99292b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f25ced1f7ed84c4f6b735461;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96f3d08b05fea9b8b41e70568;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haafc76e1f7f2d452212049225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7ea633a62e81c08752f3157d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45311ae60de123ba778abe34c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heece0ef93c9b2e6300e1094be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heff12f8569996b6df3cf6adde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd0652240cdf1c8361dc0ac10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0ebf2d2e91468e36a8ca3182;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94e35bc1d721aa36f4df425ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3c0d67a4af62b9074edf5152;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c3035c008aab0f0cca8dab00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h448ca389353f1d8d73a5d85d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd65c4c287191d87d05b0253f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5eafd5bd36365b876fa81d2f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90671157ab2c3d24735fe9eb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h550afbbc8cd450d9e7a991ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e1a6c7f7bc438f89747e006f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc598d4fccb4ad0af1d227c377;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4d64864d8448b7799d3da15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h318d4fc683777aeaf2ac8c021;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe5c8fbc43339da814356c562;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb796108ab1b7628d4a74b569;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdfdaec0a09ca217ce8cd7611;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a184a5e417bd4d7d2cf2fa0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fc52ed217127118b4a4eb087;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3d9d35e7acf18affe99271db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e54267472153baac8a672d71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c424e586afaef8e5170263c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3928b0d786f13483de5f54cf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83393badf84d10ad841d89c2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd31af875e556a784b76e52fbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84a697ef361eb38dd473eabee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90a6fd1e8c8aa043b2e6f1130;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57786537f5a6dae1619da3c15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37a5bbf5754d759546669bacc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5db954296658d7ace057266cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38677682d0b0e64b2011c72b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac04ba9a30929da011c116d6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d9040caaf1714c0876dc1ffa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7512c5ebe4f7588254fe9364b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4aa3afcdc67e7cee2e319a96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0ed762332a4ce349b393a792;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42db744a85cad54ace0cfbf92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92911f240583492924f0ac424;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h987d78de508269c675553767d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcce89c878b69688fff0980937;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h705fcbc123370ab619ccd5459;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e8c961a0d6286d84871954ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha22ca4286128592719166c1e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he03ca61ddfa00a2257a655dc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17fd7681b1046b925c6d8c79d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8d2dd13276b96c3585660a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50a69837897b5bfe867705033;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfefc8902bc8cf84d76bb71fc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdef7cc41c2f323c6b0393e2df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef9039d83a7c599ec5649248d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5b5e6757133f3461f0e27931;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bacdac46f9aa8e9f4e21f71c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82085986e2493429be2910516;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6511a840de16074a0e9170843;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9220f4f366c4b032152f70101;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h592a93b92f3ef1ac3b264973d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddbc888e4744ad3803b9a11e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf99fec3167b7764b7fb34a7cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c26a92610f205c8544cfc8f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2aee7c3d23b24d39393519db0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dbf93a6cf7c1000d5d58841f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf3e9e8b77637f4e19ba8255a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cc72fc6469df72d45d0dee88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12626092c478097bd48e10fd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8b510374aeddbff5bf2ae891;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10cb0d560f84f20fd25808e6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd24e64ff93c0c6f5b444371a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8c2f640f00132377520ff061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39e509b9347a3c6eb5e42cbbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb7bab6c5c431da1ca14ea16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf72e242ae1fc48a4c06dec5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b66534e3d486c9f322c29919;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41fd98ea7b5cdc529a738a33d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71a3c02ad561d4b3897dad38b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84dc2e0699ffcd67168e8585d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc93d03f71b70874a902c17143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f8345c4eb7b192d931c1f959;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f00a986768bc0e25ac653df7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h276dec2d0f19dc5b59f5b2f1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf38d9f714b37364f3591ec0ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5832ea0d01ff6745989c477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8527d4316528fdca90be9f2f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5baf5ed6572d622038f6242a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f264b231894e7383eba61be2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b54c3e7039cbfe4aa379aa3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fa701b4d13362a1d74cc7196;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdb4e821cb1b813b2dbe831c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7acf0a973f70c6abfa440f513;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84c3012ca96e07a566f0d925d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd89302b7f0d99d863eaf1d7c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbef8ec549a1c377db78c41c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf103ade9f0773f7d988c1f96e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91de29bef9f123267189e2f8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha59f360b82f63010731b3b34e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9bbffdc5c9adae8b6272d9b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he78ea08738ec0c9839b4d7dd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65f0745d14549189c2f7af04c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h267bea96a972ef1849d66b4a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bc3d808e40ad3d6c9f226f97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h366494d2df19c9b0e1c26d1c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0080f3d3c14c05d8157e535;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e56b6ace14aae01b5a9fe63e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ce8a058831b3b3fd10ab71b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e98f7205936b04d32b1b7de7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bda08a2c32ef9de0c643852e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h246fbb08cc1df2adc81ecb80a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32757ac47c851dead6a61e75c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2291637916e7c2ec9e8586dcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c7ea2ee8a44b9108de3eb7ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8be1563c4f6c7b1666b6a1b9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb41e2acd26cbb416ff57c02e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h807a69e575a24a93781b8c67a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1c28490d5d382aeadcbfaf1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5808d178ce9db29d4f3dfc8e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ca039c22ec16358594672176;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h525522092daed587363b81b85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf06396940ba0ca9cd76a2f70f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e0032c2d00faf4ac49c9e986;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a4e8d2daae4e3138f2b08f02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h427490841ec0f9aa73e23b8f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbfea53253d1426c8acb7334c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he098a29962e6dbe7470341305;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb2962dbfe4235a45d3ed1cc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6db64f4548b7cfc243b44f9fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h398a7db509ab3e7036015f8ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h668ea899bcdfd4975eb88190d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfc89aa5dec9715eaa00f36c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8b200a37ca331f92b526e92c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5487f3870f5de814bd6988063;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e517bf60e49869e27e9ffbdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83a41c1d0a063922e0bba9be4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h813150dd435ae38598a6345e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c25e51c406cbb6b97a6c5c44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h572ef68915917f04859c0a2a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7985cc8295242eebe060433c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95dc4821f19110ada93def169;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43675802bc45cd149ddd881e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78f62f744fad315b5379072e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha75d8cdf31756fb86c9c903da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h753c04a2f98412b2e5eaa0fbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he56c9f006990cb6e18b0d0b19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd1f3326652c6fe93fe94c490;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb724ee496cf110598a7f1c27b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca61e4a3e4e1f6df6f0c9570b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca5b50df3808cb53d000bb213;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h547626fedc683507ce8661e70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h570d83696893575f739ccb2fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he31bc944a3658cf778bcc008c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44697ff397e28643fe544fb4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab1f306d50a6c9cc6235e196a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb28fc2a22c748f3f335d184bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d68f6556634e99ad01cbeb95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha505f6bd0a94c32db620465c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39d9bb978a579c1418ea25040;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h967c60f03e92359040b6d9b2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37d33d2120a1e9c1ab6e80256;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e3be4654f7f6b857f63df702;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d81d9f15dca31deff89436f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c0b1f3c0bae3e14ce31b3bb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea397a42024bc901f9d132a98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17477a9ee2085b9537fb67acc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fa27e3b0c38d6f0f3e9369a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7ff314d65948c71cd261cd2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ea686ceaacfe043c9c582404;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h687cf6ab32a3c0c4c147ba9df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11b9526c60ac703a4a72eb41e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48bc054d7543de6701573be83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e71bad33fa9cdc9f40bf9970;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf7f5d47d7faf6099d3bb014c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26543859f5af26041915db8cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4af5c598413cee48cb0406f2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd21e0875e360595577fb55210;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76643961f72ad51eca74fddd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c46b4fa5b46277e433f1ad36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f144b350bf86b988f7fd56f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef31c46ef1459a65706c94fc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h341a37eb67c885cb608685981;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a3e8333ed3d6330280d6ae3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c896ce7038f83ce32c5527bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47be62d399966a93e473f3492;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d3232895380e03ffadbe4920;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h294f52aa0ffea1b2b217807f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9063209606586ae63bbbab1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e0c83bfa4bbf7ce93d41e143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffe8a5ebf89603a9e4eb632a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1940c179361cafbb9f60967c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a7813fc5fecf8b801cc33f24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90ecd66c2d0ca01ca7d60ab75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h610aca4e5cb0233db683479c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddc27627de8f55ef1df4d0b1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0d80199b21b2fa58dcd2d770;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf0223e711bd04a6b10eed62c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e2a56bcf40c41adcd464fb3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd3d06602b8fab1a1611639fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf23fec5b24c3cb940a9e8c960;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2931ee4de29ddb11af52948a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f90382616814978aeffb2198;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3aa951c12178ec43bab16997f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb6c0ceb137d468345c17a4ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb996b6ef21137b504b5a955f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc93919c14d85e6306385c702;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc82219d7de1b35e596b6ffbae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb78876014df32b22022612a36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h900a4b85c1e736fd151e7d715;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1ffdd11f2dc1b177132cfada;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha32dc03a50cee9a24af57c1fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fb266b121a8b634958cb2f11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a7b5364d0e60f7dedcd1bafb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h425fbd0912f4856eddd79a9a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2f6515b5f90433a544184e8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h832db7c468153bed3550914c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb63d63f227a10da8dd2cc9747;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53a2087f0e1324596177bdb3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c8f0f7bf050743f2f6993950;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3e9b281c6c69196033ddd680;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h283c04843001dffeace0fddb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcf1b19e3fdd810eab656c9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9491757980f44278567b2df01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h537bc982fd94e021a477f443a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dadf74eb3587ff55dc1f36b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71c873a3a9dbb9498c042ae54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15f444c22ec371e59145dbd4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc697f7cc549fbb735547e020b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b55c694991c74a1ec0a01874;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5305bf6a90f36b57ec9365dbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb63046551619ab27c231d853;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he73f80f2876b9ec8379e1fec1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7b40aeb1a5579bea11c238d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd90865fb19cc18b41c86a9a32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f0c719fb9a2cb225a6a82939;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4112d3d6849f7a0678905244;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haef6e5a9b0d4130da455bdb09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he79565b136f87df592c7c0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dc3e68e20b41c25f59426271;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h289e557300682af1cd7a7770e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a10c8e04271e92fdf5eec186;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h714a230fdee8ee916312a1462;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea83bce75450a83554294df9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc3c3543ba023925683c7c955;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2694224cf84aeb6f790e6a5c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h238622d98067f97977dbe4f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a8de864aacdad72b2f3ea423;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d7039cdbae771e991af49382;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7955517daedb95f9cc7832307;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c1d3d5a3bc8bc7b934fb1d28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haca2ffc682f1d8a1ac32da01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda2c11ab5f3fd420b6f26038f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98d58bef81ff9f33e19003120;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h486f776d97f641a906e27c121;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f23f32bdb10b79b576bad42d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa003ddf4645e0ad01a5be5bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dadc2220bd244df77e743125;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5fedff52536ad22bb539d2a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51f8cca1dbf407e85ea68bd09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7a768988526d23737433f7cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbf67a5f80ffd71c35941db52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9696397034fc60612c7640110;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccfbb4a2a891eb48568897b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4164c74a5535af0a9552d0b06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91922edaed04325170ba33da1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57bfc029ebd576359214e792c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8d942612853235fe1b6c5080;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fec30d65aeba08adc3529a27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80753450ad6b93103c711fcb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71cf3b02fc43f0fc3b2e57450;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9e6063d232f11f047f2ac5ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h396cedc660004498526356888;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1eb2ccee6672709b76d0137b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc409300d636c6f09f619857a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha596b029f3d5f03f83541d884;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21a1516bdd001529f00ba695c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h779dbba1a9411cea363b588d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25c1d40910110273c5de69b05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62aae38fa3c1bf2bea8bce74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h568b64f1a477f1aeac22d05ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38bd9710574eccb8c5c0018fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74ad68c2a02b88c9f264c32fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6e7fc4343b9648726e14c1e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcf95cbf316f09bfb6f68dabf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he520e3862a0288c8e17a92d32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefed6f55832ac825c305fa144;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab921be78f80ccd75a77bd608;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62cd2de21ef1b5b8a934f5b55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h269d4f2097a62da995a2664e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9bbda730d2ac36bfcfe621b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4006e2776f3d5c08f593b4396;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h565479922a3f2e8825fb5b756;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h431f28e73a03fece7bb1801e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ba218d950cfa8a15c2c67e71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h143c545b3bd7456bdb436c81b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h401206dc892a3097ca7486e49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0fb3cb61eac4a7ff58743308;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha69a4ff5287f11b45133f5474;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h466361c46ca60c4c9efe76037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2022087b3fa7c7b7b06872618;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e3c895e5cd4ba09ea48a7833;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32ead1d9e0e08488776bd0ac5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2438adbe3ba3b12087cbbe82b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h470f9e5cd2de96965a2554ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b60314fff21badc1e1d13549;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef973172622b6cda6d5672ae4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1918ac84ecdc915dd908ec4f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca90b322d4af17e54b4c4188f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf51e541ea04996cf081bbdcec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa97412c6cc68d40c9875faf3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1f41708eca8f4512a70d8b7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7e5409675e5fb9f3e3f66658;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a5c6a9af19115821eaa0be02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c348a2ecca1435f5f833dfe5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6db031121e51387c8a00060;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0b91b18df11919d99d6a4c37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he56afaf39b74705c7e23d6318;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc47ec1783c235251b1e060c1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h899cb6ba4bd3b3825bc4b6d2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4612ee552d26d8f60c5220afc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4d2027afe1c288836de5cbb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haae1e1eb1161e12587bcef169;
        #1
        $finish();
    end
endmodule
