module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    compressor_CLA54_16 compressor_CLA54_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA54_16(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    wire [1:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[1], 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20,
      output wire [1:0] dst21);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [13:0] stage1_0;
   wire [16:0] stage1_1;
   wire [22:0] stage1_2;
   wire [17:0] stage1_3;
   wire [34:0] stage1_4;
   wire [24:0] stage1_5;
   wire [18:0] stage1_6;
   wire [18:0] stage1_7;
   wire [25:0] stage1_8;
   wire [26:0] stage1_9;
   wire [18:0] stage1_10;
   wire [17:0] stage1_11;
   wire [25:0] stage1_12;
   wire [25:0] stage1_13;
   wire [17:0] stage1_14;
   wire [23:0] stage1_15;
   wire [16:0] stage1_16;
   wire [7:0] stage1_17;
   wire [7:0] stage2_0;
   wire [2:0] stage2_1;
   wire [7:0] stage2_2;
   wire [8:0] stage2_3;
   wire [11:0] stage2_4;
   wire [9:0] stage2_5;
   wire [11:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [6:0] stage2_11;
   wire [8:0] stage2_12;
   wire [10:0] stage2_13;
   wire [8:0] stage2_14;
   wire [7:0] stage2_15;
   wire [9:0] stage2_16;
   wire [6:0] stage2_17;
   wire [2:0] stage2_18;
   wire [2:0] stage2_19;
   wire [0:0] stage2_20;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [5:0] stage3_5;
   wire [2:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [5:0] stage3_16;
   wire [3:0] stage3_17;
   wire [3:0] stage3_18;
   wire [0:0] stage3_19;
   wire [0:0] stage3_20;
   wire [0:0] stage3_21;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage4_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1406_5 gpc8 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage0_4[0]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc1406_5 gpc9 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage0_4[1]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], 1'b0},
      {stage0_4[2]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[15],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[6]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[16],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[17]}
   );
   gpc606_5 gpc26 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[20]}
   );
   gpc606_5 gpc29 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[21]}
   );
   gpc606_5 gpc30 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc31 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[48]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[16]}
   );
   gpc615_5 gpc34 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[49]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[17]}
   );
   gpc615_5 gpc35 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], 1'b0},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[10],stage1_8[17],stage1_7[18]}
   );
   gpc606_5 gpc36 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[11],stage1_8[18]}
   );
   gpc615_5 gpc37 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[6]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[12],stage1_8[19]}
   );
   gpc615_5 gpc38 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_9[7]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[13],stage1_8[20]}
   );
   gpc615_5 gpc39 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_9[8]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[6],stage1_9[14],stage1_8[21]}
   );
   gpc615_5 gpc40 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[9]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[7],stage1_9[15],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[10]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[8],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[11]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[9],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[12]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[10],stage1_9[18],stage1_8[25]}
   );
   gpc606_5 gpc44 (
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc45 (
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[12],stage1_9[20]}
   );
   gpc615_5 gpc46 (
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_10[48]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34]},
      {stage0_10[49]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc48 (
      {stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_10[50]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc49 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_10[51]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc50 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_10[52]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[17],stage1_9[25]}
   );
   gpc615_5 gpc51 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], 1'b0},
      {stage0_10[53]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[18],stage1_9[26]}
   );
   gpc606_5 gpc52 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[8],stage1_12[16],stage1_11[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[9],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[10],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[11],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc57 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc58 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc59 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc60 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc61 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[9],stage1_13[17],stage1_12[25]}
   );
   gpc606_5 gpc62 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[10],stage1_13[18]}
   );
   gpc606_5 gpc63 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[11],stage1_13[19]}
   );
   gpc606_5 gpc64 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[12],stage1_13[20]}
   );
   gpc606_5 gpc65 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[13],stage1_13[21]}
   );
   gpc606_5 gpc66 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[14],stage1_13[22]}
   );
   gpc606_5 gpc67 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[15],stage1_13[23]}
   );
   gpc606_5 gpc68 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[16],stage1_13[24]}
   );
   gpc606_5 gpc69 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[17],stage1_13[25]}
   );
   gpc1_1 gpc70 (
      {stage0_0[48]},
      {stage1_0[8]}
   );
   gpc1_1 gpc71 (
      {stage0_0[49]},
      {stage1_0[9]}
   );
   gpc1_1 gpc72 (
      {stage0_0[50]},
      {stage1_0[10]}
   );
   gpc1_1 gpc73 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc74 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc75 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc76 (
      {stage0_2[48]},
      {stage1_2[17]}
   );
   gpc1_1 gpc77 (
      {stage0_2[49]},
      {stage1_2[18]}
   );
   gpc1_1 gpc78 (
      {stage0_2[50]},
      {stage1_2[19]}
   );
   gpc1_1 gpc79 (
      {stage0_2[51]},
      {stage1_2[20]}
   );
   gpc1_1 gpc80 (
      {stage0_2[52]},
      {stage1_2[21]}
   );
   gpc1_1 gpc81 (
      {stage0_2[53]},
      {stage1_2[22]}
   );
   gpc1_1 gpc82 (
      {stage0_4[44]},
      {stage1_4[25]}
   );
   gpc1_1 gpc83 (
      {stage0_4[45]},
      {stage1_4[26]}
   );
   gpc1_1 gpc84 (
      {stage0_4[46]},
      {stage1_4[27]}
   );
   gpc1_1 gpc85 (
      {stage0_4[47]},
      {stage1_4[28]}
   );
   gpc1_1 gpc86 (
      {stage0_4[48]},
      {stage1_4[29]}
   );
   gpc1_1 gpc87 (
      {stage0_4[49]},
      {stage1_4[30]}
   );
   gpc1_1 gpc88 (
      {stage0_4[50]},
      {stage1_4[31]}
   );
   gpc1_1 gpc89 (
      {stage0_4[51]},
      {stage1_4[32]}
   );
   gpc1_1 gpc90 (
      {stage0_4[52]},
      {stage1_4[33]}
   );
   gpc1_1 gpc91 (
      {stage0_4[53]},
      {stage1_4[34]}
   );
   gpc1_1 gpc92 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc93 (
      {stage0_15[48]},
      {stage1_15[18]}
   );
   gpc1_1 gpc94 (
      {stage0_15[49]},
      {stage1_15[19]}
   );
   gpc1_1 gpc95 (
      {stage0_15[50]},
      {stage1_15[20]}
   );
   gpc1_1 gpc96 (
      {stage0_15[51]},
      {stage1_15[21]}
   );
   gpc1_1 gpc97 (
      {stage0_15[52]},
      {stage1_15[22]}
   );
   gpc1_1 gpc98 (
      {stage0_15[53]},
      {stage1_15[23]}
   );
   gpc1163_5 gpc99 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc100 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc101 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], 1'b0},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc102 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc606_5 gpc103 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc104 (
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc105 (
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc106 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc107 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[20]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8],stage2_3[8]}
   );
   gpc207_4 gpc108 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[3],stage2_6[6],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc109 (
      {stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[4],stage2_6[7],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc110 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[5],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc111 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc112 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc113 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[8]}
   );
   gpc615_5 gpc114 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[13]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[4],stage2_8[5],stage2_7[9]}
   );
   gpc606_5 gpc115 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[4],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc116 (
      {stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[5],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc117 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[4],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc118 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[5],stage2_10[7],stage2_9[8]}
   );
   gpc1163_5 gpc119 (
      {stage1_10[12], stage1_10[13], stage1_10[14]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[6],stage2_10[8]}
   );
   gpc117_4 gpc120 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc121 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc122 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[5],stage2_12[7]}
   );
   gpc606_5 gpc123 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], 1'b0},
      {stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[6],stage2_12[8]}
   );
   gpc606_5 gpc124 (
      {stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[5],stage2_13[7]}
   );
   gpc606_5 gpc125 (
      {stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[6],stage2_13[8]}
   );
   gpc606_5 gpc126 (
      {stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[7],stage2_13[9]}
   );
   gpc606_5 gpc127 (
      {stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[8],stage2_13[10]}
   );
   gpc117_4 gpc128 (
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[0]},
      {1'b0},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[7]}
   );
   gpc117_4 gpc129 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13]},
      {stage1_17[1]},
      {1'b0},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[8]}
   );
   gpc1163_5 gpc130 (
      {stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7]},
      {1'b0},
      {1'b0},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[9]}
   );
   gpc1_1 gpc131 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc132 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc133 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc134 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc135 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc136 (
      {stage1_2[21]},
      {stage2_2[6]}
   );
   gpc1_1 gpc137 (
      {stage1_2[22]},
      {stage2_2[7]}
   );
   gpc1_1 gpc138 (
      {stage1_4[34]},
      {stage2_4[11]}
   );
   gpc1_1 gpc139 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc140 (
      {stage1_6[18]},
      {stage2_6[11]}
   );
   gpc1_1 gpc141 (
      {stage1_7[18]},
      {stage2_7[10]}
   );
   gpc1_1 gpc142 (
      {stage1_9[24]},
      {stage2_9[9]}
   );
   gpc1_1 gpc143 (
      {stage1_9[25]},
      {stage2_9[10]}
   );
   gpc1_1 gpc144 (
      {stage1_9[26]},
      {stage2_9[11]}
   );
   gpc1_1 gpc145 (
      {stage1_10[15]},
      {stage2_10[9]}
   );
   gpc1_1 gpc146 (
      {stage1_10[16]},
      {stage2_10[10]}
   );
   gpc1_1 gpc147 (
      {stage1_10[17]},
      {stage2_10[11]}
   );
   gpc1_1 gpc148 (
      {stage1_10[18]},
      {stage2_10[12]}
   );
   gpc207_4 gpc149 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_2[0], stage2_2[1]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc150 (
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_3[0]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc151 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[1]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc152 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc153 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc154 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc155 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc156 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc157 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc158 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc1343_5 gpc159 (
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[3]}
   );
   gpc615_5 gpc160 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_13[10]},
      {stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage3_16[1],stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc117_4 gpc161 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[3]}
   );
   gpc7_3 gpc162 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7]},
      {stage3_18[1],stage3_17[1],stage3_16[3]}
   );
   gpc1325_5 gpc163 (
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage2_18[0], stage2_18[1]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[2],stage3_17[2]}
   );
   gpc1_1 gpc164 (
      {stage2_0[7]},
      {stage3_0[1]}
   );
   gpc1_1 gpc165 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc166 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc167 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc168 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc169 (
      {stage2_5[9]},
      {stage3_5[5]}
   );
   gpc1_1 gpc170 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc171 (
      {stage2_11[6]},
      {stage3_11[5]}
   );
   gpc1_1 gpc172 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc1_1 gpc173 (
      {stage2_16[8]},
      {stage3_16[4]}
   );
   gpc1_1 gpc174 (
      {stage2_16[9]},
      {stage3_16[5]}
   );
   gpc1_1 gpc175 (
      {stage2_17[6]},
      {stage3_17[3]}
   );
   gpc1_1 gpc176 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc2135_5 gpc177 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc178 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[2]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc135_4 gpc179 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc1163_5 gpc180 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc181 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1163_5 gpc182 (
      {stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1163_5 gpc183 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[1], stage3_18[2], stage3_18[3], 1'b0, 1'b0, 1'b0},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc184 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc185 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc186 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc187 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc188 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc189 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc190 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc191 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc192 (
      {stage3_21[0]},
      {stage4_21[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor_CLA54_16 compressor_CLA54_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7a58852e9e4d08b4affab80c4540fcd864d6d0109e96f0bc53f9915e4ebae0b16d2269c23fbd852c35fb14f8ba3e462b415a4da40c3dfec6fdc65add291eaf87f69566d3ee25baa29c8c688d8a8a21e972e57c264e92679a2ec61979a39beb497f33fe78f789dbb7e3bd38f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h31b802d41e4727f120421e80981b023bf3a4b1d790c3e44a2fdded0f160e29249a53e6dcd9382c48437374df031e9ce27e59705a1af94f919ade31684d4803227bc7eb148c75b16930fae542f8016a35334335b269d9c725daf94c9fc6dbd0a24d198b5c53066a8d9bd2ab42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8acaf65fe44630b4111549b507451e726e92c3ef77df1754f7b7a12e31f0b3359104b09d8154e22a1cf3f367e1f63494ad8579405dc3523245b9ccf3b1422fae565c28e11228ed2c2df955a11b3afd7808748d28cf4370edba9f1f1e58e3600b2d8ecc50e29fcfc820080b87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h54a7c9901413f3c1e3fd5d980488e74862c045c4748fa70f64d997fd43226a48af03d454073c1b782240832033f32a280eaadc45d48822e3b6de818e10d6edadffb55fc0759b5ae1ad27ce86325bbbcbfc17948e4d4f76073a142b66d6099597bd9bf1103e728605bcef01cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd14430a857e8fbbc5b9c8e4804a92c0b124a5a0e9e7e5c238b2484b7bc482370f415c1d9145e256bed3410021157fdf99bc738aee723173ffad56c5afd20fe17c5589c931c43d24c71ed1292cfae8589d67edadb284c8c181e0fbf28909d555acb9cfe2fde5a954ece0dc91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he759f5d9e4ff013e30ae42c962035bb73f7bc7bf14e4e5da1abbb9095671d42a6fe214110d9b507eea5f21b1fcc592cdd4cd7e3d5b048e0cceab4bc01b32e79ab33c7c6b0baad246ffaf3c9bd291d378fd259e496c02a0e84fe1821d9f3021785e8da10dd8cca82217a4f036;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h52a5f8172f233264700342e513ad23c0cd4b586b5b5d64c489c1ca033c0f8e0402479edf9a2e8dff624d3aaeada9185c43eef7690058c5b296023afa89f51b70ff0911ea13c8cfc8429303811e2ea780a018c3af492c915936aacbbe06d60d70b451ba8466a80e916949ba98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd4bb9f7907bb57e74b6dbd3398cf4599c3e169a6d95ef3f049db4fdf7f7a96c96a9926b6dde81e384befa6a90fba20b51364c88293be94a0422def613c5f458a6e88bd190082d732597acebb343e0ae14791e5efcb6af379bd29ab90c54cfe8d268a6bb2202182b06ce50aa8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h845ad3ab592098380fc672d8477abbe3f636e74066f65e2c242a8a434f0881979fde91ed9224d8d84acdb297348b863b47afc33a6a3acf539300b97857b62a3864ee94cbe16b30a58705b3c8667185908bb30eb29e28091718eb2741ecabe06edb56a50ddd9791a7c29c7f43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he8806421364b742f773354c3456a5fb2455336898ea97ddf74040c795c97dda55f6af027bb652b317a4dd70bc1e738f1ba82bdb7e0ce1a69e133daee09291c68621e1c922c8edf35a53d9367c35fc01eaa38d7828b071c1d7619966ce9785f9b1c3c0998d180979e7db87e43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7fbcccb7d98227fc454c497f41fab6d3c4539377cacf7c27ef5e07ec83dffd23b485d2621b9cc06d0eeb71a6257892f2c598c94947eac2a841ba57dfa39417b1d34de9cff89be3892bdfff21570047ac8e52f0a056bad0f37b73b43c357ee0515f26503b7b27f66958590f30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hda625376b3e4e96649dfb88099e1ad079573a096ba03d773ca0f497cbccb8d5bd598a4d6f29cce256a6052863b662dd05b5912ea37b442c155a5bde7835cf4bd77869b522789bedfebb162f40006dc5b20e9902c2f6ed6154d748fa325c93610a893c57947ca01306cdb8c46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb81f7d1dcf121547f8a3e61cbf421c2c111bc1a1e2837631916efb915d40176f4064fdd3df9bf500b14b8571c5718f8407903acb36b285b59bdf90d7aafd2294c3b88d8eb5879bec1006532113852bffbfbe60200cf18e2575a3e0f48792595be38667e1fe0ba711a001c497;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6d57dd24ab64f86c906662b738c5de88ea72d8095d6346c136b20a62ffa0a04df2d9a7e694532e2ba41709dc85a6228d07de3230cc01423e1139205eaf6d50dd185e402694275b63c15af48a39ec22ce6f3f4e2d49609a014a3dfc72211940239698226ff35879b7e805d324;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h50ef91de08a3148f301f72c53de1d161e1fcb6bb3a0e44b25b4a63108a7fb66c219e4ca3556520967bd82c1b7a78a7e5ded1015eca244997e2f018770f111f63b44a0bc30e78bf6c9920dd671f5ca96a059287c2d80a4b6416d128f1d989637be44f9e9fe63602fbefeeedc6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hec8957557a55999bdd8fa03d462fbf71c4e38bbe831dcc2b8c34fd9993fedd85e547638c737592096062ca393b7060d377067086bb2e37e69d8eb5ec3336b90262472a3e142fcbfb92351abfadda7f844841a2453c83bc4776cdde0927782581cccf4d8f8e43ce07e33dd67f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha7aa835594fae277d1199e29628160c5d5d29e755f7a269145bdea59eff9a6c68aac7b656ead098925d2e2656805f7007581e7313aa95e46f2980f54d10a6fc4b26fba5d2d35838b4c472598bf4fb7f4b2d636425944d3b9f203b49f24578c0e4df6a875f379c1d3f64d4a5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h16f6c844d0744c42f40db9483c13f45be4e400f621c0705e063751129a59a95accdcf556dc9248fc543d8632e37bbfe9c5fde49721080e3fad8a67ebaf30a521a04a24a4169a77b670d794e0ec63abd4b8bb4e64c0b8078d5b59c1bc57caa26fd9bf29bc60158c262a2fda0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h74c769825867667b33cd8401a71b1317cc0eadf4067936e8ecbf1257c7c22b43330482f0ace6e3bd63db0e02ff2983bfc70ad01f5ce13cda4002c6c215052662df22d277ee50ab1db6c1b280612edbd3b562e0c0771d8d1e2ea6dafd7f51029a98fed42af7288801201fdbed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd0542a37938b6324d1debdb601dedce8ec045f2e87e2529da0accaa92a5718e7e9e59446b21e26b354549cd37d3259f449bb7db6e8c5877bc3c9cb4cda4b3757d411d9b94f204edb85d38fba24fdade2ab5ace83d45715830fe4d804a1215c91efe0e170cde07f600b86b75b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf8f8f364ed2dc151d1738a53777446c82d2aac4f2936510069ae6ae2dc797f858a3e78c9974b118477c59ae9d3681a7df2dd49130596aa72e5f8830dd8b88bc6f64d9a7684ab16c207d3697054a0edd1be95660428d2af576569011bac10a6cf30dca5796ec8885976b1d051;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha521b8f6b14d96ac1b5b0dbca8390a96b8faa9acdf9505467d5af897c31fac7a97bd594ba031a61d88f272e5e1de56f01e279e9ee06e752248c32a057ccdcab6559ac29d2acce9d0f040002c6efea713bed07da352cea9a4b312f5d05823bd56317c3946e9b539bdeaa24f20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbe989b76638458da38cecba3d39b7e54cd332c82e34f015b9c5337e1b6f9c10b277233428c9749192ed79df2b699077935c825e8cffaee52efec1adfdf7f8fc461dd29a6fb97cbac79f14c3c1f6ab338b5daffb61397492aa63e8a046530e5b51046d5d5608deff058dc06f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9626170071630513f5e856419541e522fa9d9f631b95909010d68909570de0bda378feb71ace4d0a85fe998e90d71b96a36436596324a607957e7c09f4698b087b96ae49ae6fe02d7ea41e0ba8b916123042faff7d57298817ff1e1ea7f4240ac08f20cba5528b39de4292c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hfed2944c4b7b491d1878dad5f5119e407d513a843d2091707d26bec992caa321ceb94c5caf875fcc8f8be5f45a8ccfc74b6e92d521a476d913951fba6e646a02edf7d335312ad815e91d084278433e0ab7f52c66176fc4e9d824d0b5a6c134efa3d0e9cabd1c9af654575133;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc2f36e961f0b99ef40ca872901211b3ef1dcbab11e9d15ed84d1bad08fc7db09248c7c1ef7ea1fbed7362e69eb6aeb2d09323f40978f7cb821573a768f41b97aa1a40011f25df1ee4504b9f70a385c4d06bf347d85289a04b6ec808c993250b0f6758e741b8b8971fb5905d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h99071566a97e288e05ca4e287bbb8bc37cde79780fba1a1d49ac61258cc55710237508a7be209f0c71a2e94467cbcb739e28f998dd0147ec83ec1c06976b301545ab5107a3152e4804a7e16d11d5f2ca51204352d02f7120f776917e953d1ae3f49f69412638601f4bfb8235;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h482e1dba5893a4efd2bead5dd38a8cee94dbfba4ce99f32764c78538bdf92fdcfaeec8b0aa6b6be3ae06f770b01d826633976c3ae1fa70a27d5f41725ca6a05e8fe65fb707d7173ea89e83d785aabeafe88ccde1f38ff9c46ba668c8743dabd1c40651bc69636964631e3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3118229642c39787d8d6d68ff5d1e3b068e9edb4340f4737293a9553acd30259b68179645037f5aed5239b5ef198f2ac50f429e866be15fb1d01bf08627121aa52c1104a16719930eb68d7c8f4c919370ae494d43b012f9aac6b9d63e240a7b262baa8ce92793f3e5587a07d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h22d960922f0efe3bf71f5cbba8c6a24a47c1627e0a4e40f82f91a524787e21b8e9ad4d2c084ab350afd2a4d8724a900c87a9ddde49005509ddbbb1a31bf9cb5b9ce7a1b22c41b5ac427bad01a4e1173c9246fad5c41f1d54d9ca7b96a2fb80edd672a79359c56b216ba56f37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h97e03202c3ebf2cdb2a9d3deef0e02578e23f1731a727985762b6d8a3d3c6045fe7b4b13ad93a4e6fb566e2b249dde89cb9670796c53dcb5fbd478818a22a18c915e02ff21e88ca6f1964adf0079b7d8e5eda2f299581d09f9e2e471b779bf9053305d61a7fdd0e4bb875346;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3d0321cb0f4ff094a7c2a7d5a31f04c40442a7b996608762cf2f9d5cdffcc54dcdfead0c54b54dcb5a3236870d37644bd35b5fea276b318d46c28afc2a3a7ac3dae6bf94c2a049d322cd75157ff7e1efedad5f7b0b8b6b083bd96f13a47816e67b4568ec21a4894d3864ef33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9d5308dbe95a0647ceaef1ef7b3a9b8554a426b04f805caa3b55c28a6b2ca4d235dc6021731a04d8f5816d5a59632c8411bd6050170193880f418f798b868b70f7fd6697e60d8a8ea051095885b3272cc436675993498be118cecba8554cda30e5c0fd369eac080ab0deb0c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc2280a4df4008e2ada17efd9a51da7231834261c71ed3f84166b2c3c87ce66c42e7f00f179f63482218ea1b990c0eef69498d9466de05d7ab39e8d561ffd43662818ce62ef88f9e8e0ebe7c9e3397cdc2192da1a8130ef2f8651913968ed3a42a5c80e66ac3c19a3a610ce7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7bdd10f06c8f2c273406f08f7e01bc2f4f354af744c05e9b3d58b2c4729260aadcb7b2a3bf3d3260eb36b06d4a9e92b5f4a050d4b49f4e3a5ee5e26c227970e480411df7dc2b33a42ba4757dfb3b31f5e1340933301a5a4ee8d092fffaa06e2f887d98eb48077848630bf8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5ac13111c18f6883f29e53be57d193791bb3e2b376d969fce1ce0541c28fa60ac4ec6a6753d2865dd538c366216a23e5e5b7ebed94771f35f0459a9417f961e0240da8219cd4837ab1cbcc2a442650ed1172b702ab00d25d5fdbb84140785538c2306c810d91820fe96dffe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb8e57816420d47c9adc43d3e93eeed1548909ede5bb54ebf2f70eea346f63f9418081cf733f1cb60781fc4552773445212511a125490ac82b43d0e633004aadd888a55c0936d9c3b5dcf656f315213071e2900c8708d497308c017b7e948c0d36cf316c2a2023420cbfe5cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc9e818ebd6fd7eb671ad2bf2c09ea91596f2eb2ab93cba7b44d4472e3e8802fbe0b8cb3d414dc185ee52e927330a0ac18151864086776fe227a75a95677c016255a95a317014340ca23018da3b285639442889ada58503e2b8ee916e81c36b98e3858222e197f006696e7f49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7f678822d826271ba0f6727982d11f93b4b67667a4a01798283beec9423b845b7a2addb5c7d9bce3d483fba35db3740ca746258bb879f5e8e37e4536523523ddae1ac3094198129530ff0580304065e170579949bd5fb35152fe60c9f998f82efe6067efceb190be623967be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9cbb33f328daa79dc94fea1260ae168f5f6dbd3b2619ec1a0ae4d40f11e1f16eb9a10bb9207c96a015dcbd59a7a76e4ebfd9683ef9c1f05f7e94a4f644baafe7358bba50f4ec3dd6abbd77b38d71810725956bbce04e20d9282d5563208c86ab6ff9864f18986e462f0b8836;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he626b40f936ef813cf430bd7e232a33d4818b2c89066e4e5970e8653b731bce35254530d34fa108cb2aa9b9dec48bd57055256499dc9de1c0bec7715adc1970b5f097773289b3853f1f17262cc68b6317b54fcf43b74a1fbdf8c8e02ddcbdeb283aec24db406bc127658d46c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9c97984a294862c01e792f67cf6361df945440c04c082d0b7af7a131bf0a4b0867078398b3034e237feed5f9058b8e317757c4a061531abf58f3f0130e7c1e499597c48cdb603f138c9f490ece22fd54385eb6c2ba0a7e79fb78cde9dafbcfd7003ea8dbd8fd3c06767fd1c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h278e37bbd0d201366e1551376ccc83a4fdddf4c05ffc6f979a9c3f25476003cc638677b563abf7d218c9e6946e6f4b5379f651c56e8fb9133ead2ab6a096f9d2540f8c4bd762a7f1d458992654c281472d857cf04f75f911ff889b593df7fb7ad55b1ef337a26fae8306bf56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha35b32a06374cb8d098770cfe410e5215ba9fc24cee9388f4fb56714888e2022af86b65d4b30a8633c5502b9e74830e055c7935b5e018159d50a7d09ef81f1cfcac8fd6c7520a50b44cd30450d5332c93144238573d73d70f5908dd561880a0f733ffe828c6974f3e564d34d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he031ef0be5ca540275271995ee2c005422b595dbcb2d2223bc3b2f657f7085d0c009e5a6e9fce39f5c9c07a25d58c3ad23bedc40cec6a0ef74a75ea67ad67fd91a2cff70876f0a570daf487a10a25da0211e4dc1be8a1aeb063e4904e2477373364bb5e8f050ec1e3663733c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf1c9c56aad92f40f77fb1330760afe7ef6d53365e134d5c236e32f64380f12babe75e5f4bb52f3ee0758e07293be95d72149c8e4c3fec9fef109ee0fcd5bfdef1070745d6e181992a2eeebd0c5c838eea417470d208cdddcfbb760c66f29544449125c889861e5ab5fdb0424;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7cac8e385d350a36def69de9cb5bfe4ec5580d836cc39d6064b2eedbb45ae05f79bdf3fa0c3142687f407edc7f3dc885fd59ae3b165c3d187868bb968cbdd31d30d07cb28b459542692d278c3d82720abbf2251e767fb072853adb86bafbaf0f766a67a1bf974fdebaeadb4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8d0b3867e7173f7dcd26a7bf6199c74a432e27358ccf3b5b304a0e4f5f8f73cddf463b8baa6221938cd57707db11e056efd30466a95e9d694631d2a763ce57bbb4e706157ae8cdb926a4ca9c2e4c483c1116e4c92955056b211209d1a0eeaaca7f14f4b6783cb3c6edeb2c04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc7e6d660f64ca4553e88a1fd5c6ac5f2b071e50977880da30eaf4b329b0a437f3f3965f37488afd1e38da3c125e918dae7434c04938561f005888438d63b5aae9b539e723b7b464c1420a58daab3eaaf1bdb81ac8d688a286ef482de8fb5869d89d8080c619cfff163b64008;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'heba4c09821be240eb4c12c1b3c9d2d463ab651b7bfadb19310d5d3f15d8edb3a204edb3d7f62f2b141eac7f572c115e5ee5034c7588bc8bb2429b8dfb833ed3b72d780bc9a8e231756abd34d01a8b4375da109910d4d64bac5b1c1db14c25ceb93a440fba1aa78832b757843;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1541a38a2facf19679badaa1f1379e2dc07817445979282fc82568f3e47c717ab37d61f88b7024a85e9ce357683691669d713283642ecca1cc076d3e38b61117bade3499e908b338d5b661f996b5b6d6db0b2784598a2e2d324020a2a002e1d621472626aadf7bc364f4f50e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3c3f0375669b66390bad1fb85f3e24001d451cad51a8b199f09961d2366649d8b7ae3481c819e72c7d5c476b878c81d01f160e7552cd7d096edd838b1f86132234366b2270e5002ed7f69fffc1efcd176cb7961986aaccd81a90608eec7ed94fce89a3e9df829bfc748ef9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha6e2ca5a29d5e9febc406f0c6c927c246d6e9fa37cd437cc7f8e5344dd04263a913f5e237bb5dd8d5c7e1799373b97c10569b74847f59b4eb988b95e38220ec25073e17b5b88adfbbdf8776a959da94f2cada0af8187c8434a47a3a5cc43a391fc8cb81354d493d8ac70452d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4a9c0edda51f8cdf54c80a462cd64c4e3ab30ffdb4c612316f3bd99ceb7001b1980515da02dcd626f065d8dbb1686a0effbf4be1bbd723dd3e0cd04670e4161a0bcc88beea0d1a2569d33bef8378f4455b1ff4d4f028c26b02c9fe2758ffc6924243beb77104a9853265b999;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5f72460f8ffb41f4d4190c8a2d964a8848f4e6afbc4b6b5093c383214bd5a24e596a51218009ba52c1e405136e2a36181e934b9fcf60f2a348daac7dde19e123b75db7af8f79c78c6082fe8334cf4b1e2cc480ccbd5b2508870b12a35e03ed35e79bf41dbef491264310eea9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h738c82463d4b9ddd517e657a824e97e6c17f5426ad5e2f0fe1598d5dc8a6fe7b401ed1e8ca16e586e80da292eba1cedead7c1bab1aed4fd843a8724ff8c3b132eced07e2571df4729646025e4600933e385f900314ce69ac8839939418852fa1e78c7ffaf864d22f4028d2c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9d314b94a9d9a6b9e5f5ea30a5d6b3a300f0ea8b36a0a147b8b37d7772fb0557249243e6e0b3728e8aa077e7379c565b2a816faabf2eacae1ea7f3090a76779ad7f2a18fb45b6098cfff5181ee81d372574c685389e2e9fe51b5dc8fb3d78c8909a49ffa1f0595546ebedf4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h67c70c4b3845140846d202882d189748bbed19f6111bc4ddfe9959e4d21cf34ef832719d018f65315de136c47c2e087cd29b3e7827d26cca0fd9e9f35421e5153b0438005bec847d577a3f123fee64921410786eea8ea5f24037e6ad62798966822504950e2d4b98dd9a9e08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1bfe224178fbba2dd4280fb88df6e5f5db3ca5dd227828966f67c0f170bfbf7404800d9c689820815dd12fe276d02f1ce52e5f00c7e134773806e53d89c9bd764eb73a22ae6973f7d8e975384175f1c244341c3f6e67318ffc0dc1e6b41ca0cd370ed8432995214edc6ece62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb40c18fe98cd3b1070a353303f7b59128dbe39a5543573c90e7772b9987610c40da0d538fb30fb369f59e02003f3c7164e5b8d90472aa7c8908b9c7d1e47ee7115fb75fc479e6aeef9a02fa8a22dd0226fbac67e9f8c331abd6ef69921017aa3b9f5ab37ff8e52aa68c062ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h36790d80c774a6cb63da01a65b73db67795dd0f4f9fd6bd54cd4db5d5a7d6c4b02c852a75f2b623b8e4df5c3707ad5013cdc8c9aef062d91791dd6a27065d8ed0eccf30b1a53e83d71bce8885bc3366bc12e2e7a4739a0f8be7a58f69dcf9b02e8d57ae9c6a553249b216190;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha5f732704a6c843d30e5d59d00a5be5cab261cf63662b3282b1a853d2ef7df3edf3e0f49ce19a8d275115fc980cffaaa31698f225dd4b8ff956257eaf863e028000a1741aafbc1d6b4afeddff5f92d63f8526fa34bd9d538a791ef6f035f4b9deb4456c59234b0f1402cbe47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2aaba6456528738fe65cc81dd4cfbcb417e5a39b6a3f0da4d3e95818a245975d92aa0cf5def3756c2d0faa04f2d8cd000be8c3f8420899c702545a89e8e5b02dc7455df270d8dcfd1c7dbe7fc1b11293fa14eefbc8548ec8c3714181133e5ee05526bf854761889a883a29b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb52633f18f9e6f6df31fc3306afb7c1cf77953a0a01f5962ff5c10821f883d28346c8e142579e8cb3fb60696cf09b584b6cf74382a4200377f87a889d967760b738cd5d89e595586d76e5e08ef6873f144faaea4b7b943462d21152e12ebf705e9a7d872d1f910572372634c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbb99212c9748dec0de873350c2607d8284c916d2bc30ac0d24705cdc789bb7401078261f912b061d8b3ce1dfb0f85fc8141c60f38afe357c41cdbc6b2ed4314b75883920781f642afadd07d23f1486877629808d32f96e962e35baa52a71e1c65803a324e76c2254270919b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha7f88af5ee84ff204c2927cb4550badbbcf4849cdadd2f719dda768d2d536cd0fa80310c10cc4615c76781fedf81ad08e793823dcb0efb3a4f0a982ed3e90813b7234a7af0cc9ef3c6295806935f303ab48dd66e44755a66234b4837b145ba0705bd0af2fb94dae2bc30da48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h112ef76ee9367b4ad2015cc19fccd4dd285531718edadd1e4f7222c73ba34f559dc9f1fa336aaffa56bd977d8eed18c416d9c7ed3a72841edb468e88d264621a36695bc837df7587d5baca6fdf0d577567d4ab6e0401287abb8e7886b68d6d23ccb77f963d85034a7533d0d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha783dee74bcef1da079b037e801331264d1525b6eb063dfdd9202205ad3d9c9300e3166cde6c4f0abd255693f665f826557bfddb729b334c6540f8d780afd2a9ecb7d83eb24d08c4e01ffa3c58a2a7b97bf5cd7b1a410ede8eb1424754de8ad3de09a81c10de11bc1263f03b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h52f60dd12b82645131dd9458e3b735cba886f4e78f8b59bfa3075eea6545f367b7bb26c204ffeaa80b11a6fd5dc159c6e3da0e69ad9b29af1d1828c2c3b043598c86134e187a412719373b3d27f7b1a09a74a255cdbff1497c119fa05fce671dbc314b412774e10ead52a67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb3585d3c2210dc0d709eced5683bd58ed36ac82bc846f33ebfb936498ddd7abf1cb7c47c75863e79d543a16db77d0b9af3722168237865a4a7269d35decb971687a794b5ee80878188382f91c5505c1605f814a602b734ef9f15350b8b5ae64bbde4cdc40687c1e476accdfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8236296e409bf8f9bc00fce963ac336e8776f7c927fb3a2263860333d4fbc74f532d902b23373b2310674196958947aaad55c45f4dbf63c4b09e1567945de9e33ebd77981fab8bc5131465830176936276a4d2fbe29c33a27d2e20788163db031c6bdcdb7cdd81d93b209d62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h59d4d660a7c3826602ff98f6fad25c74b707106441bda8d24636ea1b7277c6893523e118a199e5fa520f9b61ecf85871c3db4498cbee364bdbc9e23a2255c4fb864a8b991b26284712aa402f835a84a0eff927403510f35f3c35b5063898aa1ee5de95f5515e0abcc8ae6fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4989fd5644e814cbe0204eb901e87736866c625a3fb6924fb4c6d9036c20a4154f6fb86873a334ba130f860c4a6ee5b7ee5c7889087d8fbcea8708b9cb3383ce9dc962e2b01fbfe1a06faa20e9e06a2df4a91ccfef5d37e5cc8ad322ad6a509cbb992497be36af34a9ded874;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8ea37a8b7bac747732b903dbe2b4513ec1e07133a0909abc80081bea794e681e288eccdee445fb5472c0ac2bbe22801e6e11312ea18a854e43b7744d165510014ab6dc0365bf6d6a078354df4f86d1c996d9ec922272d2b8f0cea96933807bbaf6ac0dfeed1279493bc9e8a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'heb39f6587abe3814749205e9cd0ea274d6b06d0082f3f15c6b8743b55a34d43681d96705b95af905fca2fd84602b47f9b03072b0edb326de98b173130258ef3582605799d922ee8162d624ca196816c49b6c1c9abed6627f8e98a0ed3a67db2828b8e59020639d10892f7342;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc0830b3aa6d0319824645bac46ca605c8f685eacd817a6be13b0f091764a345a8aa2d997ea8533086748f7e60f1477359609fbfd3c104359e98816319b76e76d44035656b65a4568023cb8eb7128841009b74eed982fdb1f5eecae0b1b396af5d9deaff73dbff24f5a8db716;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4cb4a87c4e9b3c3b97386a8c7a4ad4a9ce94b09cd55eaf4f14cb2a82addea71a91fc0ddd63f33846defcfbf34a88a3c4abc4791aa1db6a3ed4544d2470082546f4def4fddfbfeb0c7c4e43bddcef89c334cff6d59dada098f056451cb13d131e7014ef93e144192b5f1918f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h349a64693fb4cb757e778c2c1b45443f82319a1a2dbc16f0613fd30858be069a77085ba0cdf5898bcb5488adca6a70484e77fbca85fa3d47fd9710c0806883eb1f6805960c5bb8b74b7ebd120e04cc86694341aab33eeafb10965723da4c29f4eac31238fadb7a05802662bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf305bdef353b220f923cabc86b1d83923f1bdc85405cda50b8d3834c57d52088eb5a7ba810f7eef96e206696e9d47f59dbdb0576ec7159a6db34dc1723f0a6ff87310ac7b1ef096e995f43f362eb804b53f82eb7562433ec92530dc5707285624bea4d3366b29e0e0d3223ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8e5923e3550fccca09e4bf806ee3faafc89d23a2cc54c91546a5f2225f107f8a197d10627a0d0ef79c4ccb5a919451416097d174bca293d9ac4467c144b2999fe11ca0901c906afbbe7362b69045c7b4976871e7a9821d895adf787f7622df741b84e78e7471e1829b5ecb3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf24f29c0b5ca2f4364aaeeec64be4beef64c229518ee1c08ed6b3f57e7223d638e46b633c94685ba7fa80604295994b2292060041138f918b6141f47cd03a030ade1831acb9ee08f073212171f14a133a058c385be157193597743ad218053412ad9dda8b763a2ce84be5d07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbb11ed5285fce2e70511ced0a9dfe29961713653356d926a50195e8125657722ed7c736b88bafe6b9fa913f21eb8e9d9b7f27299591ea1615924400bd32a05ca3640012f0cbf519ef9d8bdaed47d31bd724f9841a1f1dbe87978369172dd9dc5364630e8a6615970c5e91a7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf594baf34c2886a5764935336362e5d1efc57f69ccd0c25321da0215c90e11d264dc55d60d667ad5cedcc059c5447fd7f22ebb25a0dbcc1a5f06c8a21937dad950cc8710dee4d1e3389cebad46c1b6aad40626eb440779fce8c314878f32e1ca28a823ebb09ff54e485134de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h51366d88b919e127adc1fe52df991a283588214c0025c95436d762dd90d7508dc1302bca40f948ee159fa9e09d9c54d0aa0cab2a521172e39f65dd7c1e16b9f125c8bd2bfcd6dc18a67059c7a144cb26bb650c34ce8ce512fcbf8c6b7a2a0fc88d8438768803f00c8ff40b8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9c987f8168967b1de3edf2aaa3d0a53dc3ec061b673431bacfb74ed96b444c26874e50fd0fb0277704f9b263788f3ef7bc70d57883be251f5b1ca0bdfb26e6763788c439228c1b13278a82fb44bf83b7b2b4374f0f1398aa31c0638472521960078c21b2c5a6f62a1eb6c792;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6ffe2f14f9c94ab55017686a227419611941e84dab133c8a3fbcc0810fce179ad4667f256717013845515f4745fb421b6b355d2e180c81f345f7f811bdce830baf94de773425624c0f317aaa550dcb6953007bcb8b1f7ea9826afb44950eb221facb6b323a457202c0e86fab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h36e38f3951b78ba3c86e8cbd62e2fcc71bbaa49a09863dbbde502b63d071cf3e12b8a97b249b6ad45c349adec0d24709cae382760df5ffb24d8d90e5dfe2a99c940a88d6df18e57c5aaafa3d18be00b5e47cc184ea550c21a9d38fe88cf6f09d40799ddf1a67de7d0a292b15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he81addd6c6ebd109987c69bacdc1bb4ca1ef4042ca18716c6acb2e8db914b609177efefd5772a45d56b3e80e9839b7d47b3d1aa608de66ecdeeb188ceec8017941b6ca7f7c095dba4cb1ba48198e3a60f3fd31fddde4200dcfa3926285962fee326853c492279c6b3b2b42cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd61b12705df788851f3993642ff201ee28695dde904bf1406a5a5a609e4a51de1b1fbef8c34a0b9a9c2401010c4f67f76e58f51ca5b3b18dd31eb84e4abc103bbe3f56ffdd64e5b9b1622e427d129be9b7f60625e622d2322a8267e322ea5e72cf34cdc2575b988de15ffb58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h963e085ef5e4932ca08d2881ff0cdd868115d46fa0f15950823f73bcfcddf6d5be7f698db6f82f9afeac55ec8c69cf70af3c3c71410ff53c039291e40cafafd542c246dedcd6afd9a2082bbe1a1445eeba16e1484a05e8a21e82455188582a4a97c02b56e171986e95970d51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he50c1c0d19a7ae1da03984a0726a6a12b3bfe6a0e16dfc99ef7e2d383786a1b260218691e43e20c1224f7c7e1a737ea71b165e32df3b0415f6901c02908c607dd3310339dd723112ea48c9865ff3cc5a9b315ed1dafac8fc1d79ccf049e518acad536cff3474ed58421e0489;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9fa0072eb73096fa8a7a94109a90fc88c5e91a287bac2305c04ab446ead1f2f0a722c652b1b3e2f80c25dee4a1317d1d722669cc0788b46ac92afc743143362ea0d849f9b243bf7f07148dc32819b2f0598cc6aee3f2d0064fc716af231455e847967d6fa3b8a13ff730b39b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc29bde4cb949ae77f77ad478dff75e7d3151d44d6cac4791e1efa5eb6ed96acd48f7f0b88f715fa37282915b37f0d357bfaa0a3cbd78b383aada87ce0dbd390079745d17e8fab9e38203943f4a815461ecd8ad38ae3e22d76b0db6d420a2c2ba6e1ddb66c2e2bfa1208746eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h57645bd9adbaebda70bc3b04fbcf3004d3851292670d50c016b8784a977498514579dcf48f5d3ea85240ad8f2e27b65ab48b01c9dd7bb359652d272120fdbec9a5e6652d50ab1f7fbff2a55a8974df2c3410ed43f4939c135a5e832d532887e1d3513023b98ee2e1738977bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h44994d80d8c048ee4db5995d2a8ad45842712c2bd7fa0e7a402c39506fee06524d522f30b11fc9522658346fc2ee89dea5f281390ac48d283199424c4bbd1552058fccbee1d4a418203a63c03774b51e37f605fe493270f41eea55c04883968b67a165494ba7ca7ed702d06c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6e120eb81cac6854a7980063e2c4027abc06493d0be14f98ba39bf261aa6188c7e2c1d93e0884c8c9257b085264ac96467764f8dd1c00e0525461bff2aae0d372705d88404d87fb9447e3dbca0dcf8164931fb995dece83b91d25bc14a1171d27ea2ed043e593823d3eefd2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8fbfa99d26b075eb3018463150ae2555bdb42e3593f4a24acb85e52f5b60dc9e372b67b7b2afec19a79d05abd9a9bade07e903909854102ebd07ede255533e581b153ffe949d42084b9add964a2c260ae113d53cfd5d190b93d6a461623bd1e8250579c412344e0489c2f86e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hff5598dab1cf638e48a540d1a02d5ca9caca0c31b28472d823e8389ad7663378c323e90118c487c19c03ed10d38f39513575b17bca601f141b69987953c6430a0f4832b4e2320fe3b059a02eaee0471235ac4b78cb1c811fe9f02f64cc794d34553dde4abd521a9598ee0dee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd91d726b79b3a42b8a40e086b0fb25f5fde964d8cb95d64afbf8c13bc7bfd4ff59eb0ebdd6bab6d19fd33c8e55363001f02d0107e4f6e17cacf364b1fdd562be5a7f12d1886b09f91c623bd1fcc652df9ce5a41ced9683a54b29f2a1b31e30c40ce8dc3ed60a27b906ecf463;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2225a440e926a2b4951626d134896bdc38bc48aa29cf0441607deea79c2745ca07222b63357773ffee492600b8866c9c899bf5c0f0d86ae72a83535a13dba2ab16c98c75cf021ee832b2f151cd82cf2d360575d7b7c71d875fa7bcc628d794775496dbd9a3aa787abefe3898;
        #1
        $finish();
    end
endmodule
