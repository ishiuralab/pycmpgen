module testbench();
    reg [20:0] src0;
    reg [20:0] src1;
    reg [20:0] src2;
    reg [20:0] src3;
    reg [20:0] src4;
    reg [20:0] src5;
    reg [20:0] src6;
    reg [20:0] src7;
    reg [20:0] src8;
    reg [20:0] src9;
    reg [20:0] src10;
    reg [20:0] src11;
    reg [20:0] src12;
    reg [20:0] src13;
    reg [20:0] src14;
    reg [20:0] src15;
    reg [20:0] src16;
    reg [20:0] src17;
    reg [20:0] src18;
    reg [20:0] src19;
    reg [20:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd71502fdbcd1ee67a9d115dcf10cb022f17e679de9c43b37ad0b13a3981de8c616e65e7ec46273fc9ea92b86ada353caba347c5d587da1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d74ab72fc5c2e3b716d51bd9aef11afec98dcc65ae6c54af953faac499e99e90dc4f598e02a9ff11c294b59f17b8b318f3e7f63c16e65c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf7a767dc767833b604cf5faba7865bed8468f8254b5ad3f708a8451e749111f698bf5bb70b9d3e691195c28c58ab52c6e4fb4fbccdfe8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f3e16608e37a4bbd0da79a64a0769ae7876e11e2f735258faef3b809cf947618c0ba90f1bf17855fd8315ce425a5948c9b8b65fa073d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h878159fcc6a8ff766cfcb018ff8d299979a38d232110a406cf0d48ed5562f78cb4a19ef0f704124ac945382d0992e4ebb94a2b6a12e6c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129396a40f0d229b7b0e8fb8575adc23da7c503dcb597bcca448aa8a3bd350519c2628babaad5577caedcace62bf9c7b714fb0b907b444;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192eebb4c79bcb668a790a88247c5954ffb267c9cb6f87549c101f044d9a2377c205125fccc72e8b7342d0323a49646b8081fc70041b25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19213743f32e91f51a4a6a0963645afa4160e948b830de218659eefe48b40f32f5bdff5018b6de13d3012603b78637664947334a1a846c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5e8aabd60d50dbaa69e3af8305ab216ed0c44a1c1140380f1ca2ea287cf17c470aa298eb6b7935314ae3876d82ac1852c8b62175e1800;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4192e6e378e32edd123bc6a65589372911967b4fb293db66be0a4ef35e8e28774eb42038caa2ff5983209fac6d9ce03d6d184e4716512;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef96ec7b89bb227c0d4c77a18ef5847a17c345272e92844cab1ff2806127797105582d2e59e516a8d390f938f846cb6921cbc1dca3486f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb0e45c7ccc640799fd22178f2181db778f56487d64e9ff08a2d47a98bfa0c2bf22f99d5f402953ea11787a838292b15228a2d11ed7fd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17331dff9193319a5de53a2119b4e0a59e58da5565cb05347b578a6942b05f0c727285c1e627ef43f7c13d196abc3b75522f44041b61b49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114dc01519c3047c1226913590d6e13b265f6482728b7c59479603f6648f0c2390ae760f1eeb76770957bc110d1820540586f1799b6b78a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b99a7fe7cc968efee412e77115c4dcf81639c4a9f57cd8afdf95c57c0376b3fdce0f2336f338865cd22fdbae544de0c5c7988c3dcc27d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9ddb77914bb1eb4a99f06c6bed6ee43dbd2477b4037fad1547a0fe20d96111c442e3bdbf8105125ebe5073fe484df80bf88a9dbb5a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cef3a617f52b32c8bf62d119a4d5567dc5ffc67344f57a9d3078a9d11d7089e06ca3427176b7ae84fac21c7043b8e03b03b7997872b3ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab0b045d7b0b75af34e108bc306647a90eb3bb90274dc683064a3603860deb0d787b9a59521b3fd455c26236105306865e31fe0732f38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he045a4e99d4ddcc3b4c194edc60056066f0c40ce1111581b995d7c80d99aca5664f48e3fa2be2261a41bdd01e398252e04f749bd9ae322;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b3f0b438cd702edaac8a425fc0b4c3a88a5099bcb40eda33b02939851734b2e230f388566ae01f66deb26f16fd244136689872c46cdeb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7ed0fabc9c62adb1af18bb7d34f1555a0ff2234df85c095fb77e4c6ce262863b473a1245660789e1a16aa26d8f2db5d41053b14d89155;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24a5585622728e7ee5ba8bb1b7a637616f420caac27502f494f503ecd548cc8d78a384f08ebb8ddacf71036ee5e40ac33e75f3ca36b646;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34f844b9b1040dd4cff984ad1137c2f609c997f2f5a5d1fff12d055e6c1e57985bd21c7b7b99f9186fdb7c9f6506b98787ad905a30cadb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a421ab087ffa7dd6c0b0ffef784f59aa8982affbfa1b20a8c5bd86860b628d4cbd839ce8849400ed5160d4bfd3c06d106b4c679f0b051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed3e9b1b58b030e8d6fcc56c86d26bf9b3904e80b3496b58439de063b70f9cd5c6fafe9f7dc731fa12e61f12211e89ff36ec42cc5bbf84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2763887875cd8e79eedb94eff8126b2bfaee51211b41120043f3a84e9b09288280a70eec51893493cb77d95a125bf2519af70e22e0f7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1d0ccd94e0b0c073c7d2db73ceac8a970a2ad819feee9e77118abfceea2033be714cd5cd0f0cb35ce39c72bc38434bf0b3401e0a6c924;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae097e7f3dcdc7d5d450ebf1caafe3154dfcfd1e83abd1a1b5cf5c052019d785c74f56ba8f1a6c2c8ac92d29a7c2d474c5293f5e8ce987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2752d3b1599eecb24119a748ae1300ffd4d2d6708ce24666a7543850219034a4e3de7cc8b8bbc74d9ea04e0da03d201ab22c2aa84cdaf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a67d1a2c15ab8b14144b17067af0352ea98dd8216557b897450d0f70eeac439cf6abaea8eb24cee5dca4e310c1884396abd1fc3239600a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb78e74277a76c78263b1ebe6e9b4579034d2a7811485e5db55c1d52e1e8482f10534a0c1173cddd56503f8cdb26ee5e162a7d59744f00b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbeafef97522a994c772ce93b4ad11527bc1d15606737975e584fe0fc70f6413bba0013f4f6abced8b7b18e912878142f490f41edf62b9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a1939313743d70fdfc2d72af4e50269dd823a3abe1ce7c4769b618b56bcf7ed623fc6f70661a62c8a02c4febe65e559bc5700baf3d386;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h864e9c23f2486783b1b331a0008de41be81ccfa464102bf27a016b4131c0cd8d16c46fe16b5371c4b5e8b99f0bcd2bc60274dc649c914b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ad7dcd8d0279766d8b95b3fb113a77307faeb1e09ca2de479e20b56d7df1be8ab5c21c194c468c51f55bae299641172c4d7c6620ddee0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9541ad66b757fa751f7e0aeaa353f98dca69a35cc4d469a7a444f8172a997db5baf43955a87f1493a4510d0decfaeee194801665607a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4b186ddb746c54eef9fe2677cc454a6cdfe153b9733c4a233be7df72d58abdce4882db3deec431e0f1bdd65acbf6e3847b7035d5bb88c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194124507029b718acf18e45db03035d889855d0fdfbfe05024832696d92db424d8f4fcb6c063814854750347a925e5a99b6a042c0b5221;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b91a2ffd16730cde6c04c165745e2552f17f890a6d226ca1a90d42608590cc931001e93837ec92796e64b1032163a0a7f6ec3f44210285;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cc1c0b416f787307ffab23324216d4ad2b2e6bf44d9da76110ea8449ebfacb8419730313e41289227dde38a4ac56a4359bd11aeed0c5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a723d99b3caac26350fecabb3aebc35d29d65881eac690e7fc918cbfbabcfd49968a90e81c31c66c7e619d0b8c08ef5b8940d65a680f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf3e98027f7fdc9848adbd5bfb8f40f6bc5310e0bb3d8f81bc2efba42c6092ceeda761913259938ad3b4786739c1cef7dc70986025b482;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1222c18f868b9bf92bc58eb3b9e1989d7c2d4e372eac7b2ffb3dc3a2a70f4de3683ef429e69887a47e745ee5b6fbaad2c0b594f1406a62f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189e03228bc7906d66c41d304c46ccbfff15bc101d2e72556fca38c22dce20604dd16cdae201467cefed187c084ee0b18c137f24cf30445;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194d11983c53c3913d3768388f8ed3f3270ebd3351aca1b5f5d92c8fec4f4972d7296e9d5c4514d1cf9853dbbb12a80f24c934f0a211e08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e76e4c69f3d8f3b5f0f6aad86e26c9b411ba05fe8f8c25fbca643bf46cb5a05d9ce9642412a9af801ebf646ff7855c616295c309326306;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13de115dcf51cd90654e094c5f0eecd0f2bc7ad7531d557c546b5df4f1147444d278f4e5c9a7fd1837f056b3aba8cb247531ed3c08c4a01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1831d06833141b32637edca6f61f005dd4cae648832e5a45f71ed82cf0b579079f2d42303da861faacad8907a08f1bb897e9478666c7abc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6cdc45fe1f64e82efbda4f9e660a91fda4d21d14ee1932f9d9cec139dc3e8fc34ead2a29f8cbc7b52850d7a6c549118c82b99bf63faa3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3f4c085ae01231eee0ac6a14b0c24a67ba43e60b1a964c15bb1be4d08632b760728a52e6bd9f2318933c1cace8ff56742addf707733a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19613e7919fef1bc4bdfb3f3ca29da8fa5a0e122d1f972171f6386f0466b7ca2e93b8d1ee74c9c768354ab2979b0742916b32ea07d85b40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde6d22c4031425e91db4417e8784bb0bff77315051ce009ad0f8303d75c9eaf40a8fb1377b23eac38a22c0c10056d4bd801640e17a535c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28c00e5955f8088704abe96633580d3b2f46cf15c591701818d826743dc2a9f4c1784238840b2334f876d124bde5c9c880a71b8b29e3f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a03a0b7440b6564879143f89276940d55c6545d75ef0c7c17b7a8b9cb4a92d17c1fa8bfbce97636eba7df3f51ef6eb2e6ff2d8c28a9d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0d5edabf212d90e14597b3a28d5c12d9a58c4f35413074fe649390611f50bf5d1f99a49a93bd8b5ccf4971ff1de50c2c0c3e1efde2749;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h747ef301f61e8ab0393df8a55db7dd9b81f25995d84fcde4d5715dec8cc7717e9b37287d1f7033b243426eea1076dd44aaf76066ab590;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a8054a0934b90ee8f2c6e1632988d7e8b36c0d946ee1bbf804aac0007651e1ceb0f50f02cb04378185671f5cd0757780b787da7910c74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b6077bd38cbd6c77a8ee37714cd6d96a7f15d5d16a79db5e4afc259ea300a33c78e13deee3d459bd8e407eaf6e058475849c7e455e8dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff0b45448334d987244518e7f8b772889fef4430f4ad1d2d429dd9149bddbbba10e35beae630abb94bb7d8137c78044874d43b67ab239b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c025b619aa692e9a33b1c260878843fe055e3d10c72e8bc39768f5d83b9b7ddcfbfcaaa4cef7e41c9afd4de74973cf73599780a4ca5ba0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b886dd73715f4b3fa216a31a3b3db6479ab2dcc7e82e652eb7698850952421859ef6d8cde91298dcdcc4897b4e2c6315adfa36288419c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab25e3e8b30f1e70df3b730926e07936a10b1dc5bb250e638c0ada8aeb549232c284a34ba0d9b7a9fcd1105c86cf0b96a5e74317aa9bed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82f31051e40a54bd840921c9ff3990a9d920181961951e1a73045490d5d581830940bb3c5d646aacb8662779dac99b0f347baea3214c88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb244493446f80571894e6187c7e151ab7fbbdb6c115e4dfbe160839a6967ad5d06aa0ed13c27f577da794652e94f214c30d0696735ae0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfdb237194e158e19ae33b5a2c9cf7b099311d1fead175d898d7123e19ec0ca510bc418c9744c0da6a2eb39cb9bdba2dab3bcd5090cfde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3ded9397b7e917cb5261abba11d1ce8d5aae31ceca7bc5e4a35ab6789ad176f418d6e402345880c490db69c85530aca435df612965f1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d299913e91df05bf95e447b2877b2e34860cd5a66d0250850297943de625b159f7dc93c1a5d1c6f5b5d3a898d3bf0e594739f47015f27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b203b2228d32bd2d183918fe1e015b1b346c8c940800bcf30bc12cc50d00d159770cbc19f82fdd104fd60a0a0efa9957d2ce0b859354f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he65ac80f3b61e8cca7f3c49f9b9e374eea25fffa5502a6b2ec5c2c063429b17388d262a2e85c81ed51d6f2893f63b926c62ba0f1262f41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc17a9ac40d6877087a4eeb497937167992af5c20b58233bae985c011cef35f2f41deb37192e6ef8cb83104ae159a52da49ae657efbae87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haae69d0d9b7030a804794e9fbc53f22cc03307213ef7978776b28c2b14cf7fd3814061d3d96a99de28540cd3033ad9623e2faf4ce7497;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f422893fad41d068249332e35ff3ffc0608a54021b84eff5338f1828c55255be587987f26890fcc71beb5991842120cf1366ab42f12c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b26e2e7b6d888553d0d2cac25acaf0a62db7663402936e83fba1db10d19562f027cbd0b9d4570ea4976763e1992d234f6c84e3b46d3ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4009937a968593e35988beb74028c49db5945adb0eb13dcdad5ca5a347fff895759d021ebf47afdc9832969d6ba35a1f8075d5a115d2b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h637aba324c83110308edcda90549ab03d21a2ab3e373a0a0f1bed05a1c7b3293a79e43c218698af06496a52a54a158baf6dfbd3f0ddc72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a3652a824b4bd5f1617315cd13b0448871e9fc59eb9eb16919d21b4d56a5d1fa0784424f022d548c909628b0a5796f6861a9eb6071780;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1536e25ec47db5a51871b667f29dac632ba05dbe2bf994136f9ac2671b1b3fa859888302615a6e7d022e16358fa8afae6eb7ec5ca34fb08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c89b8ab33942c6a4bddd6316357df69856a344f1ee52b555a6ecc9a4216c72d2a68d78c76b8825c10f47663d9b4b8be8e99781fc885da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadb0e6fd3904f362381ae4256a2a3a0ab8351a23677b4a36bf8d26e19604b673bead10f3f51a3b753cb1f503c6be867f3e3d996d006932;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1414e09075714cf8b3b85b8b453413bd8fd2e748a915af68f4fb45086a18f15d388e49954f32b823c9f25b26f112c7979ebcb9310ee6c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92da263281e88c507297c07bd27c1aa48ca16c4401d16a821cfcf6eb6a7abaf302650c790228af58cdf9946ca7e58de75b6f3948ef3c1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3e0c4a858e86d88a96f810f0da318ad56fab22496a6ac4da357a4f41d5593d53edb40bcc20ed325d0593769e40cc0a605cef9c3aa6d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0d5306ff6af87b6372611a7ac37e0813e8a8797dc4096588bb4b2d97309c95cb59a36fa5bac839282eef772da8ac90a0275b9bd6c2c33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7ca35bc94d8db07454a8df3c96c77acfa6ce289ac1aae2413b71b0df8c2ce45c909176d4f54bccf50c6d429f7e898e6432e0ec520788f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162fc698847470f009400740812e5fcf2aa6c89768e69c4cc3b36faf55460daecbc0cf8a11c5b7a3df9b7c8a8c154380cf45cb8c3f60260;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0403627261c072fb59be4d717decb83f03d27b47c4ea22e609086b5ed6ab37fc183f2da20a26b5ad162e536df297433d97bba32d8a991;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144047b9419fe77e29edf66594c8056dc4c14da60dea7e875eb3818ebd5987a87e991522f039f7670cc96cce1c7e5de3640f563db1c6203;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha080d7199e6ed3293f51dbe27714a9ec0c8c2cc8069b39ff7ad63c0a4c5a2bccd0c07304c37efa144ca146c88a1063fce5a18c5f84ee0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbdd148f52b5960ec7ddf084573741d76150fca4556128bc6e262dfd8db574eb8accc8552418cb4174279d61752af33af62a864e8e65127;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120e4afb51df2286ac5d08581ce25aa690651e359382515490d8481bc1cda4ba141124b3d22d7cb0c0410f6004e3fee4068f9df3f21c304;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16602ad6c0236527b1538782cdf38d24f3fa4417f86893046104e7b1e5ee833b3f04ba6a9c526e1bb1e9bc2bfc713b2f9bd3538f3081abc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf820192b5214678d7956d96927d99903b1e3bb46c52bd90fe42234cea3455202c27ac8dafccdf57615d20f8ad733b48d899083efb1a2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b04aa5db921c0caace282a933c6934095f0d50a031bf17bf31e1840040126110db4c64c4bdc10e1cf26b7eab73860ae8625ca232a511b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee36d9997438d9cba713d9bc7389dfcb07794f61300038270beec232effba618b862e90e92f13a665ebaf4332061245e91098cf2315abf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bf31e2f29cde7cea16a0e2d849f3ac7aafab9e01404d4a9df42987ab838735557dde8a3cb437d5b80e7e67ae41bdfeb1e908ebee5e145;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e2d1aba5f3cd32b93a8f23f7b8f7bf6a47aa186007ab2d6baf2c443492d06b685d2b9c8783d98f78c52a999be06518a323a981a15565e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb795d54b2f1372286e83e46eacf3242bc17a05c764642ee94ef59eefd627f825b35bc63620e32a14b2cdc0b2d64615eb80b74ffd88cd9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3831d60667dc40be826792ec3fe61aa0968a7dca137b89f36b8eb983c56d0169ece98603944577d33932e78288c069efcefb6417419a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha77644f192724008a14a49980be0992d9792f6f640eb3408e3fab6bffdfa787919af83c4962db43a2fe8a9c659f701c5eab411637e14cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1faacea15ec5222a5803eafcd3fb429834026f523624aef4d99f8c7ce2d6d32444c0c88165ddbec8b21c21399175bd8782f384aae7bc5a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6af5a31c12f4415358aab6bfdb8c68cc6f420110c4ec24bf7fd5402a544291e7557af9b4eee8cae211a824939332eec56212a3c95c0da9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0b4f1cdb971d3e193cd5fad5d7b5860947ffd111f3657d06a77e5a430d68c0b86e7ffed8884ad93eee625d5d55bd710b58cba7fac52dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30dd3551412c3b4dcf3cc8667f00042e54190c976867dcfbfe400a5092ab4928a8f432f63dc369e4bd70d9f1c46b333757718bc4eac112;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175f23f84ca8a5a2f48c9341ed08092874d3a754783371296bfee4a1d511d2718bea78786c013d19345dfd4beaf5623b80db3153f70eace;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da8bc8f79f34c4901cfea2bb8ecd1b993ba49ec6c4a02b9bb1e02de54a83d15b26e5c1e287d01b8d570fc5a92cabaf414b0e14505fb77e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb789f357474b662f6f9f9807e7f91930e61c32abf6824bc546fa6ee3d5165af83b41e418da8fcaeb65a607f689a7606846deef49a49acc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16769a11c85ab2bd042dc3e53094aa9aa09862e5777f52d44193c5aa13e934afd902e8063164747f07781c70247c6671936e5cce2155727;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43426b2dea3fcff576b79d85606eaeb300663783c67e7bcd69691178dcbdfabf76d34b501058a4f752527a8195878d397b5e0341cbc72a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1342815abf298296256d7642bf4e691ff60dfcd39d886d9c09a553853228073de5fdad9bff7fa2dfee3a4bbd0f938bc1a80ce1b431ba256;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cff56e573509b4983f656fbca9ec37ec56d21b16ffd27deaee511fa7b702eabf1a5eb76f7b3e72cb5e2d897d38db66e1af331d1af4cb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114727b7c5aad87743a22e8ff4248cb68aa1636a584f785e8ae1319bb1abf7f23740253d068606930d99e5ce845d8568394cfffdf81f2ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1887242afc245a945570cdb09d7dd0074595fb3961acea4334bbd45300a7fe6de7f5c370a44d661de2a057deb797f2ba6fec30b7628566f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he32d2f27f0a616682b61a373d235aa87d4a89fb287588097a9639f0c6a0caba0ae72593d941d9e1f4e6fa618f734bbb5cb9e07f159a190;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1133b100e6e468244653a412e0482ec9b0dc7a374749ebd9610ad71418fcf18c7102baaf3805745b9e0c5cdcba001723cc1bf3d698d4eea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h214e193733f55faf8d026807c8b5320f7adbbb6ff71700aad168ab0cc715f0ae09b8dc1e00ee637481f6b1603dea03212cc0a0d9bc165a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186981ecb921413f7b3bb1ea9f3257e29d0f1b992dc5022eca8f9c53959ab143fa99408fb27686c8842857bf101cd858fa54874c2961d13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1bb45ac2fd2c159375debd7afaa64c8ac4b5a7df29874b5b899f795fcbf8c38f56bfdd97acb6d03c61739d83dbd441b35624ca4e7ca2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb518ce03e0736a7de667f95e1fa7a067a33cd732a4df396e4cb3932a178167ac7efeafa5fffcd825c55f365ebd64a03bb1e43173fe1b8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8727e133760b28da2f6ec957685a6770518558adf526b7f4f574e30fc0f6d65531898f2236da78f7d1be0892f910d350244fa3829fd62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112d9bb18217d823a55139d0826bc8a2ddbad1d9958deb0c3c59665f2baef2ffaca9ceb47bdd81780c1c3161bb83f71d527a5fb4f962c0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h704bdd7516561c20921fed7a7a751d1bf69566c0a70e84f195009b2596c159980af62b08c145e38c56425ce8b35da646f5893213406343;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a3dc77da7eebd478bc5d2b9291dab3e42509e01254a6fdf3b5d6cc48fb95fbc42a679d906c5caf4b2d6074c0d827f55ce8dac49d1c80f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8d3a653807c22fc0663e052f767d90869eea3dc1d171ce876a638a9eabc7af3b1bd91c9c245b570e7335132a42f1caf98bfdf0708e752;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74c35c3b652269b763362849070b63b70455f1515e69cf6d08e6c5d0608c7434a2c49061a8f50d171274cd08e7e72f8d88a7ea12aa5e24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f08add5f62630392005216ff95931033f406f0d050d493c6da5d7d425b63b9d98c03a9c649ab3c8d95a9845bfbb1bc0e3dea294b1f4da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8479f202e341bf25a949789c50ded27ece612dc35a8626eb4e376e1814cde7fe0a10a3aef1ff23bbf22dd5186f34c04d05392f43db845;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c00a7911b506bd4a31a52b60bfc19fea5437ef1fc9942b1cd5119c6a95a74926ec92bf5b607c8ba678074c1a147ccc872f85dbb6bb1980;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfd3a2849f8c548c4d62348671c102b96a18fb0ee7922e9a11bcbe7bc245e758074547a795e3192f71b83546429d441b665f2b261ca8f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb7099d512bb9198f5ccb0199b407123cdd6259fcf3e1b9b1ed3d9bea55e4b79fafb269f3d653b34a3d4a5a85bcd635362a745535921a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94c8023de9edbabf4b946265aa36f741c04f5a12b020d83cbfcbf360e509c2253cbba132b79e5be02d9fff64c1c28682816734f42af3fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbccb750718fa73080ef96e4a4d9fff3e96e5bf1fc11d0a6f2d79694ab08d15d4fad852225a708d1c1bdd6932864189f1fd0ba5201d750;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15686a858e7614931a73dc3b9517034ca6069afe508f6d7ac980bc060581b615b1e7bbf5d7bef8ec7116e4ad8725c7399152e702d0ac737;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189d59eb819f60a2d40b276e565de0f9cfe1fed7868ee1a01e1751f0520f0bec8519aa167a0784622ec344b96cadc5e5a91b130c37c33cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd88c6cc5171ed221b032aacfdda3543d08d225adb9e0a1832a33df8fb9c91e2b90424a763a926de60ee6b9a300317a3b9f0cc5bd0aeef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc11ead619a76ad7d33ae85f68f4d65665a885db31674f81ad5237a5680a89093641fd38b54509920c12daf7fbc7d7d47979bce4165f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habc4c8e898f6a0e6ff7467b4329079022eea27a6fb4e2b120c538ee8897aa9933c3f6b2b6f5574ade5b3400d87ef8dcb3777f219268070;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137daa58beec58fc613f893d54cc933d49f6b6a0c8730c096579d274ffdae8a4f7d35adb4b99ca6f0ced14406bdfb21d7bbd3025fdc4e33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14924d9c4ace985b6f90bf6f62d1422d170e6a48b42dd3f4083d7bc5bb43c913e40164e0cdb4babeb7a9f7dd4b02ef2aa76cab140db764;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195500f608287c01b0e9cdbfb39f9e72ef3edaf11e4a7f7a43ba064bd84f86b42946a3a062696a64de759b98882bc546be95f33657fe5cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ab1a96f755d50f70a3fec389c3e1812a78b3edf6279afc88e87b3f24be1b6fe342dc7426bcfd1773c207cb132b9361a2ea97ad8a35382;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h501607558db04af994e8d87923c05b794b3cb84c987d803e99e7a7fd07ce611bc81c956e1b4a7c4afb2ac046c582da9a5e3f7fff330de4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd61b218c86a02689c8685bc44eeb69d850ded5cde63e08847035b3c639030e5460d41e994985f31e9ebcb00a897fc1f0f94412063ca92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1068612814cd610f14cf872593c014f38c6edcdb1c5d412d7bcb8fcc7a440183f581379fc9bb7c45e26bb46414a0f941b93c973880388a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127444d671c6676a6786c6bb4af3ac24baf546cf305eae2a22cd564d39e1b2d2ff53a54a117a3fef96832ab00edad9d881103900782ef5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118ef868a9b9556ced4395116eca05cc1d618be2e5d744a24a8bc16ae36a74983b88b8cfc52825c1d132b81b959ce93efffb426cd42dd77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45b57d2e62c712fc01817e962be938886c8ed9948491b8b62d97c626bb1945df5aef541f3f359f951904b5740cc923e7b0a742a06c7cdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e40f7d538c03dd3f9c28e441cd2c4c9027377e2cb6bdcaeab1d6e2c6e1f004e01852a88d86c2456c834a8e64425910664f63210b89ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf97242fb2262acbf1859c5a5733aedbe3449c019752b9d003225a1184cbff67e841fe519b73bc12a8fc05057288a3b4fbbbe5bc9ca570;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199b9bd5e0a67a9f1c93e927f81599e8c243925f0e33496017a75eca9d634011a99b5b589d590760d40cb630838b31392ab27314f25fd34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf8a87695eb36ec29d9dcc8e1ede896ca4db7e3e141b4b18e199416a6a7c53d87c267d0003960ef0c33e2dbffcf0d33a4aba0ddf8e291b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5fa315bbc8ad37d31937fa1c946e8549e4590734f281039ea3e6572483ad1fb4e72759f3266315aa21ec29c87ca5cf6573ae6c7e2b511;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha314ae90273af0872284c357e01196f7418ade277c6cb4845102d5ded57e139916898255fd93fd6ffbd5591009efa712e427601ff30c45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b481f5478703a9bae4644e19ea43ba502ce1b55b1d6f5ec106c88f3469409ed94f6e25548a6d597534bb79457f89853c87aaaa5b6e6d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d17497d20ce46b3090ab872c87eae0781734e24e7a3dccb6f769440317f207b182880d71c1ffd32a002b8d6365186db35e23a9ea1526b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb21edc26f2ae552a4fce5639b9eb154b41ab9aa4382e9f07fc3e4e30d746f60ea6eecc6d494e935576f92d245b5d90b0a0c11fcb73b3ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6008f20603036356e4c23bd3e0a8cef30ea933fd4aed600b6d1f0dd6c12f5a8298800698c209db55e61312307774991277c3cc04ec12f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he17765ae8e728cdc9e621a6f7ccfb97a30a9fbb7cdc518d1d817d459300c5a7e7a28c4c7e1f173c9723c2c8c792937575e6e2dbd121c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6855324bb68b2ea7aa74b498c766f3da05f319d59204aa51ade51e013e778c303089ecf491232c9213761ba6bb0e0a04fc5213d01693cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1810324f4a2b86818f313a236b157f9a0b0cab1bd6edec05a64c890209d4808c94259d448f296c4ceed5ba244720cdba00b45b787339075;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165508234793ebd9970a6741e95b51704ade7892740763ab7ba56d89dde0bc8896187758b4f79dfc89b75508eb23efbe857679986538837;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef12e8a2010d49d418966915e6f115a34a63a3159d1921621dabbf19c09e472a3ad16fdc8c6e16e0be83b07d83f07e0dcaf786b8c06da9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124929437a8077788cc16b4ecd62c9086370e265dc7fd1b43efad7f91e10b0f9a273a089d4946717a5e45aa26081615c70a4d4448ad5e15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfa9c8c6db089136d86aa66610a74c898da02b1caff486d4de9cc61cc823ae2abe3deb47e082c3183644adc347f75db4d37857dbc61f22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bfc6e825077508d5627485458c43d17d85c5d8f2b97025882f277db5603a490d0c95c9beb91278f4644b116c1a01c020185682c8920fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a5a59d0e3bb91e02ea0b725b63c9a3987edfc05c0e4901a27ca646068d89d733c76f50a03de4cce2cefd59f5c86fc42d5d7d3f00b3809;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1231990cb035828c274f8514961938943c7bb74862d4054853db992cd3878df2011250b517a7c89f3e65a7b38719b8d130b6a22cc0953f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9c27e2f09dee16d6ad366468faa04e179464619992e539f2b94db1bf200714e06a234a2d7a1d14ce459203d7e3be901b3807aee0d044f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1f7f51c65f97842c7d9d802576b98834f3bf1d3aa964e8c628ada9df1cba4ab0a8eefe1c27d77282150ed0745d165de51c0987b5e1d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159f633627c3a63670e44fe13d59fc8f4d29d3571f9256cd1ccbf3f967b9fd5b7e924e2bef282a4799d7227026e733c66d78a6d5029f3ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58809ec05d4f3d2f5bf914cf5284db30e842952eeac840c610716bcbf47d09c5fc5e997f99ab5196fb52672d9e17eb7ae2fe51d5ed7bab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h260371b805559f631ce9d43665dd5523f3676b3fc26a4c42c20d0ce01ea8b2577b56bc88328ebf0b586485e7db64a9cacf18016f1c47cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150aa353d699222570ecaf06c4205814643f2c31fa6c111de0332d5c679637e81135ba3babfd7bf5c441c955daf4bb2dc4ef1dcee8fc2db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef5736253f7de67c95b9c9e11a7ccff12010067bf6f97109dac540e6618d859e9b26d8a5a97eb71ef8ff8ed7c18bb5759d8b4a09d2182f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1695da468e9d01fa65c08b935568218375e9aee4fbd657009b2d7d2e6d73d89bd76e915ed92aafb21fcf2290d087a1230a112cba89bb196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8602c7744186805233fa0bfcc1bcb543735f91e951fca92fa0ce2776d650e324d52052e02f21adebf32e2c9300fdb991a0970bfe53f21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7d91f780f92d04405ce502b552f986f4a1d9e31a4acfd29d05c66306f23771dc20f0517a94675ba076cf97bf8357f084c1ff7dc0d420d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca79b2b3e5e811a8a01952aeb8bd2b0dfc323dd5680f7d834791c63e2443f31a15746cafca83958e06d957f4001ddda8dbb70d8970aba1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac1445bbf70a64895aaade46096cb40c8d16c972bce00f962df56b00af19f6c2810314fd82d42f82f62b1e7601cb0f17525604ef28474d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b571a95e21cff7b59aab2b0b8e7277d543885ed7fe950af468cec1c3462f13f15205c5f58266f368c4943fc657fbac2ea825366e992663;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf82ae0030c28255493fdb36e12bf11c19dfb8b1ecf8f1667dcdcad4e8a4bee9b5b9cf7ee613607a3b19b1786e847ef5ccea4a2b1df275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h693f3df9d4715e466e098405551da3de48bce982a4f4bba4a9bf147574d288404ed57b847cec911018bee5770c207eb8cbe57c324ad3a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b61c908d4128a3afc169794e8277fe26fd1974c4c7cf401757b3f1f0fabef6af4477bc7acb9e88983a8b46e232d902c226d5bc0de6b8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83dd96e06f28edd263092c6a7ed1cbfeab38b44a8698ab7642882b09e651c644a0caf0839811f2dcdb308173b299d18c6b2fd5aff33b40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6b7bf01ec4d3c6b2804a1e4cd4b9598dea633b3a0c2614b78f89792f27537373806944564ed777a334198a31f99c07149139f083bbbf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c49b66bb27d5dbf0d09b1fb0e654933f9a276066fe3a7d29370c144eecca5a8c81dfac0c4b3bc501817621816fae572b341d209c9e107;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18777e3431bf4ade66acc3328e76ad1c52c336249d5e5857d9aa599b06278d668a2ed07dcdabccd05eccd53830f1369104a7cd4cbcc513a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4027e78a61b5a95b775893b122b5130203e174201c61060649a0dc6bb694eee59ec2df14ebfbb0e5234622d508ac8c5dac7e52ff25b83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c2705c895c736e8fd87452722146e7a06601a54e161f62c41509ad6e7ec6ffcc2ede7f25df21ac1a96c7d9799dcd36e09e4c64c8d8a94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h506c769222793b4505673b3dcbdd2d9d47f0b5c87d3d12ecfcd1592be799dbc61a0bd51ba98aec645fbc8c6f3a6086b73818044669fd5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1292b8d90881c386e5aa339d4c1c42ce94c87033339a0b67c63136ead1b7d55c08ea38efa829f26faa441e75d91f772e322c2260890708b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d929435bae4871441c928d1cab9070036c4213f18f999a8b11048cb3202e503553ad2155ae3653bd46d3abef106af87dc10bf4e3ef2d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8fe058275115760d78ebd2ba3e74f8f1937a66b200b80d0805d3695abb2cb5e67585537c5b6536af3351a8edb9bee935ac9bb8bdb28ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc00293590dd2641c843569c8b67570d709386b3b95957b980a7393d166c5b4b7a3e397c32cbe807706d3bed3d1c7793b14d3bf067245de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2a33dde080699498457ae6575033e751ba7317eb1e72510a86d00787fa7825ce519196d642dfc54d5b6c5a2c575bedf52bd5df44e8e83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120cec52a079e8389612afa02149e03d5ff3f826243cf203fc860c2ddaf1eba477dd5d22a92a75532b05a5615d69891ebeaed7cba0e7a5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h136e2e001d01b49703dbd78aee24f65621ef375fb2bef9f1b59068810e01e8d41b6426f35e6c8a87bad4e407fcc9e87d6c1cc91cf0fe7c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcce7fc0c0a1660d64fdc92aaae470ad4bb4f9fa4cceaebe21882dfb772eecf96ef5a8dff53de35f83185e159ee7d392388dd37d9674f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h806b25da9beecef2d80cefe40a4387a151f7330dfa3ce5e9a3cd65c26e590e740b46f0e39cdc523019c9b63344ac67a31aabe1568dbd06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6c7271b4252a148e4c959f7060b03646ed68abedf33457b438d73841ae16e380e18849e1cced17bd5795c4e73b1131589bae1e3963579;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha11ad8a6e5b64456f7055d940af4061518bf498eecdd2222a1e25a4552af591cd39eeca624d6d2b0e3ea923896a6d9b5214ad21e5e9426;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha77b3112b7caa96ebe4056b1d584277d859dcc47a7a3b35f513a093d89b986a522a04837d4dfbb92ad05172f605d7356c79a479ea3ba72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd60bfb831778bd59f15957a730c22c72fe804822eaf666c4146123d2837c55029ba4fdabb858f88a3121efbc285dfbf9c4d9f81b665466;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99ef702848f80c90eaa8e56d46005df613dda6c968f7ffe1a258e785a03ba4075c507518b5fb185b62f2b092bf32787c52e525e989d7f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b59f87fe41fa077316947926dd681a7b8b58b6b9f0efa8fc156e65e7dd9699c9b44f6c532914aea5160871720688c9feeac0a164777b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80533fec1c6004223340801fb2cf22c08735be628495f569d1aab72e271031d56e44b112786c6b532abe69c20f4a04be3b0797424b628a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f2b96a38c13e2f789c22a36461b772d2cc6c1e7f8fe96ff1f8b16c06c7b631b27e5353039e9a93c34fbefe0a637ad13e2baecbfdf22d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad679b1d56ac11738fbc73bf2d4152c0113e0d71512a78393cceab10156bea743b894625ed93df6982f0d508980b3fca37aad9f5739b17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7058dbaa9d06cbf433710bd2d3377b690c7bb058133dddf30482d0e36ed17e900d63eb6f892bf6dc43932d834e1aaca4620b66588ede8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144c6b0dce3d02138457d72e02d51795d9693333f5b5eb4a0297d4ed71514985497d0667ea1cdc994bbdb5b769afbe64494152687bd83a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcd3f14f06ead96b3e6a6d9617f1f9aadd410832b69c994f739d0ee7229750ff7a13804ab146332aa6011f2fec35523095615ccf43e251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103cc1c46d6e45a2fde403358cdd64b44ccfac595e2db45d699b10c5eb1f54d58855172f12c8961dfb6b87cad6af533421227f7589258e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c8c52f6d86ee6ec4ec4a78fcd336b79701223064b29091aec64d503033202c6d7b2cf7425df0c2b8e9648c4742194099a99991cfd22cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cfb4f7e587731f2de3b2638baa7b9ea5267a64b100a4aa5ac9a880c25f0e3699debf6ca7c0212b704f363424b59a966ba06d67254f43f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ca210befeea67e2c8c87b778c7706b43ffadb3de22a150d28718224a50b05fcc26adf2092c5b72650c2d09ac613899176d6905822bcf4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h597eb821901fc7ee376b299de922dc1464aad3b80dd344c0f66615dfff65e2fc605dda1dcccf9f877aac4d8b91fc8fb2ba6a8ce969c7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e591b5e79146429c76425530ed27fcd15be31b06fc591a4ba7545ee0bdaf6bad85c6b64bc155763254a1f37899f47bb368d13fe64ca94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a0f7154c7ab7bfb261349b42d9f3f63d1b5c43fbad663f8b1ba18f9bec5b86235aea144cc686f61bc8672fd04b59f333da48837a9e551;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h663016de0f7ff187e3e9c008a21cac1d3a2618a8d02c45dcf6edace079ec8211a5f4971d3f5ca9cbd7949ba5df628ba893c89cbabd8f21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b556423519aaeb7d519616560aaa685796b7571a572eb5b32b3883840bcc0d6a49e9dd3efe742a0dc7031c4acc2c1944811a0ab2897cb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1368afc233369f0b7584980f63e9d80b34d8785f66b5b8c0cc53460bd1c880ffba2a5a1b2d7aaecf214c923f851eb8eb4bfc66fa06477be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1500a8ff2378241ed83c22760c61db69c703ef2afdc52fe28a07af5273e245f6a47d2804e5a11550e7eb3f5799dce7c66008728ccc817c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fabd2b61389cc7149c4451ade2b5478292899bf68f685c6ccafb705f98f3bc5f2ec0d8757743f5d24b2030106979b1c0193cc0a4ef3e7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf390b4fbf84b935b4d5018a5d15c1d9151a93fccc3a5b94cd53beeb49459fb132e5b94ffde6359fb921ec641de703b3d378492b6ca9d48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5693da9f22e9d2e237652ec5c614c754a6def883d9edc6fc50931bf152b9e9c03d763dc8b3a14743a6cfd2d4bbf7a6fea30828a7185c96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe7872d6798cbd40f87293fae36259e312976b471002df601d0cb15856d7e7be3e238be19ffd6f667d65222a369ab2518b5c05d1960773;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15cfaf1b865cc8b6794c67396978889872d3453f01324ff89b10886152b26a5e644b43d3309c5f83fbd3e23d1d608ec76d46b0992e39efc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8a5fa2b2f4e63e5d9a6bcca6775c64be5982afae7d6cb765fe7bfaaa4bdca04c18d0dd77c5b81ff6d18182f2c743909fcb91b0c9f6d2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5555074a7ef00b4fb7ff4b18a1b9f90094df95f835d8f638bf502659436016a198bdd578022801b6d46bc3c7df45b3435bba4becbd60d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4556ef60bedd4b36b87433c7e876d76627335c82b212f8c7a0520eb1d51fbc088871c93b9c7582319b09975acea44c31af4490c80c760b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2d241ec2d9b16f5991aa4b61b7bb2a50392b0163dda4dcd6b00b750bcfe648fbd3e6c50e2234f9b7becc432107900dbb421f306dd7e0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f437acd58eb655345cc617828d84a6584f4ef76a6778907bd10357b09c5ea6b71a51cdb2e4506b2747b2754260a210d150e835455ddc2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54c991ab4f04072b9b012050dcce9a0a8ff3233190a78198f48765b658561d915144ddf20865c51c9a0bad8a4a27a4322a5b54acfb87bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h865e572a115834a9fc36bd524bfc02bcde6ff8ffc145d48831de98be90aad3fb0c5825d906c73eecfc8415a30c547ab7de4a7108967624;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1234fcec056031c0a08466bdffea80ff27f9f9e9e372c6707d641eaea0509b06af1f28270966630f0486f6fb210d2b4778fda090b9926d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195bc3f99b96ff6ba98f5c6db9e621a32d463e32a7d8b7d51722ed5a7f2880a73cbaf086e140099915422cb043fd7a887126ee9739aa67b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1632b23b99845bdc97d6a2500413b3183148d9c135b27bd722b3c0badab5604dcd721b4f0d54f04eb75345cbe58f56b330228ddc85d811c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c941739f59820153afb55dc68132d08a12cf569c4ef6f2763fb2152c289f03521175601988f0e09d6ea31173bd75f66a2b098af41ab3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eac23646a6f032cc1feb32bc05e26e5d0ee5558b2c2eac7a9a62e968f732b4c220f8e9719d08c49865d22c62dbf25200eec7ed26c71162;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ed5092f78a05f794312e30166fe5c5b7fc69eccf69cd12bf82b9e5cedb4a05855232aa38c1f616ed5cb171dfcfcc6aa96fcbe13e6c025;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b63231cf9bb5a04e14e9d095cd3b10c8318b6ed780fe7963302a142cf4c45dac8943288f5e59379c4ed15f75ec6cf50913f3bcc86299a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb137f0bbbf3944057d1615203c0a670b8d92baa67bf9c5eb2ed0d5fcd91abf9431b735ac8d8f5dfd7cecd74af75e7290575208ea513be1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd2f289a31c408fea2f31153b97a13112e0fc1e7df36b83306e58ca70e6b44e7cf37fb8909181fdbb9c65d7ea9888c4ea01e4bc4722c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cc13e25b75bdfe9a24ce63ba6f27a6a9e351c21b1cb7f0a557f9accf4a81763ba54dfc0d8eb3aaa4db77b2e7a26dbb9552bb8de9442d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1618dc5c8bb3a03bf67c19c192402bdffd4a0f08a1c6a120c2ac54ceee9439a356366474b44ea8c5b65edc504167ff6bde3cd2e58186352;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he363c23af17a0efb5719555462ff70ce235aa7aae275c01f21ec5d75defa1bf4a7adbc93b9f0e591d013092ad8ee66c0a217344c29a363;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f227f72a913b1a6007b5e7e25dddf289c0ea36b397c50dc78dc6967316272595f881ada0cb8cca0ce926b57606df5e68bb1b2743663bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58f9bfe89f1d1e75856aac18a1693fb8831f847e4ae63efe3ab6b5b8046634f998c5bb093baf96a42b71c8daa4abada06127fd0586fffc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf6629ac11be1896c385c9873441bd91aff206598868db00b717b272e140bd480a99fe07342b4486048f626730d4f633ec01542b6914fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3a373a0772aa39b7bc5ac092ed8f50f7a121cd76a69b3942c110a94c52dc8f35791bb7c83b50216cab1ed4045c540c07559a8db67fdda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1c22dbc2110deb539f08a1f0327efed543f081ff9e1e72189c87e41429a0672f2a1b567a5465ecdcec0feafa6d402d21c92e89da84a43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a680ddff450aa2645dbed27b5c7c2c6221584b468edd5c10274d51de9fed8a84dd056b3b69023962e4c5da672e422087e6307d489fb6cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a5e2e763768d0dea03159faf1c800e3127fe6ee50f9c913233a4df128cff86af64af58aea4bd7be1478dd4bb1d86f04bc24de6cf6d6bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h975d5292ecc1f5bd869b5d76dc178921786953c02a87b062430f92140b9f2656935d7617c2ea08433157076205b1a414c3706a0cab30ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1024aa5a3b51c1eff1d9aaf071e9d45854a34f3ee2539b7fa801630b422d2f8e79c2f1072a9b580586129bb19dfee060877301f74c48cc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1f29e013007cd7295a721cdd43854af702a6a045e5af4305a90ea739a044d493460a5c5fff6a92cf058636773100e73b535f1dc8316b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34ac75a117c8e33086228c237fab2e16595c21b8b26ff6518696b85add4ee6184ad528c818b2f0771098bbcf8aae376cabf9fda3643e73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bedb45c1fc8e7e8b241b35e9ed2e68afaa8299af22778f8caa2b592345460f83c357f241cbaf876296175ef306209b20ac384f723f760;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2f9654ef627bea51a2af597819cbc70b91e069937dad3b0a7fd317107484fc31e39e568783262a253a40a4f5c9c17ae0786f95756c002;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181a8153aa0bd881dc724aba28fecf0ff96f9b2806520c39ecada396b7453d006c53387b764f4722473c27357c96034c269e86d4d3a4ac2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91684da91986a04a7c52056d53980d05fa850359514b1b62c89ccc5c4c2ed5afc289822a439746641ab613f989f26bbd4563b6520a651e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14aa77aab2cf12cfb0008efa89dfd2ee76554da12f4ebf7c6f1a10267564048b558b8bde681cc9ca7bddd298afb7bd4ae67bd77644702d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f75525f2eae97264add27810e3de5263e75f3e9455031b0a8bfd3fb72b8f34a95195fe5fdc35382ab8140d27941138edaa872fc263987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70dbb94abbaab1dc72c6e57e94b0dd1d5d000d8c4a475c341db42b02b48755c144bff38605d09afd8aee8c2b279627cba4faefa5738b56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120d70bb7b81845dc54576b9cfe769401d68539d16445bd87bdd20555d18a9f7bcfa1db3e5d17bec8385255471b0c0616a9033573e8c95f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5462aade36f4bb468fdec6e863a2d5e2461c49c7e2db7c6ea5977ab7c7141ce02025497923dbaf8f06309d4423a1d60a429eb8f915a8b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce4a09f90d265b31bb4b874edeeb34b757014c891193791b79357f0b8dcc283d451415adae83cc9c32d9e1b65db019f3ba138c78c7505f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbb3e63856ed5267e39b3ab0ec01f89a636d63a1b9a4eb4d53d8aa04baf60e7c5c930193133697803f200f8abf6b182649cbd900ee705f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d03608154a5894aff8f28c774d56752de30ae8f48e59a09e7a78e142180ca2b860b5df3d1249887322af89faa794ed4c8c73e8653cf97e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad30614d9e467d33feeed589752362a8bb250b339875040e98e3ec51ef6599c20d995b5a0b350fc60db85e090ec7548cfd1b4d5f13a3a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he26c30629c8625f4554a14818625f22f53bde60d1b2a8d7b8b873dff08fb02e5d36768837e6077e8cdf1f58128d3dc1696657b18479cec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6879eba1c383bd12340e7c8cb07b73becc7ee08861b20797564b163c9e043ca0793c5d1c05ce75cd66815444dd33e926673c01117d926;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a410108d417d2baea62bddd9e6f71fda286b03e92b3f306705377ccd83d71e7d7b23c9942f8d44e646ae8783114edc9f3cd0e2bbc01a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15014e768a73bf71df871dd2a283ed74da5dc7406b32d0f633ab283608c77cbfe19123da21e07ae0611308b26d012cae2061909526809b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb87c339889c7b12b32a47d248c5c7c0eed8b18f291716e361d901d56ca212cd693057c523528c497f781a066564de161902f11de638a5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3a4aabe2f999795ba0b0792ac73b4755c30bc034f5277a2d095a032b0423f97b58f1782bb2b4324898ded5d2aa08e1757077014cb1858;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde8471337935b090a980e431adc9ecbf69ccaa40fdc4efc123049d137d42785ee39769507f9e72162b37f0ec83fabc476f32037e08b51d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcf30bbb9f5defbb56e5f82159c777d7d0ba7554c6f46dba3edde26d6c95db97cad705da26c877a97c4ff8347394b3a38c406d0f798cee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df46177cde4b8265f33d946566341ed2cd0a3c52a5d1d8a56525d720b8425a1baac319315b199c06b8683fbeabfaef99ed025b6a228c95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1349e60e35d99b6cbcb79f3a020dcfbdade54e7aba8d99570f4b9c886cb36012a493d1d3ae8988515bda379c9c11ba874d95cbf564712dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea2674654322abd872ce97dddf6afcc3f2579f94bb367b304fddd818ed44a8ec325ad2223d2e6921dfef9bb6c8e2f889216ee87ac06afc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5ec5859ab6e9db65fc8ef5e776031b41fd77ae413ed7707f71e61fa49764892e6334d62c19307700c195c63c05976d47a61f177d5cd61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1df6d1fd34c38732f1baaad0c26a121e375b1e2f3944a5d2e4e145f00a1c84f954ca43b95ae1e2307721a5044f27695ab45ddd975cdc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3dbcece868712a57472c70fb9887c85938d5edb8fc3ec2e52ea1b164a304519af265fb16e83b87abbc46d696fa32245fd431629b3d96e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b28f8617b6fa49c69197a36774cd29d17c81c7ef2ea96aa17760cfea80142e99cb3ede330663229721e81e910a84b793f93cc2716930e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h812bfcd03618ae91634015930c9413b75837150632851affd9489ecbc6adc41de8562e364aa33c37a88115771f3a15e879d9d283af1c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65f86ff8edcffb7a4e48af59a816bcedb8cdf023ff70e0c69808db94d89f7353dd30e218baeed6b670735117005c9c35479b21c9d4694e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbfb0205b612d01dc19e92cca3e49b7e4e2d2e978cc013752223caff8baea449176f07d6e0ab5d26b55d6571ba750d93e0f7519460ceac5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b62d356e8e064df621c3bef8475e334db595b7ea60ff619f3fac19a068795db22c9a11eb3afda6976265627f41d284c4fcb4d9f4ecb6c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79a0db45d40dc53de047349ff2dea74b903df1bfc25e6b9d6e665cfdcdcb84d0a7bccd9be72df202024f0765d6f4fc4b91aeb6dc9173d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180d36f72bc804ac35993ed45e8ca6d588d414294d927cdd3d3bba26c8d9a8933d79efab8449905417d18921b8ab80f378db28a60d394ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb862aa1945c6d73efc000658b4754750ea23aea6f92060cd442835cafc9260b73ff3b0fdedc8dc6f68fe2f9be598041f045089ba80c05c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b608da7c451be3e1d0764f7ea70e3cec3fb6aa0788ea5ad7634bc4f5b0470e60a1da64aa599c854e7ad7724f2ced83c07e95c09ce130c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126080a945814dee8b67cd31f79086cb10b83a37cbfc916e6948a7a72dd46d8c3bf344da269e99c08b37a6933911bca253b2bf5a91a464;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1bc4e33c9d3f1edf557bc4a3578a0954e686f22046618a92ee1a6eda2b3b7d25c47f43e99d6101db1f55d21a1737fb27265d6800c8842;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a5ad4b06d0c5a075f0f980ba86fe3d0e290f0278b248bc0997d382075a92a76fd1908697362922c4aaa3be00b248e2b38fdd740015953;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17aafe8e8378dbd33a8a5d73d6f642d1ce943d367cccdf69b426c757d102f9206819c8ccdabf5d874deabf14b9da16c67f04e94cace1e99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5b28801631de7da200bff35700569784637df119a1ff2e655171438f7d84e3b9a0402010d317bf6473b4d1586bdc394c21a2cfb07df7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f4a7af725e7b2604d4b6951f5866a0851a258c6e6d55865c3964ed209bc7a9a64e8bf09802fdd74a35243f1dcd357cb4b7206d2b3209f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7855e1128cea3e7ab3e2665e9353465129ff4a89d3a5983bce1cdbac7e2307242acd7447a50ee63b639025c3806c688e55ab16cbd8538f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac2ccf03180167440607bf0ade44ce4f71464e66bb7521e8d5fd6c75b1ad4baf0ffdf9fbf73f658a34045cdcc21f1113ccbcc69ca39c37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109c7cd8aa18cd3d73d79e37f1537823be63ab6577357be8c692887ea9d4d9efb43f6ce1bd7fd6fa75fd56a5d4ff8fff8a7750526d03398;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18220d40055b0c284dbe1401042f7d25b6cf8309ec62ed3cee14f00961ede44239e0308d4f16febaae4871cb0d85f4da2cee1481b91a870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3a656cdc2b6c0bfcab84e69d29fc25f64dfda3ff8ea79331ba339ac08e105827ce7be9712159b226608737e05627a59383ec5eb14ab5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102aa92cfe8581616a1fba6624f9688552df10205114d10194912a6eb56819ea537faaa4a824b635640db68d2f4e5ec336376f2096384c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122e2bcddb09e8cf39bb33407fd2c31f1e6eeb42b98a6f7f45050179ce4846bd15ec055fee993ddab913bcf513403a9588035fe563f0059;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ae89d7e272d9a73eb40e4718ef4e038997fb30dda78a4a34c232b25068d071dc02422192ebc479931f9f72e017d024bc7fb0ea457080e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15741192186fe4fd81ce12e48bf404a53b4886d3fb2b893d0a0bd9eb63dbaecc633fddc93ce601aec9d084e510b39a23a4dba93ab7bbc64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c7919ad35e923f9dfb262075a08accec1f6c09f69d956dfb6d2ed94d416d2f26af03870402f2ab6ce88735f2f5520cf5a10dbcb7856c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dff5f956b5dae87224899a5c4dcf5ca1189dd0d4e0a20eb573babf813e5436c3349594fc4a5eb37d9118289c2e48fa733da681c2ae1d8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d4d5bb6a2af26fcc55f6f43787d923617c2561c8e249b799699b80e8f172463fd62a0e65e699b601d5d92330f4dc3e9a066756959222;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc7bd2ff82dd38ac680fe96dd6e20ab8b132ec5097c06e46cc843fea0c3bb68f34474011537f0ac218855f9274ee6750949aaf647de45d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62c173cc72b00a1f4fd3d017161dd074d2cd15aba27b3bb2352e7df2887e19543972423b8ab6996ce6c1b7a80d88b527bf44c8075d7697;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89ffc5879c4ebc0d6fd688caa4194524fb713911a7df3b9f9c4014296dad418cb7056de188776e98e37d80a23ed4ee114028a492bcf250;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4c785fa83d0b24c3b229e0a94fec510919584baac848620997b51cb6af60d17ef5033e06ec0b1a21f598d2161b3fe6227f99de59d249e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb45faa040b1d68f7187db9fee812cc199d5d887fb04975a1f0a85174bb1498bbf0376f10b662ebed9ac0241c27dba033b0ac7b9fe95c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4c4ae8c7d632a98414f9a0606669f00f9904269c269e331e50a7775bff5e11d2956eb58bb3d14ce12a10a217e5fe1c4f939cb678bba3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15185cff8f723fb47604f7887f480732226b3cf8851f9169be7b5cc6fa8569e3f81c54dde06cb3ab8dd479c3b6e93678da557179f21d898;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3174ebe2a159b3977dd9b7a08653205fa7b7d77367612374527ffea15502b3ad5cf9832f596b74e117bb04c94ffe76b2951249609c339;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f15b71f9a6f8a08184cb767d775d20b56bd1920c24b7b792560cbbab4ec12f78dad679047a9b0850e2b8d095e3033da0be16ea66961f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee7769b3865fe376909370574997a600ec10866a3f19c7a839acd968e8c4dede6bc74de58865f612a5ef1d2cf9c4527a6d9dfebe451840;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c1f80af9552c08d6d3c2368388c33e2dca1ae241b720e54153d26dff525a7da547be8f18311c29ebc871e69bc7e90b548d0461026cc81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdda4be941504384244108df3bf3db26fc0ccda154704097716f8c2e9dbfd32c1359f1ab4a5ddc22c2abf265673b54f17f3f3849760280;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f018d2a93b6e45c43373a6823f83a5a6a17c2bbbb216fe3a1d2b4ee9edc1a8b21e0d4d2c0ef5a71af0b1b12d500c2f017ec294a0aaeee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c683a5f58f2c8088a04de57d7be3559d21aa4bb4e24311e45d8c4f20d2d8390438b2cb92cc9a77b79ae4ba34757a853a9b1816dc7794;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13148f3bd4b230d8128a720095f37ea768ebbc939939ebb000492f0ec83b598b58f1958a354d842266008e80ba494427153384d9375dd1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3d1564ed09899058baadc5e8cd4d4c39fbbec36bfb95ce41910faec14cfad13cceb04e970cd4ca68466b83291150e9ef7c13d806665c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aad880eb91002ef7243b9ed04b9c9f18b0dacea28711516081ea05223f58ff5fb0e7153b6ac8ca3cbde34e55aa0da6a6e66e0c5d3fbf2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8cf749e44d4541770d65e285ef65e0cf5df2d926bc21bfeb7a1798ff211029564c698e0747d437aacfeb5a4371bbfd82270fbab551e495;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ce599bf4ea081dfbe98992186b4c69638e4ca084f493d6bfd4f1f6342b0a05084582fbb9cdd04d98d45795791430e59940c00de715f94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ff4d71dbeb22e1170f5211ec0c3d5aacb822e3d70e83c68668b5994fc49e8271205118b0f077a994a19d4fb8c202db00de2cde755b231;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h669ebf4be133ce533f2a12303ddec4890c77ab0150d3d31bc532653fe222ccd7f08b875f38d5b59294bbc1fb35e9337661d39035beae4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb61b932db410fa50b1fab7536dbb1afdb2ce3238de1033556629bec8bb5c27ba7acf838830f28fbd0d32a71cee8cc1e5d86825068e1f4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64082df9aa6705c1049c2e7fe1fefdebb43b23565d40f8aab63d5942ffbf226a37c64c0fac0e10715289605e2154b17c1c23ed4e374c99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he41161a3670fd361253bdefa701a0940eda32c5c84062e5697d493a2636a382dbae984017acb000e5a0f35237703cb192f42b8285a215;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h957497ef67acb2b8b1a8bdeea071f00fae8786a277e1f7a78e6509d1af082e08f184f45aa2e66e3e09091b56a45d41298cb43d89726e3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d51be6f3274858bf8945020b08fb5259d8df4275d06e853dbd12c2efb08171b055b86ca1afe47b00e24d546b66a9951edd7e184e0be229;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h221610ed1810fac13064e36c269edc13492e759012d6e20a0c5185ac03cb6dd6d198cb44e520bb11418cae55df9a4e8b7e51ad3cd08576;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cc4b056a9518df84af6166ecdec094dc5f5846e6412b566cde6340d23d58243d7ca93cdbd547f92d49f3886d455065704cce079c28034;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f765ad36e77950141affb1f439aef5af64418c48604f5a506d3fd9e77e44fb6a1e16eb52dd32e65f1c142a4607aea463438c6a4770171;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha430e586f95936f2c6ef30d1e664cd6ebb3346a785148b8c680c043adb6cac34f1acec69d5993f6d2d34e19d2422a9f62448011e5038d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he91edfd379f30db42b5750c034ecc40069868682dc166bc486977519babc475d075a7a890fe1f0d14ee64f17ea117cf7a9699ffe67d602;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbccb963802966c46d3568f1b4ae262a26436c08c310b9a80a58260a2002c96369f67cd6d9b57ddbd791ea1992d76fbb67917fd8e90c7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30687fa141ad319c0c86ed376e7bad58b9837160e274123215c735cbd164172de1dea726439599d4c63cb456bcfc08a6e69a52ad929347;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2e539ae2c02f0f0134f02bccab7808745ba6b2af10cee49c1d7f8f0e128a6fb530e3faef91f295305634de49e484f57ad8c63e344a5ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e24dd039f7779d7a49f4c10ddae3d35f23fb0be7f95e66a25b1c54abc59a31507e1609c7e00406d7b39003d56effd598344c8f9c083df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7e44ee85d3aed4d31c61cc24cf4d98e57dbb882c7bbc74542f8c68ffbcf8fc3cf1c5f63f770612809676f010631aeeba5ca075aec2db2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2c367a8a9290b724acf1b3b46ede30e92662c5ff6856c3aaf07f33da190e43d2eee30864c8f0c6d9ccdc5ac333cafaed5e9b61ec2a46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9646c9b64343d1e30b4594f1423e6d075a9e1f8480ff74806643bcc2f6cdd434fcb272e85821f90d85d3681d86ec7ffc7d33c7cda756f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120d07a4e127d3d63e1090166dbe6f3da47a457af71710cc13425d322ed20b92dfc8e3a6792dae97aff078a5fde13960274dd0c8eb3f52f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b46708252a2c357646332aacceee9712f592832123601b4be7a8d2d6f486b84265da7d0301942ec1deaab1c311bd0f2c8f95d4b231902f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fde41f3bb4832692a6fb3d21d9fa50a731bcfb72f3c68ee877f28fb9862583b5f27345b16b2b278ef6d70d0fb6c5cd64def92d4042939;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0e0ace8be2dec7c12042ca2ffba02493de2ce39abe9807117cb37fa18149a27385fdf7a3e80543796222954e4c2e1b42c3ef302c83932;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha808dfc162175abc3ffdf70a905e1a158aa25a49a7aa213e0deba38b0b1b10a077a4b1e090b74bcdf5c81689227f434f7e835b7f734186;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0087a9bd9104cc2d4ad900160092b6b5c48bec1e54132c93763c2011e07f24718755e8c5cbc0e4d35b9861ee96d9c50755497fed46a24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fc3eafd81e65c94f0e0bf8d8a64fbd3a23d64eaec5b4a434fe40afd09b898c0443253336a6fa655a58a3007580cf25a3abfb5ffc16c69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1949545ed033808e187dd000ce567e89d3a4fd48a0549b7adff6fddeac7883696c57dda3629c65ada7eb762b73a8ee2444321176901858d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111d1e3dbf75a8a907b3e61d6ecee5cfd23fd6838a8e1fa6bc1f02921968f74585f3c2f504034d67a1f6cdae2501f6c609c611a6d8b4727;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a8a7122f116f96facb1fe9a59ac7fa3663ef0b6f57800ffcb2f5bf0402daff8c6e9b3e48f457ad2b3333f61daba5e3b4043772c6250a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af60621401b581794ef3c6db117dbd778eaad299ffa8ca523e8f6c882868947140275f407ccf8e07070d1a8eb427f369410a2b0957ef9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b0eb3896337a755fd7aa140393259e816d3a82041dbc1fa02d4a27733b4e9403fa81cdb5147f8c62bc1290cfb9339bc45d41257b66c17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd7935a2e196813d73e60403a0983d077012da5e0e186088605d0ae814ee80c4cb6c78ba296d5230595a19086ff14dd1f841fdea84e9fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26184f33178490d33a20f74541aaa46888e9fcde0b457c8bbf5a4d0213ba7533941abb95acf3d0fa04cd22492e79fd646c8556ad458089;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f63f25b5ddfef2fba8105413da2dfd6d695346c1e6ae6b10e7abf3e6810faa827454d286edfc4ea5ec2636d23f8901c821ff42732d2c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdca788f5240d494be4bf5fae9cc57ab7945555d322c3d0b5744254410e9eed0cea6f2aabd6df5bf9f84d308994f43f0deeb2afd2ed540;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5a6028d932712d53c93482b936d46c08f16de571198b701a2c1e94784704feccf628db835ab752b1dc97c641af9d3d05d6b12eb1befb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea1f3098687c8d28e542db30ab884788a0196d676c969c92eb26927ea3af1066722d8cecf6ef70c9ca94683d631478457588a36ec05a4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fab4a2c5ae779179805b41b55c5dca6cc3af015a07e70f38a44e6fedaf5a97e2f7711b9530acf10a7922319f75f9a9b3c0079aa8f1cc3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a1626a003c1271c4130374cac344539cc621df6568895d66463d82be6ce51d15e4608bdcb5cd4a1fb572353d3fdb134af80bac9b40ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c885bd32d517a43a150e402a1598f445b14f61222b3f6f4936e5a4ee47c06d8935694af223edefe4141cdf46d6a9ce9a3c0bfd52655a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14efb88f3a94258411b766478aaf8ddbc48ab6c83742f8c13105bf40391c0c27fff10c5f1973b9bc1e35cdb9a8953f64e2b8056cb92abc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ccdb0ae9ef9cadbb7b801aa55cf952577d4ff9f18966cb371ef234596f0636dd9d865f5b03770af7087750b992138cc069fb27aa74f56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1565610980b7c0305c517a15ebdee61be9b036b917c61af21c3126015713a53c5fc4df47e7c83644926741fd50d674b385e9b806f129383;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a30e81154b096934107e7e0adf28bcbf81d287c573bef20bc5347f42f1039e0fe2c4905243c7f58b9bda4fb4d1d28fecdaeb3d1fd716e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc1df7def1d82f6b2f1c883ddd590cf8144116e8710bd0a4b0527a31a2d7d06640b2029848ca574b7fbce22c2529d558f94317df36f125;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfc04236e220eaedb16d2d7e600ef562dd4f25b522c5e76b1bb0f7d12bd7812e94d1591ad301729117c764d1989207cd0b65373eef4c71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f6dc80cec8c458bdccf8b12c8eeb1381e8c42ad7101271ac499efb1115d8823a4af145dc23526e2107ae5d03307b7865a053dcdfc8e0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd79d431ae9715915dc6dc6e1a789d453cf025835f4e9f6118d544e8d3d1a15ea492ca915273a66ab17e5a4d70187db6563b7b9b0d7a5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2892f01333ebcfed76b6528c9e12882028925e73bd6cc8642dbd1302aec29496c2a0e593d49f428794d6b4eeb88701faa6e35e583a49eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac4da3eabe773c5565072a4692842f4ed3f34bf33a5ab38bb22b94f7125183f16f61bf277ef3e2e991440cf8fb7fc385e2c46c3f143fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d5b10b9775fc4b77e4caa7bf136de72c99046fd1a5371abb72cf0371ce9f41283d56f81a7da8b160966bc60815e5133ee330437f2f89e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180432a11507dd7e79970af64d8d5867094ff60f133d87530119f2b0f7dd1cd8b9b40b56b9d91d41e59fdb1ac18cc8cf1138a9303798ffb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30d09e75b84f820b560c7d2a59ce7500a207f2ee8c7b891a65444ff30c47d9bd9bdd81795cab78d096128717e03892137778d9766ebbcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddb11ccaf10411b8bf18de46dbdcaa33637a0485dc3fe43963560ff426e97ed090c65e31f2ff76117e26c109d4da709626651fd282e967;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd50afc8ae59c85f1a54c0b7c694edfc91d99b8524d0edee9ead440057374c0cc8e4f427b9010e06bfe86753e3846b148920abc66df7a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35cde4686ab3adff85d7eb367e2d69487688b4048f7497ed2bf52bca05ca40c05394032c054a5260392a663978da9263d7c091b5178593;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf040414c0739324d3bcb6d9a45446ba91cec4f828c22b3a5949fb261f48a621ea1dd47e559b926fb42afba496bf1b5b90b1ce40df3d7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he939c511b01658a34c3475def2cb446b5d334f68cbfd37879de091c850eb7c9b74a2f61c84be622b1efae90d72253debea85b9e7271615;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19efabb218ee22c2c74b1fc1c184619e7010de41c40d272b7b18d28088c0f095e540c63ae55a98b6ade9808202d0228b964576cb8149e1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ba686e83cb0ee54e370c6b2e1dd724f78b8a9c6d7c228eefa4cf67197432ebacc932a22131bfad2ae00b77d96b6911238def793fe858;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1204e481fd28c47878e96e415920a618a4386782751f5fddc21d7e2da4531999970b3aaa6ffdd47f773b38df86c69e5c0e7290acd2cb935;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db6a644dcedfd91efc387bea96d54390da7969a237a514bf2aaf13c1c55cdd22f7584591d63424c948eb91341e6aaa7e6049639f4f1f9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had4b2abc4d407fb55d9cbf88529205fa43c2ec917180388313f61a4edee33c12a7cff35443255917a2cd9541b234ba5b77d5a1314f2aca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79c94ffeac67e09d072c0a23761d07600a981f846a424a2ee104f410967044631f1dc47058999ffec203bff1d1ba14176c88d0dd6e2622;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd708498b13f2f502face0fd6a91fca38aea38f853adf824b2c90515f3d0d99138c5c4a8988381f1596181b9440079fa16a32a36f6c6b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d1bb23b0c8fc2c282c2a19e2936cb05d186a3cd913e5f35b9e751efddd28300672f78ff06277c6f99631616e62bf9485c01eb78a5a567;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d295a8d17139705776cf4d0c7918f5859ae25f8b403e087f319ad1c8f8c746743204d75f2f5e1bf8df182b8c9397789dc1aa810c9e29e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179a3ed15796b8a340725dc53615071d0df917f97634968dc0ee162462b40b377d47d7bbc6f7aa705fb0753885ff94888d340619a1e2ce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1a326b97026c6ce9ca477793bdd24a90e0507c97fbb7ac434474072814b58c27b8b039acc6e50927759ac0b6a4efe30cf4fab12917afe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h974d1e88972f0483a75f13f69ef1e797aef77e62680b51b441ec24033ab68d5f36fc2ba3872ad40b4f0fa225b16e01845a266bd7ab6ff0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18104bb4a8acae8a90d9d181752900de3a3e021211e8b418dd88d00410fc54a7ed4fb6f9c517723f7ff645834d046e8a7134db020c7cead;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb105a7e542284085cfb2e46eaad8276df8696d4b516b6d8d8598e972f4b3780bd8142403a8262c12d0feabe49ee7c5c34a68447fe3806;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90b642924f6435d09f78d1beef7f5a45b2fad2544c3cc65817fb20df695daba3d42f184624c1dcd444628d16967fd45fee546b70d66479;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0faaadd8e14e9cd9f1ce8f6155600f34a8f9f3712ab1d0b23d9790a8a4025ff41f78d50074d145763a0082cb224c4e4a6b33d816ca744;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5632af6a19fad7120654845cfb4b6a3e85931f06eed331ca48b7fab8159225b82f494f8fb2d46589121210f59fe8543267292041215e33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112876d16a706d6d6c25afba65ff399d30979ff4805ecb3509f6198a0933ecb1b0f1a762524145dac17ef69a7f400e2291131e3114e1e8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127c42137ee82ef994bce48cc4c3138f36376234d7e9d43aa0b6c5f3fbb0d724aad7c4b82402c08202b50d8a2eb898160cf9c84076415ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f7a8ae4f29e17598dc6a3f8d36cb191896c9bc6b883a4993dbc2e021ed5b9e946af40c8f4cc4aae5ac663e5fcf46da32f1e54c63fad30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3916e71161de0bcbe54f1eeefb6cf9cad176d1f8c3bf6b1e1db51c88079ce27158e80aad9308ffb0dd4be3697508290475ab52dc884c4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40f0dad709bb6b8efb412a64845630a7808c6c7c45ba264fb6e4952d0a0bda2ae1993d90b53dcf07ecccdb9db35ad99e75a7369a5d31e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9fb4dbe9399316e1ffb69de19395f6de9592bf7d0ae35af24bebaa31853739b4403cf0885a1b34b70ed5eeb557ce57dabace5301ebae6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f089a7bc41c259a6c260a1c2171ce306072588ddc8a10674d8c478e8c89511e878fdcae8b38e7723292f7dba43c72ce88947c65c961af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5681e091a7a05fb0e14c9d55bbe8fe4ad9064ed37bc9930761d53ba1be903f60a5235fb54940e0947ee48e095532063be0cd1a986cc98a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83cd5374f978ad11b4b83410ea553c530f898cc59fdeb834cf275fa9a3db4c74ae35d1201d5a770166b0a028fd5c2e840d3ca39d6c23c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he098fa3744372d71b32f6f4d044a186bfa3a367e0d1686313576dd3aa7488a255776a4293774df6ef9394a4d79c6b0fbed7007da1c6bc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7cf8419b32af17b0904ac4e4bd08d0ead2437d2d7c8536668a5a8540fee0c67ff482d29d7edbc3dccea72e15af419ce8983aabe90c607;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ffad10c5e9e4445797e08b73438199b36450f4f25ff923d72bb3933d24bf364010a071d57a49658baaf72aa241354f3f0a5b33944abb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191ec837ac37e302bd5679848651e4aeea224249cbe66f494faed533c922dec7ba77fb97d2c6a85231261df6e81f845202bae91a3dff848;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3400616f676edf69d0542e99b46deec82a93380583ae88a305c2d7bef524256a9647a6023a6e04bd32e8cb2a29e8ec6b10ff3f19dc3ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b942300ad61a63ac7c1aa972b1aab21d9e34ead98c668a7651456a24edc5a5fba80793d9517a5bb6514ea9595404ea14f2db9396760b07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h950977b326ef9cc2a054686d6d1eb52ace9cfb72ed5a6f4f5983dbf2f0c83cf1e6b5dfbc09008c584075c4eb6c74400bc05b9df18b1b66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e5221b6947bcad854c09cf7d11c91c04f1c0dcec8ec5469a2c8990d9d491d5d53459660d1a9c5b947ac7b9190b44e0972144367168768;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87ac468225702403637cc89b66c7ee7ea1a751dd5c6f17635aee17d0b78fb8b3e1bc1e7ca1883e450bcc860f9fec788bfdc5d8ffe7f37e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdbfba9e2aa141110c47427309b5907a1e171e4dce73636aaab28fcefc85558ad200b221920a2155f79f3ad2868c51e9a623b90db3855b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90146945ff4ffe5c9323d91bae1a41ff8470d72c459e8cf3fbc5ac5fffba1eb36b1109751167d13c8cd4e4f06460ab1187b2f13131479c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd297dc4993a19dc5af4e622c39d6b440a1c53e9599fd35914e41e70c550ad4538782bd606f44c1c69fc65c6d53faf204f203a0abbab907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179211febf6aa8e181ecfff8af5a41e655f3ae761fc3ce702d4585d9fee440cd99d50d6d00d9cc1c6743902c546a8ac7a4e9ede7e3b90ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f481dc14844b8deac4afb4b5d8ff0434cb743bee6adca00dfb444d89e47e481c4cae62873503f182500c6a64c96ee86db7e4c74e4585e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8a05106be0409550d5cfeed963acd03bc426c8fcea01d0baab3bbbbff8933cc898a3e3c4e8b20b1c25e5a1771b2d2b9ec388cdf35a584;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13056ce51f90b61e30ed282ce6797bf6e413529e736005c006fe01ecb3d17019321e76c0fe3f9c3c48488345778dd1f1b20b764c1c93e91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfac4cd40e467aceb6c34d31b9273c55429e8c002f7837ee692e6bdc8bbae74ad8fe5b732372ba86f1c255e4f1e6be427b9ca76b2e8d8c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1278cddda5fdfbd5c95ab972a9eee21b54eb04a4b51e1b37ed47f46da2140ee101331ae6752e0e31714adf7041f6b4c0c9673834e0168f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1796bd23ce0c928c3e8b8f2f14bdc2c196a443df2171ed2515e2d2602b88bc3ded4f24249608f857b04358cf09011297e3a56c16f598c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77203c8c6013b1c766c4657024c1f6c5e2bab783e0b5bafe719d67a2945b85c2827757371f9134b786e4c0dae8c040061b28a0f878a79b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d779f5f29b65197982d3e58cf07d37a44185615de142c939f22cca6680ce5ba121b8158dfc3c794145d75be9d144f6cd703e98652b39ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14011540e2c467e267771194528824a0caa29538eab16bb4123eeba642e0e1dabf0ae95a8b913a80d83f5d53e83802c8974cfb67687eaa7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ac8bb7ee7df791303d36b16f706435619153b549b33dcb343d58fbbf260736afb985c7d810f460fe4f715a4797cfdcc83c714fd3584c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfdbea95574cc7134f7d84d55e1a67db7f913ce54ae4fa14825c6e757fc935c259b5fd0b7d90521631d45bec5593db7010a97c65647423;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h359beb03f62b8ac3a878025694ed274b2c0347eadbc8730fac8f9b17361b3895f126ee438ddfa4281766c5f61598cadb2ad9ecce5feaa1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a77d3e26fd66777972dcb844ad798159ee22e312ebb8489aab48cf2cfff57c64906cb99f4d872a6b74b5fdd6a99305e13e51601ca357d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22c533623a301eae19b2a4b01e3c5185ccd388ce89eff7f7c5b74d385005331ae02354a26596b739476ab9c8f439803b5b9fa44e192ee6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1940ac03426bfcc92db56084a05dd7aaa7aa5f6cb309b178b4da5397bb523ec7be7e19c8d97a7965bb2d5e8478a0648f1bc885ff5e8570a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bfb89e2bdb3958e544eebf4c7a6913c6ebfa3198db3af9e13263746d2fed51549f328640311a6d5e3f214c3da73417d035f3c0a238e04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fb80f5fb62473639efac534a8e2b337f1e7ee21731517f70711c36cff257fd8ade47dd98a1a63f37acdc16e9e83af6bbbaf921a73f275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189821f4d24038de29474afd2f633880a7dbe2b39fe7a220e248bfd47f190ec1b00a9489cd607d1fecda8d1b88b5030b551b6bcc856f6cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3ff653377d24ec1dd592974d04356b79afa3a6f3fbd6357dc14658008598dfb1aade2177e3f5b0eb37cc17fb1dff877fb1e05efaa5e6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h500513a8de84a3908732052ff186031a1209cf32677e6de9a4b6c5cce0dff848654138738e9696bf5214411db46baae115eafa7c787bd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c251cd3911c0580b58e6aad3a1979908daf31a8ec1917668b23e7b9f2881d55c99ef679cc2573a726b5b7b4866b0048754b62aef573c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb37354744c5baa07e688cbbb04a72771d1717aa11bfe57e7567f045f2caeeb2eaea734fdcc720028884d378c724c2eda08bc652350a013;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b320afec376308c56101e059a1aa955ce3768d6c9c2eab4e0a3986f8d48154cbbb9b5e829aa8418f0cf42ece175cd2cd0423a677e77d7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fec958aa0be4fae59773f65956b6e289f4416f18c3c052636361f51cd73eb7f066f0ed2f6cd2e6be16de679d56e9ac15312e9346a42ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c934d9f41995463ddc6a9a5bc0005e1d4874fd7ee1de5823ec16558e4290677aa191648bb151e56eb03ca26b3de97fe53e2b2f55bb891;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1838e31e22e5a599198be314c24dcff3b9ff5575906b0be385b40ccabad311a67e665485e2e12978c6ea14dd4fc79940678b0516a6b8fd4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ed97809997897c321631d9b72b5ec5ecb484fb9fbca68de1868a026817f8078cc6120b08f8d9929cb11e680a04e933491c2764dbb75dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8bd5d8a3f0804a2224e2114847651121a95fbeb90178352ccd9525939ddb236e4b3f8f9fa7604cbe6a5df921ddaecb5e3d12ddfa639e6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2284d6d8c61f6a551834b559464d3608d6fb0492646e5ba88a987af8eef3059311100a9976b1fb9fe778f9e7fe59b5d01f5d7a3db828eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d6f99f4eea9c1322c73d842c72f53f7710f23352be1851d8d1683abad7608f3c6c695af765c6689c6e87d8342fc014e2a5c55a0de017f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1cb5f08deb0a18dbd58922810da7ad2a9b03757cafb7f175afa723f724d1465fad877e60a33674cad7c881a3b535929d16b88906c2acb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e719e20aba12b8dc853c9618f2dc1be2d01476fa7a8b20d8d45d1cea2c484e75804f2dc3e649df0ee7dd4a67d4e1fda25c6bf9268533d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124d7dd5489fe36d484070209389ca71e463b8c699c9814d85cb8e859527dcaf825bc999af15671db973b1481ea39496b90e4d620080547;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h25167be39bf261dd053e9bb10989809799b23427e6e077aacef05a70711d3574f5a717ad46d3311d69d7c71555e47b521f61ef53eaa113;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1228e7ab5a8609fd72a1855570f93dffcd9f6b374851e1e0d9dc9cdb100d2ccadafae92da3bd768f4570907c318a041964945706cefd97f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bba4023202cda78f0e8faba02744b97612d4db12bd6f25684508d288aa4fa596989e712dff4cad0646be17224b662351929ec245dc1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h568ac60297e52d02d3f9edf95ddc5a2b6f4c55a3e05157236bc35dbe5a7733e653874fd8c05a77aa35b04058c20f6a21081024d641f3e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41023cf3e0e70f92bb993e87109ffd1383763b99ef128441602dbe4ad8ca33b3d551da9dc9409f1116919da5e1d2b56aab0e0bee4ffc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110ac26e4e07de9a53af9bb0299dfe1c252a03eaeea418176b7bf78a2de7150f7fe25a8c3385071bcc0819965de94c5b3e7b2fe501fbcbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7d19c7ce8f051df9b0ffc1d517284fe2f35ddba24aef0189b1f3a07597d52861c6b679adbd6ddcb8167f5415b3a94bff854a96f2ac974;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c91f5f1dea7a0d34a860c8d4ed530ba008693216a26e94a1d452dfffd1ecf08ad6757d90d4855bc1a25a649c5f4d3cb4bd44d309d7449f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c49c6a38ed7c0359534eeea4869a2aaa620dcc96794b0c2b5a8840ee02e20c870630dbb18442bd2c35781a60b537b49ea6e1fe43ef2c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e51a6a0e7bf24c0274e2fe0f08e495a02d82c5861fc3ff8ea0356f1c6b217cced8e048dcc66c74a7a9fe092ab6a5490bf6b8daf454bc05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h301d732c5fca9890289d948c16d89ce199af80c619a1d82ecfe52ab555b14afd803141bed189fc949fb96414023650a86831dc158c067;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e113278d4bdd133d572518b704a113080c924f2582ec241a13440737b6a620eea10229fa7e27ec60323c8d2d71ee468d507c2c1ae1c79b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1230593cb32eb3273f628451013d1d0c8a79ef8d874f9dba5f6bd42a228d92191afd6b8a4b1d065217bf99e8ff1012ad7a318b6291d4962;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6065cb74b65e877c2aacdaa7994aa960ba2e399d06157d910d9de8fd353db348e4f97a201c16fb43defcaf94d1db7da4eaa6f8125c5b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15beca409556957baeaab0a581a3accf1e4e995d28d8b8667d1fd57000372f5aba24fe275510a9b2efcf5690637c69bc3b3060b0165af19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6e803325d1afbc0ddd53ce8690b4cc93910b03d269ee497d300e84f4cbfb325941964c804891898c4e3c0d0ba5dea6680fbe5c16abd17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea0a6913d42727d8c2a8d0a4879a4e1cec5e5d5be30ebe2214e4c99b559512869bd61d6466d1202076d5a49e1cc436ad0af8ba62b9b407;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd541768ebc5a1262a687a5924958d31b2b71d4f25362f40e1eb28d356f6bc7867db2404e76a6879f77bbe325dbfa5e1201e210da78745c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38c5baa0ac0f480aedcd8b7c9fe62666c97c3dc5150d0c98867aa5ce841049ea3044b92f51c39e7d20902f2caab60bc43cf4dd9340912;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e4771e6a61ed7546de50a0f21e0a2d9eca96eb071629ec94366a49d0ee0ec8b24c15c893ddb18cb0dd889c06feaff6407fa35897589a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15790b0d25d263f3bae61ab90a40e5d1c117ccafa4cfdfd4b002b2457986de51e2abbf8bd42570d11baec2171a82b55852c4ceebc22233;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha232b76862f4facce8f42db77280dffc0e6122f529cd359e8b6c5315b46a668f416a58574c1be7afc5c41b7dd95fdedb4031f9098ffc08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h250db625515d78ca68680c5077065c1a4f2b909b657bb0862b97972cd8962dfd5a6b7dbcfb4909521365993f0afbd6008b0ed76de85c63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1682cac60b9cd0682bc56f11762cb2327eb84244e6fbb6f4fcee21d7fce26d25e74b4335e76daf841b1b75b6b417c18a01b31419cdb0e30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd957fb586de4edb3540c1a68e158e7a5bb85bc8410033f8079ab2f5a64c40dc611245c9f0f16cc6929e3e2b3550ce8694e89a9a351e7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd0d3c13350022257f1547ff3d955dc30f14df9384487e534a75058403274d6a0a373303c990577d1e6f253f52a92283c659d8f62135e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a118f071eed5a66dd330cdb53c4ce5172ba134a8dc485f4c60cf82b4f81c0c54eadf5b9674cfb8df2ccac2ca72191b49bea6f67441dfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef75ae81b53d371440265376edfebec317b953593d924694e255b13e21aad69fe555bb059a983fc72762a8c09364e7e7113876fca18dd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f0a93ad7325b40a01c5f2b4e90fd9425f5800253fea82ce3eb73bc8b612836884c0eb15753ebf6422476aeccd532c05f475cc1b722b33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddea24eccfab9d00e26839649cf24a620e510a9c50199856b9495d73571625399a8bcffa1b52fb60fcaf5aa5ed7dd5c18f460b510d1f03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1791069cf333384b3c5692eaae18736283cfda975bd2741630d5510a9849bf37fb87729f0de78c4ddb28562da0dfda5d60fa457caa435d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119da266e59da7010ee7d86c97e7fecd68a1677e37c1cb82adfd67a9f58a6075d5f62dfad1556c5c0b5c0dbc288bd2a43d371c420c7c2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22bff2b229be37de9ebdb4a2d86fb548569870f0a5257d56b8f486e89a1786f6b92538904605b2de921f108cbf3d9018a17a4c7f1374e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee2a274749dd0eab2c866ff50095ecad0c984274922f28b58483cacc4985a71c88741eb2080b564b4627f3745c89f9524e4dd25946fb86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f058a5e5b7cc87f0a8084ad8438922b53c68d9e6941539d4bf319ab4d69b7cf996cf778627a2da81034b54bfdc3e6c4eda6a9a3cbd305;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab5b5402aff1e0a6ec2a59e657c3c0099eea5ab58866ea81e4a5078adebf1d985d35c64f81f7cd29e3195a0ab4ce12c7613ea6c4f2f489;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa77fd82a560127cbfb81440a87f6509968e6f7e26b7fb6717566b192ffe414b3988553400c9feec169d730f62f99235d0724cb8422215;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e09e642c2d244c34705711512c95d05c2189940da195b61ecfe69b89fbcc34e1db6a6aaedc8e8e53b2b66cfa69465c7d0982a98d63d4e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171ecd8a4c39a503fc19514f905a81207b85b3a9fc7cd401806894c5590ac41bd3f6443398b7c48a7c1f999ae3ca65ad81b5e6744f27214;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191f3d7c36cb49daaf9a4216bae1781b77cea4f075c44acaa4d179147df021edf29674a39bbae428bf3e0e5476e7923d8c3b91cfa75534a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha63fde4199b8acd3b0b582bbbfe79e38d060202301864e125d8687a486b7242b62456a61420be76af1ba68d7221027886f307732c3dde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9bb64682dd3370d5be562c0aa0f6554381f9e6eaa363d95bdb316a0d1b84e800ee96dce73fcbbf66457c7170785915627c9e335488d07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152051301dc44fb1440b360264a350c9556b40d07efa9dbffd1060b76e6cb5694729e23253d1249355fc953cf7db83ca0da2fa5b7b658f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4895fba64bf2320fb72479f54a699633d3d341ddd93b92f468e09678415f9a2d38ff24c29591a5468578d8eeb6d3c1c8576b738318a80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2284f5ac203ff0b79d670bbcda0e33fc5d32a080a7d44c56115ccf71218415e800dc57cffa1703f4d11c4324ccf089c3c2867702bb53e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h72a1a3bd06620acbbec8adbe5ed42a7d516aa857fd4f9c1a88a542f04ca489c113f36b136070386695677b185a3610a64cc9ea70f5c402;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e53d286466eaf527c367eb04ee2c6e050a1c6d5c781e93ca187d2dbacb8dd1e27730f410f8ddcc71a686ce03dd323c3e1a669191cc981;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1012581d3aba32c32d9d57956d30761cbdcba56b449bd55043bd520c1e84bdfa79a3193aa86e545cc1f4bfc3a1ff30ae18083d71bc594c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6bc143daa0cb1c35c8cfece405c8f465387659dcf3c753f858262381a48d523410df0f1e1b3f02a7b5522a31b46ca37f6e2dbe14b2d74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e6d4296c50788f71d9671921cfdc83fb478c7d2da98d0af84ab4cab3cec226d92f815383819e92eab0dd31797620fbe8f89de5b700185;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e1d7f901de7427e6e0f9efb8ef456653ddc16b441c263bd2aa6cc58356c0ae7cebe3b7ec8d864f49c36378a55bb7d637bc9c268622128;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77f0eec805d9a5c2d9dc04feb136f37564e417dfb81f74d37fcc2fec0d3c468ecc7773d909266ddf330cedab1bd94537c60a12c90e5cf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d85ac1c3d7f1189828696ba1a49a6263a411081826477277b0cf9330c7ca3d9e0779a66fd0948286e1e5583d5d07511e577f87b1e45fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc11fb81688d3ed6388ecdac22636eff78d9bb168dfa366c4e48f9fe31c1c1490d88d90a140980190a0d1e49cfada0c8a621384aee6ebd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64a7695c2a42f4b51d3a0d532d638af8f18b807c98c747e02efde7f3bc3c492ce4dae8d528143ab398f82fdca88915e046c65197cc96ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d1cfc226061a048c34d581d99d71b7c4ee87f3022102d4859d035d565cb80905fe1b4338099538da29da2dbe4eafdd8934d9f03b5120c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1162002bbabbca21d6131fe01e5800f8bf466d995dca78be47f10bb55bbbfd5f89342ee1ba5dec2684930d04f3c940538632f7aeca5c42f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcc348926c955ce7e765299fde29292c4a02e258fc185ea0b4ccd0bc49fb42824c7d6548caa2e71f467fa0a794d893bc0f01d961798b7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce339095978e17daef7f08b4327cdb9e557cbba04641677da9cb27205630b4ee2fce2ffe4b47232d951881c2ae9313e1dde33401799a87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cd266578595731672fa17fec67dd11c6b3053e2a077ac36925c961d7bf0dfe73e1e43cd72a8d534ce832eb839b31c0c15005a58e54b90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df44793c85859b0153bf1f483682519aecb89e33ed6342a8021586387ed0d7760eaf618e75df2640320f4b0934851fed55482d70fffa4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cce1fab3bfb3e00c50035c987716fc72b8c06ec0aba39dcabb36ed29facbe47fbd0a26367aa12cec7bb44dab7f48cc6219c50776c9f542;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d98f903503e6e8ddf8a1edbfb7a375d426a67560a1ae1744ad769304ca848cf3fd6b6817df9536d2e4b8207cf25b7e5631b27bfa1d2956;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31ebeaf8b0da347414782cf6c5054addd24c9f2e5f2542c4bd3f26baa1caac0b7a8e0e27786d2ae7047a27dcf18325a70add0a5cab8615;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h949eb63bb71bff777fdf867ca23966db266226bcd3bb308183180fb4d5a84b07e80cb56e30b8e814392d87fa18de34ed1ec7efba583b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac8a285ce526da514de3c2b39040c10a663db3f8c45c8528cc6b8310c2c834d34b5f9e8aaee9af8e1a0d5b155794bc59e6cdd434d4cd40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10685011d36b41d5e0b25ee05c4f5936479f597e659efce38d203eff05cdd0e9124a2fe76108a055e7972ccf64ba60d4b4e976072c24d79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8fefb5d63ae7d1eeea6df4111b633f928f4e132d28be86ef34dfce44fe216bc187d1a43e9a27aa9c6314d64caecaae65ba345ee2925322;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e005d4a59f41525e7e99c5ae30e7970471f06b6184532a696f38cd88a6e3ae16705bbdfb8fba2b4bed08457ac53440cd05fb60bfd3c4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5306c88e48ffb810336c14961acfc4599cda1d32b43793ebfcd3d5d73abc951ec1e67e2161b06fa6774893d1260f8fbc12b275f7a300e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168015b0e8bee516e9b7d72d77bbde58c55c5f73181f72f565e872ecdb390daced087a35a0dac0abd970a5f4c325a62720f30b82e443c00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had0920a5288a10482a6eece6e35d84ed1dc17fa81f9de077dc06ef8fc6296e7fc8fec623015f156f530ded6151e3944b2735624cefd6e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2d104a5bfb315a734c98aa2931b857ef640061e90d9c05817a5de9c78354edbb9127dab2722bea120d4b55502f2023e6644bb1e31e096;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18edc7a21770756fab317cfcc02bb9a46aab219f4656b283df0c38939957bf52f913fcf9c4b0e7d0c9ce9ae8d0ba432ecddcd9869aa1421;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1e2d8d920e1558f5a2a4700b4d519abcc8d46f01e2c253551f90d3109e6f6033346b0d168257de091657fdeb4adab127d93d44c74b06b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28c1de07b3c856d5f7398c5d0c5a3f052faea9adb4beae752f12b0bbe68f471c0a87db5d647e8946999bd45e3b50ef431fb5d24ec5d7b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10298ddc7c477d5a99a593d8a35428bc526b96386dfef4a49c4ce424e39a918312c2eaf4de686012fefc6d2d33a71a4c9eac2a1e6c7d598;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f6e50e1ac5a9af308d129563d3242b9c0bea46697e7a61084148a309e47b8703eb4df4934e4f938a9232eb5241e902a74748bdc650daa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he868a69cf73e1d7803707c0973943c792ce48e39aa62d1e595e83eb9fbcff083ea1bd26fac1fe8a6be291389ff354308a28f1a2fb5e6bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d13b29502459c118ac6e1898178f08cbcb6229827ae41b972590f5e0ec885d401c4e3bd59d6506a7ad1c4843ea31de73bd8e302564b11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdca03d94e23233e8099eaeb2329e1a966b4723c5b835b0e790dff3b4c1a836c2e5dc3edda849cffe17ee15f2851d58474448946eb285d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194464ca582ccb78bcb26bf20c7e106b60bfb22f30635f2a79325779bd5f3c9f623d1f65aeb3c165de037d388a5a393d45471c8fdc7222f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19625f0932e59136f3b99e9446bbd718aa701106a07f29ffd66cfbf0487cdccb7db3d64cb6b6d58c1e4ad005bc99adc30f29c4bbc8d8afc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d5a6206e5be17a281c1da3aaf776139ef30104565799e2c04ede0638f50f95b5bd3ce07782e060575e73134c6b2b55c92e3afbdb72c69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e3914ff3cbd238a69e3d830b38f1329f2575e284ca25919f2a6fbc7cb7033a62ca0e3740c6d7af555fbf2d660c61246abf8392fb9b38f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacfe6f974fea43875fac625de604d37da0332a690db0ce406874a55ee6c4d773b71865e84ba098c084bf4a3c336bd3489f50f849ab61a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75e61720f3bc6270a27b131462e72364117085bb16cebdd3ea9d144a003dabe1850cf2e2eb8b96b31774ede86c0fc6f304ece6833905c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h994285fcf61c3ba2cfc4e129d3d0ba1fc2764eaf46814de6e4426efb0fb9a7f9fa89f17dc76c06a9fc86e6923cf5ba5a7825db0e8c3ff2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1229c7c2782380381297503650cc4e1b84665c75ac914f738f373b634cd9f70f7db7a9a2f5c37d7c8d21ca0e9d48f63dfb0f5bd4556e7e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b1b7e65f2fb2ebd24beb576efa6b805c61bbc2db7faace7db105fad667beeb093c17801bf125c26792903fb62b5ee682357cc9cca8b81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed7cf2a52cce52e443ad9a8a2a31f773d3b4c7cd5f8bc48755e0e4393ebcd5808cdffaa268a255368be2a1b0e382be7985efdebe073df3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36c354fc2f0ed386ba72d6e4b202050d4d177ba891ecbe0587356398221c085ec3acad15e1a3b851e4b0603fbfc040810a673f26217271;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd72c83cd775f79c162c8e4570ad576bfb42abed37bc108f0ea94ec0ea1f672969f586fa6f5f17a52e0905c9b0e3b86ca39703e47d30b39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c4fb9c0163e187b77c69b602911a92629b919332d1f869ceca3f2d9e514563d1c6b712a0a78a2b3c83005cbd580434fbc405b2c64a8be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5eda0d49087c58a45aeefe657a20b9ddee124fc137ad7093ac8f2b3e877d89902c85224b7a0412c62c225cb4a14624d340064afd96318;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35e2221047af4021170f85cd274c7522daf2b2b2187bef2d5cb216c3fc70deedc2845638f9b24420e6a407133a130badfc8c50cf93ef72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc30c7a452d50b2b5c27e5d1e0f9b9103cb82c722181d23ea5b22f22307f981e99a6cc1da31d9cc0fb70a54ca5de6d4b0a6ec18ceb5ae1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac973b93b610f2a459fdd220e411af1dd15fd4939ccd2c0862bb59c3e3cd397df2ff19c1d16e94b020661ed806c434b4f60942453149d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h767004315a4dc5f466c485c44123e5bd9697f2e60fc1a1afe31f4eb7f393beda2385e02ed28e906013676d506d94b9212849c1bacfa2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b4dd747056242768b9e3b46d0d09d06e1906c65c405c376d0f459f7aa6ded3d49fba24a4f0f8a0c1eb684f105bdae0120ecf3684d41d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f65401f2cb3a95dbabcd1222e52995fb41fd817ce2f23e91cbfffdaf880b2f9036369a40fb3b647cbf6d8148cbac8c0f3a61be537f4c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d5317ad91ec993db8126d323800a7b06285205a82ebb0310dcdcd80dd33338886cf286c3c4900a74a5b891e4bb7cfc6c5054166880f90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ae4c5f1b8465e20d1f67642d9e07e60997d09673235703b846f7b8d2dadcd3c2d4c11cf0341487236cdd23a01a19e1c206ed999c537e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8ab92549760fbe6b475c2a9c1a82cb24842c3aa85ee8b894ddcd7938fdb63c801afee0c50f7bf905ac0ea91837f1aa749f36b3c636338;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f924810031d44d31e1d9ced417547e6dc412215ac74c062d8a583bd996caeb5891d9afebaeee91a67b30e0a1bed7fc9dace394fbcbf19b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1888463e3aff556094a5f8409345935bba4b472de51163bfb4e4c4ff1d20a712fabfe41361c754347910a9e1c5e2c3c93c8fbaedb3d51a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c13d70dde0a087716ba61a57d17725b0e4e34f4feff887eeb855dcad3093d69381a0ff3139639167839773e4944ca9d846552166927d54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd32a3836729a72ceba1e1e9592ce29014f2d0160d790b2c48945aa3f85ada1e30dd0104ffcbd9486e424f13773aba2aff270b4226de354;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1efa8e9f868ff76858ed3fefc222d5c23c4befc4179b5c36be57207fa4c3c42fc357e9c1da35d85490abc10a1e733758d4056366e5d2023;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b3f2e837af4a073a3792317de716aa4419f5bf7bb8e443a3cee272ce219c5897b7642a66b1525068f2182c52f73881e97ce9ca2617881;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bcb944673e74c4cb96d5949b30095b5c5b8f72f94e3d3b0c0233cdc9bcef0ef1463de1f460056a6e96f8a861e73a680b12e515dc252ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da8c0df0b44c438c88b7ae02c2eb87ffb74b6a653e122ce3ea74c977b637460a667041b33cf2fa7497aaa0d1515a10b745413afb3419aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78ec17ef65f6b589502cd1fd3f2cc418e77c19f322eecd53f841f2b3b00c97d0ac409eb8086130baf131ff9b4c9733ca586b88295bca92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169bfa2d12fa856731ac9068c132dc13e3613850c884effbc6eb068d8e42a84e8c2873b5f790c797ce0e3329ab25086fb30e5db43abbecb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ea753ac2144fea07d7d87895a9d24ffd65c9af4a32c0eda35afd557590ffb58d56bf3765ef90885ccf42b0adba0fc6dc249b41500da31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h735074e8ce9a2d8d634478e6790affcb706aaf92ba5f683bad9fcd1f722575dbaf6cd71505ab98463e573d87d705e25f1db75062b25a8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13996c32ef1f02a85e079016d85393ec7bb94bcd27a1c391ecdbff7effd8b5828e6a4533fd9de2d53cac83fe734616664fb5eef59851d55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d0b344f19d80d8c36e798abfdf942df30c1b6cbce500e435d59a20bf5b8a0ec7f6b3f14275a968eee8fd919ef0877c347cc798bb09e59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hade9a8c8ba39d4fecc7469cc38e426605a7b26a85c5c1aa29f9fef3bf44daec75972673fb7b0a460993c46bcc5798729f575eb6d88c9d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h805ff8b6564b37a013f218a718e6a563601cfaa6b602492a28a5ca16fed5d5e08fc31433349e5fbace2d3a5c7eebd9022e5621d22a618d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189f49cfa528d028ab2d7854aaca702376d501208b00a3e0cd1d576480b1a25ebc220ea8a7ea818a4d3dec073112f9a1908527db566b1ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b8a005c6471eb8b2f4024801ec3cacb64d3ef4e941e3e331b692e101ccab5735087d450186677bf87e190ce0f308030529154df603a26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a6f9e2036244736bceca9746dbdcfcfc0b2f5c9b27b6b0a9cd2b20bf87ec0e983787b7e906e26051f292052e890555006dacc956d96cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30441437451c25db807bc5b3e1de8fca19c702dd5da748ec557052d1ee8ce1aca7b548058ba7219ceae7694203aad218dbf110dcc86475;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9b8ca175e310284bb7e69e779e995cd0ddae24affa4a235642e097665c2951a6107a8352fb0e8ce880d749eeab067c97e8125e7be16a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d7475e628fe19c8b7fdc8f96220902b0c25b1d6d5e919c2c228981ebd76162b0f36b81fac819bf1d28427e92bca79ec397fe43fb2a2a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c3e956dc8159377febcce2ac14c1899313cb7382eaa760936e0d9492a5d233ae2a99e0b5858ebdf580c6036d1b6f62b70c5747beab66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha01d82ba9fad6d80521d740f1d2a3c5f2dfc6bf3de1085cf33b411a0b2d768e190eb336c7dd5828817b07a902387b2c98719cbb1e1e34b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11797fb43b3e7783bf0b6ade42a4356d7dfec6729c82e30cc15f9554f977179f2705e748a80d428ac8ccccfe5e1bc33132928165feec064;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab5daba25d691fbfa115bd765939eb6aabfb1ec86e1ccd38b2105a218163fd66efef868e45820a4e8ac420e2bbdc02f1201a211850aa9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135a8d90ce85b96e4ad1ffb842237c96f53a8126e7f316203c0dfbc19304af202f19ac2a953800c97a1e48d565f9180241fc7e082160a3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2bbeae4b562f39ee3147fdf1e13c01d9a81b472c0e2c9ee9e7e633f88d2ba317c7c76fac1075aa9837a1e87b188937ea6f2f00c17afe6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h136c0dfe33b6e04286efdced87dca415d0d23a28e643e02561a31ef588e40dcc8422ead66aaed0e228464253e64d8311a2042796d658c44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf272f9fd45331a95a429c3a5bb724d8ffcc9324bc6180b309ead368ff8ee4d8d7b14402c145e6c4ac440615459f4b747f8a025721319b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fa21a5a47f4ebb771cdff741849bff8730314c7b20334382e397c78d75b1a964b7875243083c44803d8d37c6eb0015621da21bae592ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e1263dd43806673a7f26f390501b5d58de88c86b72af8e1bad764400f5a5ea856b81c7215bf52fac1d6ca69078b681e7ede08641f4bca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1a725e1ef03d680a7e6368e379a5a2c4606848ffeee13caf6c9e34a8a11d2b996fb11e3bb37bd3610ffba33330f4a6a68756f6dc17ec9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117c12a4dfdab4fef7aa4636a2878d93ba1c587fe39853cbde4458153b97761faa7f2d0e40940b4038b888e196e75c5c1e419fed267f783;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187956c3d31164e12cba8467c12991ebe8f99b8ca51e184a49b14950d3f1075b22f2b620e583ae9ab0e2484204ca6fa47c5eef7b4a582af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h471bf4dd5403d00446774ad8c287bd20128104711d9336b804e7d36e26d3845c187e8f71d3b49e961bef81d76de81e013d8e46a1e4acac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h50256e76f44862d5063083d6e41b5571f45b845ad0ee1f3f9e97cbdb5ff12efcf3925e5818080c7f415f892d6c60a6a3ce1f49c1f6feb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8af624b9effc3e9b7dda3a98be8365fc191e28396a3ae1d612c81b3119081be89eccd6065c527367938259a6a27df91a7608a290d999cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ef142c79f979aa392e586c09ae5f5c1abedb497554ab6fafc4ba7d8f8d826db12d5f78711c03cad3a02185bf38a101d34d12fe451fe21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34461b8e4cf5aebda310699e09fe2dcdfd6949351213d13ea2adbdcc7b6f4493a2e0f67b215b9bf382a26caec4fcc97efd8489c43a9f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1142c1a6cfc7f7d5063785292f031f4656734f0e674c40f8dc8c1e6ced998823178f2edf8a07d8140ba4642b8ada655d5bc52a540092b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h25a7fe0fe71cb32d3ceb767ca5b561c40d65edda7001a3b67df5cd9eab292d28d598c1e7c7ddcdf1b9e7605486e552bcaa1ee0f6533ebf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afaf77109fbb487e8642bc2843e81c86bf80f06f8cbf64ededf9426ce1d364b8898c6f932e5878bdee7f2b9ec78a77e387b5452d161ad9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126df28488220c797302b4dffec941492bb7d0447f5ef3ef1aa239a8ffbc157748420bdcbf2e7f1ff15b4ea82133e7e050acfa8d060bc8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e23aac0af1d0530237696da4d0d81d3b1e43c319b603b0109f2769add4295ffe6eb52473b1b63bfe5ac61589400e35457ab7c096b8526;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b88e6400719441fa1a8d0286330c4167162caef1441a04ee7c6f9b3d01902a6092f98bc13e6fd23221b484bd17a3622bfe1c1f8c51d1b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66723f287ed4185796b7edd44e5699493d6efd7bd0f060dd34515402018f22d00312192136954b75b3d4fa96459f6c9d1792de7792de6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1152254c768076fe7e165db3358ef9181e4123b69725ed0ce68539061ab1e777bd9d2a96ea52fa5051377d91eebfcddb7b9ffd90099ef64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h505923ab4441befbcb89414c2e4b8d4bc8fe8089910e1cfea83ae4917b4a8cc387bb67d80b333b543ae9d268590d46a8fc13ecc918e05c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188e358f7826c8be073f75cf3cbeab80e6d8e69bc16ae1ff07468848533504b0452f2b04ce841fece09f85609d467708ea4f1e397ae0031;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166910c5428c5cd67b25a4f35fbf0d2bbb0989d2be7336ece38b418309c2c99a2825170b4f3ab75be0ce0704bd23191871dc6a82a615993;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ef7f28f06e61ad502251ac77e8abf0d1d148161eac78bd456a97c6fd9d96af414d39196977ec24da3f80e7ecb16fb3bba9cbae16fdda2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122c51f53b4bda63bb6a23986c00092a2397a34c48599cf1b353072f3a1213cb2ef983aa918c4050f2d7f78ec4642ae674a509e9eb1c928;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63f60e365e559fad2e15d1d2880d572121bd442bd590cf2028f344bc1680ac274f8b709ee355562fb714aca20c91a70be71f8e7de939de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1745f4208a766ae9dc6167f5e68ec86ef2da34c6238d8bdc9980f6e368c85fb357d56e1bd355bd967b9644942958fb42443ec7d7686b5d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha72e2ef3a1b3c0fa2b74cadbd32244ffd5b78857ac5c0295db530685f4f2e99213f7d76c21a0da8ef28689757f0537ab0670c71ef9aac4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46047e6b85b6e9ec2fe6ec5059a49954ee432a9c11425f7b6f832fadc7343ae6edf45c5a93cc641b2b70ac1f28f8c27bbe2736d0e6497a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfe8bc3af08b7a7c2ee129319c5ab7886daa433056fc8fab9861a69bc5860885bfe99d3ae566e732f9bf8dc4da732ffef253e57f05074b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcde0eaf8b5e3ff4addeafaeb683c7ef41f2a15efaaba7452d8fb379fbc3bb72f406a37980929c8bc2c3459410ddab10f46372f84c7868;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a0ee8eb3d0cc152f2e99fcd593e67e3290a574f16cd4029537f29aa89d5bf976a941ad441fd7a7ee09a27c394b9e3916e8bb61212cee8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46405cafd27db231f23950af2049b214173b36cdcb7ed52ee1ef3f2d404435370cb8dedd9ee7b3c869c76033addd4e090698f70a886924;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1616e227dbb5b1dbe4e76ccab225e3488b389456145009516cca705635c7264d31936199a174c2e82c4d0522d4a69f5d9da554ef9bcad9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1615e05b22314c87d36fc167e940c5f951d6d471f99096b8ddad29a571dfe0194cec81dc1fad8fc931ebb03ad3b9b98626b00bfa2367abf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1c34d38c67ecf19ed8978eb87f35f5e931e191667149b3ebdd6f540c47d844353b3fb965e10ebb7b9332823fdf74ea1128c164149c3ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he10fb93df6b6685afc72b8dfdb0e610543ead6bfebaba2e86b63276f76e2e4b9108f99bcef8145f40ed1a2f4f0107d24c00f3f6843e40c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec90ebceb21482df95f09cf2e49ace3ec8a6721f3ebad4219baa0548f63e2aaa9209fbffa28e9650688749930d786edfd84949703b86c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3686eac087e87434bcf595d1e96ad8930992f4c5ffd11de9356609ae2d5b4b96fab6fe6e0c1fc7f42b9b3e8a1bc106e4d7d1985a663b5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1286c7269b5f6c3cd473bc33a5f0d5c282c613fabb18a043d194be5846d8cf29546cfe249e8dfd9f454616985e909787255ac8eeee6f6d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69fa1a756776c098216efcccfc3ec743dd0163ab4c377bf6398e5bb84115402d13970a67ae781aa6ffb2f572546f515f34ab3575059b3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1325fa2743e20049f33b1823315eb733ecb43c723ceafc1357968f71b794ca9cde84393249b27a6e3db67a57c704d9cd382c3b8b5d5bda0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d9e1e71f51761f63597fa411d1da1f8670356305c16d84537791edf59cfbec277fde71ed386d1c8e673aa8687c06809cbb7b8a5903a8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cf0039dc812491ea5bbe215a43e88ef271621c7792829d3bd680acf31eea92fe9464c5964834d3fb5dc001d50bb5d3f8bebb255163a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95c97c10f75867b24af195158df992e2d22e2778168de5bd60cad1f22cae976aea19052971e957deb8d5eade3a62301d934e62eb86e6cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c1828207d55b06dab43a8a9198d1750f1c582564c6cd8cea8c81b8927248ede2faf066d9996f036ed243e24a099a2af6226a28ddb1df9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8733566c7cdc96961b873dcd1d8265415a4846cb42fa8f5791b422e513f7f3aa44ed65b823bea5ffa505912e097a8e50d3807d3250dfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c89452061113f174f1c6cb41a70743da9a4c87e0eae3535dfc7eb632392cd19f1d07142cf2b00921a325c879e675a9d88215ea09adbc59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67a1beb57158cd334e87de055489d208ff1708e7775b2312cbf6551e8c9768ecad54a42b71bf53b87a677d9e4574c9152ccf7dbdec520;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4afd9b998d63e3e4d43cc8c2ff629c2474d8ad7798fc6169295852aec62a37723b942a74b90d3469fc9f6a3bc8e4b746bbdf81c16b377;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ff34588624d1d87d4ef49ee822a896439c0cb550f8413a66fd30b9b2d1cfa64c2815a18eadae1fb796faa763a6f3139109dd5223156d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195dffdc7240fba324c69da26c30709125529647f96283c0096b40354e317cce1f26d20a410306c5435e8cd960799ff789e26833f3b0684;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40df508ffa87f3ce3ce3ab8c817d1313a30f20dd916f2def721e2e2f674e7e98c2e89902e5e8431b38bd9dc31e28c44368a3b109128762;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5efe16355fedff785adb477a66b3016112d7555f5be51ab032326ffb7ca99ca3c188833b77ad41be58dc85e3810cc7a5b7e57776c0bf85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c9c914ac087a991c4ed4370a6800420046c0da75715db97088b3d41decf3de8f088a1491f53f2ecabceda219fd9aa9915e16078fee43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f26a320e1efcc13e0fe26b1f67a43c9569d5db0bc2682f8a6d579258d08d77a4b904d8ab54cd11912d82ef84d820bc59aa59360528654;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9db4f5d97177582456e7915addfc9164ec2eb6aa06ae9b97f4dcea11c85e92b37e78dce5127555e4c699ce0584523e67655cebd91aa235;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc6507bdaa5ba073759448e42fe8547c73fdb94285ff96bed01c428eec4bb560ca6234ef5b77035607242746994141c82c5cdc6f0ec500;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf86fb4cf9e9fbef03a19f97665e9ed7119e3a88b3ac1d6d6c9c87f7ba3e5c175f6ad2d00450c7a689802b1e4829e02ffe202ee9c6956c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e5a8dc6a875d76e2776e76d1feb4b6a6b5e6758f1191af48b39d997ddccb0c0f45c4632a1b107597887af920fad4ca791394ac3788cc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd14cbe06560c5003f2cd08d607a4845e10c9a6f0ff4a0bee3293ab3404db2d1218228e8de562c8d03400ed04c82cea5e909c935930d2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0031ca16fb67378fc4135652995c9ef51e1597e3c04130030a1da13a092adf9ac3e0c6a321596a22de9300bfc325cadb686bda323306d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129aae9df3009732247ca04252de6160cf49d5d499f8d1aaca3a257b58e7c10121f4a0622635b0b5e26602d7a876887e253d8491d7c897f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d018343efd5044b308cb8daafb5edb577f2fcdb45f4dec9994e479cce72629c18ccf6fb7d8745fb9098bdebd8247c24c82f32b0043710;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14830a1d0ea1ce863ca09612900ee799b60512b09dc9188a3075522942b84ef08a947ce1097f95c42f88d9e80707fe4038d70f800f674d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4947151dd861c80a5475438f7e1ea9ec4c22162e5383a0038cdbee339b9b6f33b0707afef743b338a76f1a8159458a33e704f227e49225;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ee89040d474b4e78e91444c4601cbf672e7eecae57ec4e57a5c40466f53ce8fd8bc461d9b891550a4fe3bf5b41c12591f1daecb3884e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31cf5ccd2e75f12960e32baf14c88dedd97e27ecfe902be310de881fddb6d3d102605c43475022d9aa21b8e63406d9b706a59f50520920;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b71c491d267bd479898139965d6c366ca17ff087293b1575af4f3f1e03e08e12725c63dbbe872e82e7ca4cf5b223a82dcec51af313167;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186dc5abe69face1493690b1f70be04f08b85814cae74e9d59d5c2c15b061aed03e0a30710f5dd7a6b820bf5b9dfbdacbfe83ecbfba0092;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b266e4dbce0ed27a4d9204082112471d69c79df9eb1f2549a2e31ad5f5266dc64042d6c024dd1f41d66fb5e1c1214015572df9c7b012;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea51d8b50d274b8dcacb6da2bf8ae72c227f83cf678e8e2171016589283a1186286822cc68a96b1e8c925b91409317cc9650326e44c20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d72701b72a078fc25d863709facd5b3a88934703c67598a12f63ab758166c461b8c3fcea7c26205767a9e4b3d4b27e2ef1a3a8410e5df0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78c7f6c00d3bcc9d94efc1fdd0d1b140ebdf09af7d992645c193ffc0ae88aaeda5431c01079eaeaa775f2bd4841b31f1ee9a94c1e1973e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14afec3deb1ea92d7c5319876ba5ed534af5e61749c4ccd40ddd35ddea5232f4c2a216bed4e977410f7baa50d8cb11ccae1f86e4b60165f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16efa517517481fbf80fcec60dd6c3516be07f76f84121a5652285aa9a30e953241017312928d773a22b903feaaf7409f94787e4c97dedb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c01030ba85cdc31d7a749cf8064a1bc9c4d0ea8a2897e56933d199a14756d3946057e9d99f6351f523b55522980582004d1d2141584b88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157868028d3d01021b1e07a7534ff496761e7643cb102efb07cfcb3984be1574a221c0b9384fa1d2a586423cf407a8b09caa82942dea30e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a9a9d9c692625bc260e9346b8132dfcf1bcf209e18798857867eb0522416fd8b98fbdd45166146cc0bdd8dd965cbe167d6f6485c1c78a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8852fc6c35d3bbcc29f698198a4b032178f2c6d96d0d2390bc16df8c33b4d43add5bd2fd64fe58c3114a29653833cac8042d1258c7d72a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1675849af44360aab0e3840d59498208bd71903ada193480a2de2acdc6aa6be3fd6e43043b3f04c94135b08a1de9f12ac11cf52a3f400e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcbb6641853162abce4359b8f86acfbe3f899a5009160433daefc1a8536e430a9977cd53c5b122102913457f8209d1882c410a91461cd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114f8ee7bb4154d07f36503d631ba6722aad6db40b2db866e8efbb81a3343aa61547a0d9b005231aa945d522993011453be835966cf00f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10313ad7de11ee2195650f7f716f35a4f09eb4249c3245b5fc8baf90a0061ccc725569b14659f58c7eefa067597384c58d483a8404e554f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4c3d3b1b2f0ff25786ad83e6b639096f55ff37d41441b280586315fe2a063c2026532c6c02b8ec00b3c8771981c6ce5ca065b21bc9b91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43201efa4cf59c0662ede0aeb7bc0278f13b54a66ec16d2d872e2f3ee4752af64cf86d75a858545e60147b7c49da2fd1d6e40edefe4554;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2a9f82a8ac8e848cbab9809d363af3cdadaffa2e54d58dc9aa69d3d92caedae09323e03337e5680d6b33694b17a0aa5d39a9155ce187;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110a9658cbb281604541f9d81baa101fc260767a1d1bf2d93589e7647d3c395a6a1d9ed66af20c4e1afb088dd9ea6f78d881f9499014a2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc4d5af37ef9cf752ef2482b86a41432f46ceb4ecf66de7cbd949b502342836dc1d61e6b6690d965bb7d7f18d54a1a816e2981cac6979a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d6a032d04d577f644ff760e3b05373794cf43c303da306ecc4c90a052f613fe06705f136b597e43928bf021ee75748cf3433700275f4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16601f58f3ab658c95bd611f4372c9cd1eb92717813a60dd0aad0351a9f69ceb7790c449145193e330cac745df37149f2ccb39990f510fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101fd3eb82c77bc76ce3824b785f680c66739239e9844bc9c4590a384eca0af60d1232455daab08a9613010d6c8e1906b911ab808ac31e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170c49afbe851b7b64195b51d74a05890896d036532ed874ad6d2afd54fec41d51a242f3453a8110c223b71d4c707f9c9112c4b1c0b8274;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff69db039d46a7737fed5eb3bd38d4e675aed4ff4f90dc94c7a92a6132a759f2f5f9aa80c7f188944411741217e284e4535b3656b886ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1594500efbc0ac8118890a45dcb8bc559738bb8eaf61bf2da41b0af1a24bc81edd1ec49df6ac2d31457c4c9447438e3944e03a85a524a3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf08faf5872f062cf5062cb16b49973514dfd00262af3156cab77abd33e83f21a81a0c6c0acfd6c5ed1314065d886329dc0120ae5785fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b730f39621c4a469106cd7166b59754af082766f68494a8568fc309455ac6586638f1ce9d3f9b98dab6f2c521c3592984f0ec4162db013;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h221de8698e2cfcd3c0749a91be5d49d87659ac7ea655d50c25886717ed4e3440146c6400322d556bdc2396ce1f27d0de5be2f36818e0cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b678b3314102b08b7c10f962d0b223ffcdbbf2406e50c8fb443d89233f92ca6683bc66513164d69212668142c40a49f3a16e70a1b2b8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9428606df7568523e248f93cefcc5821c4fc077812f70be8e618ddc19e6db2d081ab14d581a9f2329404240b113460e64d55b67c76e66e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1850e06b61190bac2761123848f14dddc242dabb0415b55642a95eb743c42ada65947e1c3eea045801d875eccee25fe4a3b23a64d2418ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca9dc8141a41bda4d586fa4fe3ee9ccc9db87076a1b3f64e404664cfd302acef7e3081fa23fdaee38caa216589bd82b44ec4a748d50bc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9bf0ecd659c473f0461901920cf97933952d66624a696327f5b731721d64d8a8b643671639deb0418c47deddbc4a3e114e45c567235fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bf9d76b841b59899613958e4f7c1218bf498a9495cba7dbe036ee8808a44e4e78d916f92c01dc14d3a70476d5f024b047def94ecf68ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d6bb050ed6cb68e973ab9d3f790bd5427acd7819dd88fb8f5ebee9ff192a318d116ae25644322ceab7aae201de55702e6c99b71422099;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h516e4f733e19769dc07aadbb925d33b814a035c843260ce887d3ace577db664ad059a35127c65f3c1a4aece0b2631c87c397ec64c04501;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15052dc13390884a7f2d2c637a72513663141d52b488ad1a91a9bb8104d190e5eb92fe818259847edcad4d09e2a928cf1872dda998b64c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18686844346145770bbce3986eaf7c68e017ab741297dd31e8520dc8eb8f4c604407d8890a605bde804b9fb09fbe6d4aac670e323eceffd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5750ffb3697da831ea2550777fd1373d142eed6521474b703218f440142e17f5052434e2a55c90f9ede9da8dc785482266d86e891d2fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1f8af76d7982d2cb7026169a6615aca1d46e4fe076e660d6059349d286c8ab452cd3748647f684de8def891509290c4da767ffcfb25d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd8cb198291c2cf6021c3db3a8ddb0aa092f4b4a8f007433dad516cae4d3fd18407e94e5ed6cea38f88b24e819363e9b5f05bdead57afb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1f53d87dd0580e6a5942d088e880c108a5da9053ad71f4bb24c3ea452788ccb473ec5e561f200eda1847b24a1831ae9f9674ae57d04ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30927e35849771be679405a9fe7613d092aa6f7c7f11dae3e51868f1679d488272df0ff236394e351588886aa5cfd8585989d5a95277f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10eee3c4dfb62f68f7a423832c7ada7e83702e74ca471283133aaa0b225cf8c02d0ed3611319eaa06780ceb2edb035d9c875bd08fc31e62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acc9c5a2ef652802f3ca6afa36a6c5798d356650dd0bb8d0e020a942dc34b2aae1c45c632b798e0e4b9eeabc52cc3bed76f7cd392b9175;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63c540f1726be476414b33e23d4c2676f4485e741dc33e25199275aad9338a6f65baeb21877d9eef7fab667c5f021fe256bc5c81b8bbf4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84d9f245fa4c0000fea5ecf50e4c205f3ffec1f158197160dfefb1b9b615d6bb4a087b090b33e2aa005ae494ab2c4086946f25b6b2565d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d10a06800b2d15df5873a089dce68622dd625afe18fb801a20ae1601e5d52548463c38eae0f57d196c88d81340014a579d2f7be90c5eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h283c3f463d317277f74ab5a98ba0c5859300dd0c52455e82b01edd5b8c77c70cd547b5682a11d821419055f343b0e282c98664b97c5b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18fd399a84a894be539348570e978b1da3ebe397da17b01bc5ac4d1b49c10b8421cfdbaf5c79109557d5763d47bb32ba2604f76dc984bcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd0a823094195f4c908bd0c17d41481d428aa74e66ce3f616482fcb088b2cc1c42d1871e9db3c99e5d6d8ffc504721a8e7e4e436a711bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e02d80e08267db67bdad5232d9e3dd361f36bd8acbbd54ebe948cdb57aec9354802684110566fcb4b3a72e3fa682d60094e3b0e289970e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15976f223c5fa32e64e298a0e04bf09f00edc61ce05d36a3272dc5a4e41c30f0d0408eb5261b00ca22cf23b4a1455ac688d53fc303ba73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e51e80bc02678db346c494b0c4112e8e816748c9c45b0fe7cd75f32f63a3eee2a04962f2cde2b67686e15e0750bedfa24f3df1a277506;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff30e5959f3ddcc1c7db5ad408d694f1e0b36f8eb70fe47577590a71aad7078dae3751afec4f7d84c8b9b9588fa47bdc502da6106981a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189219a2187aa81ddcab9f66cf5189e79abce20aa8261d1fabc6224b087c75dd5b5a1a683d5f532b787de7263c7cf96a34eb35c7e04c85c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc421d98c0715dd304b35c13c6e75af0ebf99cc5e6687877c99600718cd3cc23db4bc18ae95e3b985b0a716b0ddb57dd7679f9b06aa233e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9db3fb3f87e610a81f390386148473114fc508bfd68cdffe6a3fb175ceb22a27d6cd8e1850961db560038e1be62c02b11f4d2b07111fd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h511394df1d3a16fcd4f1e25954d747342119a8940293c74712dc7d3edda6911fecf20cfb0410f0806eabaa569d9951c180495ed43052b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b2ac0edd273f0b1f7931d34a260cacdce3ececc71a35538249d7bc587d0944793e0184b569b9c502149ae75ad5d6de1dc1d52a58aff39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c5d114b71002a90af36222723f277732d74bac75dda17ab6ccd9471fb189fc8342fae5719b8b651ddfd1e9222bfe1d84ace89828f2450;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117986d841e490d064cab66704d5b5b9381963f065f5f16bed2c2c2fc45a5f7949614fa803600a749414a67b6d0d52742ce6839555fd052;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef3dfdd73198dbb405d3169485db0476e91c68759d2abc30117209ecf2d11a0fcb63a7eced42f1d6a7a5f02471c0c8e2542456adbacbd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h265b014de28a625cbcbb617710501aff2a1a32d6812606b557d1df6bb9b1a7864e14fd8767bff4b62a733a1a81b266760644717d6b9749;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49ba883b90ed3920afd6b398868f69bddadf9843e29f1a9c2216f5fcae6da92325cdeb7fbbb4ea68aa7e15c122de32cfa63f4c6475b507;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e39314e94f30c462755728e8e19c1edc819f22bd23b653a0d87b8c1859b3d22a0880f173892e773232342a051250c3c9d00d0f8d4c90f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc622d4aa52dc19fbd99183f656050cddf866ec54524e28261272819142fcf32ca1f0b8cded23fa230895dcbbb17890eb266b31b7035603;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa0b988e46cccce65d84d78a897fef6693d736c641dcf8650974a905e55781a9eb99bfb4f6c5d556871f85c396960c1f5dac03c5f0ba22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0e5487b40beb600a885ddf746ba088077a5b2ddf36e0259ba754ed732fe897592fd1aa215ec8d5f38e1cc8d184b1904001b6771515bb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117eb3a63f1c6b4243fa58d664ca21fbb461030116e2a5c82d24266cfb6334d1f81336699fdeac2471d4d905204a862506382899946bfce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18446084dffca6c2003255363c64476443b049524874d9af7d9ae48e59c4c1b7b436f0977c4c8f4d6106b9318c6872a81f90e6c7d50aae9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c3be31cdac0f13fffe9b27533d2a3388908d3ce3b9b31c8dd9389c4867e024cb455a102231429c82895161a5b9fab717798d7f1a496c51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188ed372d760d087f308d271f7ecbc675fa3e0a079388855c859500e4d5f38f3917302f476480806b5fa149d4e038520011203005ebb0ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba6b610bc925e1b70cafda3bbdcd581c2d7c25a7791336f0f9cfa412bfb661db3244d32b20dd343aedbf770f333e992ba2ba1817735367;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ad23841d02cc0feec3b2ac81882c97be8c096a7a4b7b7e33d0217e47544272bac1e7d8ce97fd43d1fd066ead9748bb0fec67462aa9448;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1927629cea833197bd90dfabf6eda3d46848807f9376f547954a8939db3c920a1393b36bbc3fcbecd5eb1a3672700afcf07445a271b6356;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10001d751856a9dfece23ba3bd06cdfebc0cd206b1714d4a81e5c79443543c6e6c3ca0e0431efd225103086e072f44eb354a970a1c85cc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7dc7f002038ad367091533d65a6074622d19a04a84d612f37b4fbcdccc4b0bcb6f13ad48f59b995397f03fc137ae3c65e5035ad9fe1f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d149dabe01b075ef8bda71a9e7f082ad465d0a71b8df239c51040c759c88e95a95d41a34f5e15c54897df4eed6554266e2e772a732c26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd4ffb22833ea18305f7b5ad898c6ad089fe651920bddba6267db70a58ee4164fe909159fada8310a237c58da3fe6a0245566d8ce7b3b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1644ac3a608cb77c14f7dba241973f2267f509c3657feb2dac9137f6c6cb965477edefde6251e82440017e1c2cc251accbbfd470a8853;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcff9c387d9caf958b4a67f6bf70f648302d1ef0467c2377b8ee7a8e4ca213f50f559073aec75e536e23bccd98550fd4989bdeb604a40d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc64feb10575f4de03fda07fb6dcb92d33e2bc27164399010f2c5a53773834b30589a78d7c090c8074e6b31b98dca67164cad5875060fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd70dba1d8236218a67e02454354fd652f2ec33c1a16575620aea304b3a500107cdaaa13469b3a81bf7c2fbcee84fb88ca598381d36e7c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e35aeba5cc0150f10e8d64a9762eee7587c9804a6bc1ca07d57412294977245b36f299b601b3a4c34f24b5cef7e9ced57ab6fba082ed75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96f805817d0b75a996558a94720874823a609eb0f0e75148c1a4d75142aced2b6da2b72fe252339c83da89c7e2add08a2dfcfe25135ec2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c3c9b819f0ac4bb1e621e279e2e5c73d6a2667cae58e811f29ff51a233885599ffe3aaceebb58b7c798afbc1a827a19800ca6de92e3b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e2a3af4e0b9b8d59070488e28c7846a66636487a4d19ea385d6782fef519a69ec10e9229f0e88553b97ce7a5af5ea4e60c815869555b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b54044b44faf20cfa7a15a26da2c5f388c7dba19a1ed33c10bef189ac6e5a1d1b5bcb7fbcf56eda4bd417694bc22651c08d99b0b3c7190;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d7d6ec970e84d017f2de5bba6150afda1fa34c0e7d6037f023dcf6f16558e846eaba8b460458464f5a6378580d6c51d8a5b7d36367f40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h921542630c4a6eb17c8e69045489001c87874e7a5c42b7cbe0c637b367bd7c1783b42ed39414bd0b4354ba2f06b3681dbc2ef2069038dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3380d01abad2ebfa20a3b9c743295e8948175af8330a8f2bfeda6b7e0b69fdab70747c5eed8d65bd87d2a6b5aae5538536d9b45ce07e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b98e7e470f8761d6a59859845de68f1a55aebde7f0f44db5b4ab30c86a52cf95ce30a5a28c164648e0e3e3ddfd5cdbb41fa9171ba4c36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94452cd9cacc19b8ef2ffc8056436b4b4c890cfb08e7ab8aab68237dcee9685621e67c8a88492e82f34e02643ab4f80f3d9c1394de43d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2704ce61e40a956b76ed5c2826d1e8c178d6d6e7680cac0bc2f6501cb73ea65f8f42b6998253cae0e4cef634f6a4e919c02532563fa297;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db4df661dcc01f710c1bba273d125981ec22b8eba8e9c35bbc5536f397aee09e45fb9800130998181091459351b528e90ead997a7b5d68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb8a6f6268d85d36f78608ad8150f64da19aa0eff6e69cc5df16515593a61c029857dd639fdc0cd97a201fff9aa5e02914ff6727968013;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196d0fdd0289a41098fb23f25158ddd24e6779629cec0c6cba2f45c877f4b8710c81584d947b90fc77b0ab42efaeb4ee2b4aed5f6d90fdb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h837971500a4e5baeec22ae085415c24f049bc1c38e043a829edcc84e52096932c2e53e38ca932e39502acc79184cbe29dc16317f905d5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9286c9611f4d9416d3747ae6d2b101d6a8a475dcf479fecdbf827f3f9f5fbed8f2ac0c7102b08a368bb870288c7f02cc17d8f26522f217;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h311c7beac5227c3078b20386d7f733e8d2f87e709308a328decc2ec4b3ce4ade628f828a295cca29b81f88379c710f158c4e4b8a87ea74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ad8f6030de952852701d33fd2fca0eba9e80b1b01f7ef662d2d5a71d72b976a42109538877d71db55b5b96d66ca766f18635377cfed76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8df21a5869366dfbc4d1623b7bc1f5b26b1bea808afa47bff415c642d3576083be77c2170dac1df7ebe48b5208cb0117f7f55661ff5787;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a443344bb36171a1847fcf75ec93615a854282a1539521216f88272711add0f2406fa3fa9ef57da4458eef985357f408ddb7a562eb6a7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1055c9c0318ebb7c2b879c99b283300458f912169e7ef6d1968dd5011bc4b83bddf9920ab022f893349bb85f4958fee9d2f8f34ca2d54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe7ef234526b429f2e0aaff9f586149dfe8af5eca3626f78db7120635e407a65c09cc152edb93df541add0a519fa9db40f15cb207a82a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112540969cd58b77154f11fbabb924a9b111db911f9aae7a03e19da5d92007c93c53acc07d87b3fd3ef3edfe1162479125bf6845934ef25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dc81c7035765dbce638480ccd2a9b5b9cf5eade3d35007a610a270184663e4ac71ae72eeb6bf8d9b98d937c0d30ff487f0c6db292e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df69ed99f34c847364251828967b7cbb08eec2229eb03b7233f2c69820330f9d4d1fe4c2f9ac31d8071d543b14e1251bd376d8787c9678;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1755625f6fec7f9e9819c2063b84108f1883da21e8782f61dfab1aa798e3faa336b187172a405d50c5b72f81505ba295c3cfd1dd206cf4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a47f7b8334afb543f41e6132a66c1399b21eae681a055afb057173bca1f2b2f147eb54161196d6a47176276fdb7ef50a5fde1257af137;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec46b7c63fda174a09ac94d5d7271cc810ed863603ce771087abdc000f3366fae1078022735a6b8fc80e2f41b111a08f37ec5bd6911039;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a39407565eeb65d9294554bfe7cd5489eb7b52c8d3aa3bb56f1dfa585e9d480c2f5a20de8ae6133c98b0bdc13c35fe12617f28fd26f93a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a9d51382d004a4a9d81a84762b5aa1e609f48088239531c05a68b184c3963d2a908802f17700577be5084c5b2be8a4b66529f9710b64e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3afad952579835d2d38943b5661c569f3ee8ec7434065f15e709b641ee4ef46b091ad87690c2d7dd4a8e6ea6ef522aa1960afc234804a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11199f2cd6ad98124649e6150cd432f942699a82ab2b6e70cb11b1f2d63d0831bdfd32e68c4d12128dd042cf9b21e6e5a40e20c4a7a181f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf01e3f68d1f1a485b17228a773075ea2c38e6d86cb53d4fca1e6797fae2aeb74abd9b96b0a60b3d829aabaa9154bbd9455a4913ec24fc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2792a1f550cb681392205c54e3869bffdfa95b55cad94f317ba35886451f5c4952705864a75e202e0b19d0e78c68cbb2a8e9d02039de2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f1d6bcf040740d43f4d34f317ae975d77b37adfd0a8a0c6b1e4e2c99ada6b8a3eb8a924190e0727641149a6e1e4c98b984ad270e8e82a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8bd14f33f32ecbaf33c9e9b91eafc05ef6abfbb4eb20ade1705e99b7cafddde601b351c53812d55fa47455ff901479c058807cd1d51530;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e322b4acdf95c80c6e26c2a5269c470e911e76cd920b5bc72af2b5206839af6a151f4770bdfa52c05fc73f73b199bbfdca04edcb0fab07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab3e58320dcca8c5756053852bfcc5423f3a0d401e361949136f5711586dbb04a04180fd35e9aef4cd62af512484e8fdde6242ad448b94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a97f366db7db30a613689e8c3724bd00a0392c13ea800d1e545836b91f3758dec9467df3e6b5d825f6d3edef49ca4f2d79ed5bce1ef264;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89361373d6190c6a9c86ba1c4206237244e02e84944d679b80275ca9deb245902776961285e18fd29e4ea325a9f058d68db0611a5ed2d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c26481def2c455463083ce07d659d9ba2077bb663dd9d9d02e2e58e115d41eebd7e6c7cb88a360bb9f18cd727359c5b5b0e02391fafb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb10b7a5aa868a9f4e37194b9401729b7eabe49ea15b976931305ed0b1fbb01774c9de97e19775390a142c57486a8996849b085e5f647b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a05bc899232f1b516ba16b60a5500f9dfe838c5b77e6afafd6eeb39fb4a697f2e7e41abc1d3093b45c077991c89f06ae843f666c868c03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4c8bceb0dae604203ce2420663dc1e65e758fceb2ce7e6c6149546049a208e593ec359a295bcc8d10266257a2511b8ec79546ead1efd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55958451c8df46e72d901e7e814417326cba4d974f2d163503f221351faaecfe68fc292dd91f9e98aa7f187f71c53a58f9ef0dc50f8d95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee3fbf46f47c8603af86f4bd07a14f8ff6561c4c18b0a608428ff93448392d3161eded9f49eb376ba01ce13c5326c918509eb9f6cb229a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb9a9db63719bf02b8e767767064287a0c3d0ce5d8ecdfba5839c4c1f3ba3dcda98717fe339d00505bb76840a77d75f6490c43d1c41c6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb72e9ddfdd361cab7237c9b6c44800c9684be3bf977897efacc558270535608bcd809f61ddaf8a441a26d417c3b7116dbbff8ba869d75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11198201520201ba3a6a7fb733272a724b025f7c3fdaf7048f18dad9d334a69dfbd032571bdbe383165569796637375258bf0ea68f4ecf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e226423367f34b3644af0dc8dc2e7a881af672c80235ce01e62e652b5e48050ea626c80a553cb21d3ac1795921761fba80d50996c2e2e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8685efb6048971ea1735aacc62fe3df2e1bf3664af8918cfe4e4b6ab1f715b1e7701980c3744467472183adf9c71fbd0e53f479e0b089;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173868657f2823c0105b1975fe061634ec5e7520350def79e891171e0f086d35e31642f56dcd28ef988bd24ee7801ba1cd92fae41589105;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1448ebc8a253eed832ebfef2dc1213b92d4b433b93252ad75b10673269df1eb388a5181a0bef903d177d91b547c25fa4c93718dbd0ae5cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f6f322655fe7c733f6eabd731084eb09ed4e31944f47a867d805fce3311b1392db126cb915646c936003af702bd34d9c5c5cb88adcea7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cc3169c6d0043c675b8bab67709b5e40dd1a47dad77b0a06bb89af46cc0fe8f3ae88c1ff5de477aec9b6cb3f81c448527bf4010c316f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e33d7185d70a12ba303b7cf30d3d0719140b6c952670fd7748831e07f8786f2085fe527725ab9f65f12d8ca66629a0ff90210ad11e3340;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1974406ab777f94761c4658211fea5848b013341d789f3f1649518bbb7d8b0602143c0c341d83cddadb538ac0d79b8fa2e0e432c58156a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc40f5c457afd2029a55296015da53876617ed3b899ab4e948ac75db69d2728848494eaf3bd91c74db3d330edf283c6805c40fc287d52f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcb242b8d1873c5509fe388db52b778846881f4bb0014296c4cad2a637c381acd80fe002490399f216995da81d20692a035a29e4d02ece;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173754c3c6ca033536416abb5bf71c9b36e3222d218d844d6bf22a3d914892c5e90e1a8aeb9ae3289d1913bafe800becfc9bc3ba37fda40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f5583ed99154ebd03beb0117e80c5e000f549265d11106fde64eb4eb4cd98c3e2192ecadc8f90915e1b0dd8018c107142ce4896576676;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c8f76504d390073b1956ca13c7244cf16493e24ec1cd3e97ac0f9c70e1d0b7f91f744bfed7edae83bcd1e235e6861050f4cf8a3a809bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b812c1fea32408e67b8f353b59beacdf68e88afcd762272c15161bffd9e772058fa1359231ba4ecb132e971ed28494a4bd4a451d8af24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23ecb015ab36f9212d5c2601be81da6b0f2c5e4e6cd30fbf508cebcf38dd7a0b015880df36b2f1cf77de327cd57e9274af2cfc9f3a74a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hefe7432a4f9bf961e9939e272e4a85ac0441ad9c09feeadcf7172efa38d5ebc22203c77625162cd288001283ac4b9a87f0875df07edf57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a80c3ae1ef76e46381e1841da9e4be1bfcec4920fb374b11ea04603ffd1d86cb5a17486d547319b07f77eee1b3f3938b267b4462b7c29a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdf6b16a88a90a5751c5494835615c01d61ba8208bddd5b70e868d651db50fc5f8c939dcec53315693987988826a2280992fa95842871;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac3f54ed535c6330905e4bd03600ff9abe04782f4150284d17d609a7462c25c926db9cef43724b97f8b98d7fc7f796077df97986048bf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc97e66a8bcf72c5d2b240d10c4f670f15981c223958c6214fb951b86542737deb1e9ad76bca33392a0d4f105b7ba3d5cfae4cf731a2fc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1581e9bfe329a16f4eada8fe181b171723203174fc17f30073b7b7de66b79b953da867c8844a4ea34ff7b8e4df4b7bd36d8fbbdb83a3383;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a939a77aa3396d2bd88fc9959dbbb5e6a713682a5d77ac4efeae50e6b7c6ae2d36eb97f4d91027304262c40b25384ea22b309027eb6b66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f841fab8a840d5ffe50545f1d02325ca51795643a0d9ea14ff61c0a1673a2324be7af741bb682e064abc73252f545d11e89d3a05bf7f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc20ab879d144f1bb84edb12d6a05c24da7429c2e0e3b3dd59e5cba6c303527e762b7ec211c6392f96f38c0e3aac0f35306e16e2db8d6a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h669b1c977bc139cd7dae163f539122ecb72c0a7908dd4b991959a9331c5327f6ac958ae71c5b44c74240d54acbec95fef8cbf150c45364;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h37384ddd0bc8a4eece40ef853698e850d2b9e916cef3a5db185b49a6c1ffc1b0f9b8cb9ffe2d0434182b12a66606c1d25730f86f11a042;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196a6e6bdf4f90fafd6f4e65d6877ebd6f9d4ae3b3b3ac31ee59d527d93d670ad443ecc24e7a4934182ba64e8c3d0b1df4565b5618b24d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ac3260210e108eb01b01ef299ab9e919db770929357f24cef290042e0e293c58a32df7b98a54ddfc371c7378d56b9212687876da88a87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed72b5b32feea00e54a5ef272bc0d5895f2f1dee282156c4a044d3cf29003b9e2502a5f8f47b430082d4413b9d09e0502082937f068090;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc88bd4ab435fa964ed046d44f18f92dcc33aa62fa5397ad0ff7baee25ffab5ca7ca18ea2ed5a4ea1c0bc6ab1ebfa1b6d56e00bd73e730;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c88a4f23088298f6139a9e3c42e7ea3b0b4d0c3484db2f92592b533a4b404dca5e169e7aa54b5890d2b895a080d4fbaf83c2f49a81d7a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc428b5276334fb04ea65ff83cc399d45e755c7389e3bac32b000c809ca39ad82632e5d7deb56a1593d71c254ee2a9c9223bef5e3bc49f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b3d287eb9d59e6720343122f5c66539007c9873b5a78e484dffcdecca4f6f6ecd58d958a46a35c3c73676a51c48862f81d3b6c699f412;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29340e0818963e7c9b04f29ea100e229fdde581ecdcf1b546d7b2184c826e18ce1a513f002e8cfd1bdd7862655477251b9c019d20309ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d40a2ca81b5c49c80b682886a3d459c4ba403cd661cfe93e0b9e626c36ae4b27fe69eaa6ed5a5d693003bee606d4f819f0816d0e283fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6b7e674dfd88359f8eff68f70e164dd4dcd78b943778e6fb26120f9908c76046f581ea886bb79a6b8346bdddaf5bebaab30e5cf2b5c2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197497f9f9e7137137d374377f8fcae71e62608cf28f0b4b78b6230a0b39a9e9004c371d7fa102ff1dcbdbcb81006b6f177013eb6475938;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8e44ccde078af83668999601320bd4b6c8b42349784e908777508e95456aac7f21524eec9a43cd204e0922c1f737daaf3fbe99280ecab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c7db0370369f974fb4b223bb2815a3c5217f954e82a8f6b86d6fdc4d0d70aecd69c87350e3f49248cbe449da7f88f2044fcfe012f9b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eb671219c47f1d54b5b5d49863f204cbcba7b041064fa0d922c902ba925e80a9bf5057441f60fc2755cd46b8336634ffd6e5a0ad34c82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a094bb2a85e58316ab2cbc0eeed0da34e81e53cb5f4646acf676fcfc8ae8fbf29cee6ffd854fc9c2feb3b860c98ab51c10494b5e00969;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9525ec39087c971d32a777a44b6e479dc48126d343fde4716d84527ea118933252e460721121850dae4ac11412cd7fd99869fe4f93100;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a459b99551bf79b4c0ed8c78e627b92cd65cf44bf9e98b8adf1567ebf12db8e8ac25ee9bd65ac22cc8a1eaa98a143301182eb28291eb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a9ff64172adc497fce4d22aae7e50f02814b60abbb1358da807f48cd5021ae440d81bed48ae4e1a8a9f309d69e7785b1f6b071626ac18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dd8a817e46e5c1645b1cf9683cb91900e963d07b4469baffab6bfb0235624d9852d26245461f8be5537a4060a465e49f974ca10b21a31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134e06a3c0d1eaf790597fba9c065a07c3c3f173e61ec0c1dbd6b1c4dff34c27ddfcadabcc6826a3e62db18fe36cc0b2fbebd1e064ee315;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c5856e1291b911793820cca31b6885655040ee234114cfeff54ece3a50bd422b030fae8d6bec932d93fad8f7de3ab7d38b2b3cf7244c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3189449685a86cb52943f71ae571a94848ffad8aea2ef880fb82d714cc22ed2179cebedd7e6da1591df505bf6f8d48fbf1b90a30fb53d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haddef68435f0c1928e4be7ff44467c22eff17763b2628f84592c6bf72b7edf03161f845c8a10badd4a29f9aa6f70bfd8edcf881dea7b4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10dddb7f93a910c1bcf334ec69bf7ec336aca514e6bacfde6a123279bdd5b0c9a7855672efb61fdc5098829a8231ffc96041491cba9ebed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c27affe715437954626e6ac9ef9225feba8bbeab0327e9c996e7f475711c601d8e439fb0ae2ebf4cf5e63e9e36c1980087c0f76348fcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1934b95c359c7761c8bcf15d04e19c0528695a3080d7206f0ccb7bbb087fe908b8816a609429978a6342eacb5c8565e9bbd3470398f09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff318ef4db36504a9928f27a69932315c450498fd8f11dd62275283d54d0d3dbbaa5687389311fe682eb220d9565166a688a96aff4df87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2bf53755aa1bfcbc8ccb5700024033fbb3801da7187e8952538f872a429a336ba618ebde96712faba613a6ff78127ec38e63a2aa39644;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha146a584b490df4ef8f5de28a90cb7e5d2b977480149dbabc3c9ca081ed30862614d62048d0fdfc8d97797b713f687a8824a49c61b6c54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1981622ea2b9b67960eff31054e4fb57389813ae212de806ca97264a7c9c5f3b62fa911d62b876610f2c1ac5c8e6dfb8f354fef1e72bc7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d43ffd1f7b956130c9e8095561bc056ffb381e4d1c4dc0b444b5acd54aa73109eb848199c7dd5d2b556c8a5c80116a6c18e7c70148554;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1858a0a5c163ffc848a0d487807020b19d0895841a96e5673e132c757e8dd19cf44f27edd01395ad035eacb33fe485d6645863d841175ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117603d6d5477d3437033143291ee0c57f01e25d49fd6ed3513b1a9e635dc2c9527743f222c607acc5938c136a14490bd772af7d47554f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176055bb346e6dc488491961881ea4aa7a52ddedbe441223fe3b0eca70cca0cb52327289f3898056576c3fcab2fb74c31c146f7a748ed3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea1e0c10bd6b48c61e2392ee7224dc2ea23f45f5b9c25d897c859751203fdb448fbf0c12281988d389ea401c73cd478c0a38b796b7c478;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75fb683e429cad2562efcd020c1e1032e96c09f1f8f4d380d4a68f87c31326fd174a3caa5b80f04c99d457f169ce9a9d9dd220770be204;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c96c1ea309391cbd032bd308bdb34fd6bf32eb7c7144588b1b61c6a8a83ad4cfdf5924c02e206e246ca43cbc3a1a0727d9c72c7ab04b3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153f215152490014d05b230e3e673036e91a1b5aa5b82f975d55a00e8c6b79fea6ac421f9d0098d042931ee62052de4330d4980a91f3d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4fff04b9c7271dc60ba4752bd9942cb1b39601b8f11945ebcae49e87ff9dd8cbd03406b9a720081ec172467fb15d0b53848e493740908;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdac589ab1014ae2b9bbc58389e25c277ed737b4e3e96009c794714b35316e374218983eae6661e602ae4f0c410aa5efb5303bb20fe6ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdd62172f982dcf24b635e203df6656c436dfe2fc532d61c1b63e5ed281798387a4fef680d8f72866ed36f86365fabbd02cdba7657e8dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1534ce8f0774e40b5ff3676a20b30880d3f970ef4c770cc0208ce3fc3b9eb31c6013ed9e6c9849df5fcbd1f6f80adede021276e69de2cae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0f0aaec60fd0a551597f9d225ec9e34be5aa63d97ab81f28086648317d69be2a3b408a001247a79bae92b3d2c2ab1fa2ffee5d046354;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9ec5a8537a6b1df698def53d3e011039c68bc99427fed5296a33c6e1efb4c0f93e25ebc158440d48e584bd387455325b21915bbe8956d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4270e5377d24a30504eacf5ab0b0d24a5887357e877ca7d58028a765e47142903120363144e1b50fe3b17426159facd47c600316074b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf43a86dc515b6250c44712e3dc2e2fe80966afd1965f7fe21a3335e17bf0739d688761c05f874883f5d1b973ccb4025d774349dd726db1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d07900516f21a3fe5a6163447728ab8bc9dd17382a60ef957ea5f374497ab55ea408daa3f2a05e70b3c17c979eb2e70aec12a36d585ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e652f6a1ef0af035fae4107a64fd889b0a86c6099b8974b2686f1ee99bcf2f8db3fc27e544f074aa9d762ec20e911384dc2897302810da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bc3c45aaa169bb8c7e03295a20bcbc365d101fa293843f4ebf888c273ca54b7f72f4998dade2aa0b8063e3f89529d643e40d2f261545a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe2ec9db086e4d69086a0d68ada318ae5a59af6bb16fef6ee2bb2ff476e21f8dfb1ceb01e8efca474f44f4942b5f52b57b0202bd18da22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b5cccc5ae64b57f5bd1c754262fecd9fdf12a61104cbcf6fa010a1bac74c4ff049371b196bb3483f57e29b3e28ca682a6c2e0353dd1e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134b8216be5aaeee50e75d5380833b848541ef632c006555ffed1a74887094a7c1aa22e463111b884d7b08797bbe28a857cdb752a7386fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e916744113ab8366d127233f28b84126777221f94e9198c6ed0fd626d7bf53267af43ba6f3c35075d49e5ae9001bad4d6dfc550d20db1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4573aba1e0d936838614746c5f3b5486bca5a44712aa4f392218de1fd64202c32384bf189e6a24c819d7e24aab750b2f11bcd1ed2b5193;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4fc0cef657c78cc8024b0cf3499ff4824584a1b7da1f112b882fc6daef8b42b12592614c97b71143e2dd9536ea4e6faceddacd5977b8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6f44320efbd4d6e1c123772928b1b3d2ae718fcf7d815f2dec86b7b15b1a13ce7ec1c1812d6997d2e1d3d8fd9774db907109a87f61c8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a86828de5ebdc316f1c74f47365cd4b38f5a440d5828dc49e2cea364527d9a413a47d24dba5be13717489ab9239248e767efd0ea4de8d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f875cb1ad09c9d6036a30edf0c7f092cccec97216ae5605f203f753db322ee6377af21da2133e40dca42e5e3b2e72ecf67d97b2535ca0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152c8aa3a418fbcb4f757f9c9fa3f653c48107a473b57f8d627fd8188dbea582d945b6f2fbcd5ea602ebf6c1182386834cb00def093e931;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1169dca6b7dc4e51479611e125f5d887fd01b75a6a0131d39c7e4065b96078ed3b52e24ee98779fb4d331199bff5034e09aff14cb002b24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8a3274132a9e32cfdce0f8ff928d52bc84622ccde63afd8159223bb1657c471787bd241d7f8c5ec64470d71c2b2f2c9a546f86c33fc40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3183d1b5d2507f937ad785909d0fe05ebd12692387225a602632e934e0020b76ff50eecfd3d6968a67e96988f017c28b1b633f10c9484;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2cf45afd80347d8d5d77747674a0304d91c3010062cc1553e5d6d0ecd8d5d76c8a7f8839f445a5e8b73a7db5db5489a1e292877a948b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144b4ad653a98b6e2656fcb459efd41c5ae13691d3c553ede6756c16f9318a57dd9b96735ad81ed7e6404c50bb32a17a017f8d68318f62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6ec2e5aac8419beff211b4c6ce2fc8a856e01956e2f3956cf2effc7c950cad271109c7ed7a1946a820bc22da6a0bd9f42bac5c4c571d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11683e1d2c4092104d3bec25f956caebff576fa55f549eb5b2590a0c9267574b7892a186c49e25ce87a1ce7e2b25a5ef7d413e5ae8d7500;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9899eda95149ff3ddb3d6ae7926648cfc47278bbde2a894f370dc2e993b85816dc933e62068df00744dd1880afdbba862a73eecc234bae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8caab570eb3ffe2aca8fecfe2c1e5e750c056f3d8f491ced8012980ddc38556197cc829d688230db6b8e093fa9c239eff8b74d285e8fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd676a899266f7b8de5efc25da5765f0d9c4f8bae5122edc1adf264614639c6e7fbcea3deb69811b461739b95f125923a2964bf2e66071;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c1ad771b1ffff5d68450b19ab06412b82e7fa17d729c10ec7885c712fd3d919cb250d15f62d1f676f97a54014f5af703e41064875475d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf720e3f6621865b2c6408c0c51e958259d87e15e11ec70fd89251becba00d6261ea52e3e9578a9e81e7e122d6846dbaee3c03c50801371;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee08c0b9c3fd9596db92bbcb01e961cb41e97a4703cdef491624c405438bfda763d1f80d8e3670d2b11cc8af5ae6be8418a12b77faf2ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha17058063cf53d289be9ab03dfba059f1c80f9f270d41cbf9c3f7e0f80a8d574696b17625a8b24f8d5f66744ee28718f56fdd6b2f37933;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbe706cf13c75da4747566a1b2d5f76add0e95443e6497a28e3a294c5419d48593408f5fe933d298f60f13b4c214dc9de5c77c46a1aa61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df619f332f703d8f5c45e882f2e977f7163a82bffd9cc51882ffaf31d036e6d6eea3300d76e64007c495ed18ec990ed35f083a6652ab7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151fcb8412f683b2e497149c6f675ccdf4e395c26bef56f1e7ca215b403f368852166178c0e8039e3bdf14f4701c16dc2da3b7bbdee0819;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3673b5849b74e5fd0e4e9b53e4406bdf4e11f029b79b377c3637466c77e925f11a01cb50e189242f143e382b037a4be7d77902a24cb0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a161d807f539396d8ee0547cb4819a9e221a4abfdba262e5252c6efba8a0ee15e470e42f0457031030a0d97f948d50b8c53f9320c1f13b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16bf02438f6d52eda65563c11711bd43b0702677c70243547a2e81fbf6b1a9584022d3dd3c6e317f63758301a367d943de20da50e96fff0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afa5e1599cf1664759cd4f2e3ac1a2e711004057b6c14bcfe69a29701d357518d29b76ada383b5e7e794256bf69fd924238cf98ee13528;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a8f5ae69d8689aed48e9a2248ec7ed4209030efe0f56d26c75326e6e4538238da4d4f2a15f2aeff3e9873fe9f27b9c4d48f49da289650;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f71b8efe701da457b88d1fa4c899e3b71eaf4f5b964f40977d1f1437012db457fc41389501f436786049b010fdfad89f5a44aa3f30a34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2000a1ff5e2863135a3d85ed9c96a9b50e662a46a9372291674d0df060f44e718fe6b508a2b0c8494d2352e652959d4defc8f21cc447bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168b6a7335b6930874c26ca652af2572dc109ea72cecc9ccb9c740164c118edec65823c149d28b7527fd71995d3fa9525e55d4cdc870f69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eea7c3b9d4087f74ee9285ab3ef9bd7306b332d5e339f5a157e6d011db2d0d185b9e527dc8e6e49096f2093355b150d90f20def14235cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h456b62136113231df6d88d0ffcb40b081c0e84af7a5acc3275c368fc830e80e756b3780b40661a8403d42fc2046bad1a1d2076076cf234;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4661661d8f3528de47c8c97fe017b520b1147ef92e58e4804449f57370566859fb298de01ddfc124dd28e1d052f66721f5a9ea236524ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c58fef0a877c52136117d5a2bbf4c9b27336c4483e39eeb8c757100ea1fc547c242c9857d778664241e5eb09a5df64b7856ac57c24ecf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bc0d5aab6f834b304068f08af7733ea2fc881feee671bfd315f120f40d201204c5067cb218c8c3fa8d2082070880cc05bd16acfbb17db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112cd027d360cfdc5e148f942e0631dfb3fcf0d793690074200ca8534e54be607171d5c736b82990d9a49eed1bff63f580715662fd1e79b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189e3462741c2a81d2af50a2eca0ad6b2aa04c6893e2682691fa3a8fba74bcdea25d9dfb85ea634489c7336accf51879d969ee69a6cd43f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16589bf73e089ae1e7948e9e500aa18299e2972b46fa8c720ffde7312567b8d2fd03fb63f23f8f3c94ad45eb0c74109a3f00cdc8989fa77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9af2f5b0dcabf67d91114ccc1b9aa74d3305e3649d5157753904724598f5601449c4ce3c11c095ad27e4356c630e3ef2ae144c5323c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5ee2a48df7262252d00c03367a80ecbd14e2d7e9a8c8966f325bd0ec6e5d29161a624c944b500df016ba8bf810a4adc033c405b479286;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb0541ddb48f82d1b6442c5df882034b0875defaeb56c3774ceae7e97d7a06f1ec309c3dffaa869753737db2148290a1a8e5d3dba3e9e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff2b2e7ebaf7ec6eaad605508025bfcc67471964599afa325ed8d9a8c388b4705944928b8e4d63e17ef04d15cf3f545f6e80da2b2c6447;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha07d058c0a48866ccfb020701436a9a350222e7cc99923e77499d026b33b1361827be54d756352e6dfc17e483780108164c8662bd5a960;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132855579bd5bf415d5bc71aafe2533fe2ca632dfe396bd39be4284dfd71f15c0aee26e242319521cace66a15867f2279b9b5f0c03768d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dcc6dd5aa658767144ca34956791385c934ded397156a52a2cf9b44821931ada9582801bc3920f193497bec1b175916564a4a20a264e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19651c724be74c05139eef4352a4c2c96ab365b464b9fb532c1a90e5b36f233febdbde1e15d8871525c1eb16f62a13a626db73cd31baa0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9eb79dd510a08fc4d2b2c942d09a5d993f4c66c2e3466c52a0315a7ab735073e3e9273eeffabdf12afe5aa214d596570fc62e3404d7121;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e352ebe195b09dd6bb31701e4a1156f6957375b619a9addbe2b13b237f6a2204df5cb6d62b2e918dcd30f64852341889a3a3f8c2966c39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce518b8d9e6f25eac140ba20ea0090dde82eef1a2fcb0b6e13f517c59594e36e11f154900ef2a771842aa5e8a1a2b80f08d2f87559e524;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23a96c04dfd093ac6c53098fc30c1a282aeacf6b6f8dcfd263696766d841473231beb71d2338efe13753c535b9fc4061010032eb2fbef8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a91d60c13e6034c742bd9e0a0df7da639df7e54bff4855cf165302035eb7ee579cdeb51b571945d8556b1233713545ee374555d5500d5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8d0d3ad9ceb9df6d6154fc7ed817ba13223e346f7e7ed2e9cf1f20d52978e339dc2e75493217ae6a52680809bc1cfba40a7c0788d6ac1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175dd6d29caa24be761345dcb14b60464bbc035075d900a821e9f4f79d21449d981c4e5871244fcaac2b3e30371b46b6264720cd425c028;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d3dfe4cc2eef11b41be003bdc8b0783339bfd0f2d17a5974d9f2acd4e24eda0d3d02b1189f9bfa397014ea3cf61439568830e2f79a1e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8192b97c58173d5c08d199c3c4907cfabbab5d58ecc105e951f0434f1a38a6be1285a3387f1b22ee0209a0b3d059ae94df8d7bce5c537;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d2ddc8b98525b9df94a18a5265708d1e976fc01c23f5b0f1fdd2e0c8f730c492bb703faa5a8c57ccbbb1bebd0199abe73ecd73004758;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1751ae9393491f97fcd1fd3b001d6d7ccde013c5d46c621ae8fc17759e6a3b744208f40f6f59deb81c627d9147735ce3b4a1c1f40e275c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88d72678b43d37001cec9348a5d7a5531840b03890a6b0eafb2b55b0c586fc05f3ae6071efa0fd7300a7ee9c5642f599db54ffe528c7a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1393c5525f242553db5ec5f68cbfb74f701cfea5d0a15580d604c9a59f0af6604c9883ab3f5aea5368e9076569f6460740af5cfe8bbe1e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d430f5e0dc3c41c15b3413f1752df7ca7716fc2fa31e7c778ccca4929d9e43f0d57962065e86969f6e2640d0699885f00549d3e99d396;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10501f16ab5383addefecc48532a63eb15e47220b1e1052897d729db8bc9d3000eb7928c9ac9e41b77e3423fe391e0a306096e58ff5ac54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf26dba49a1f1643e1b1f4ff379848411fc118c24159ecd5cd5e15ad7168aedaf3d747452368b85a52e024465fe5f09150756b81a952e4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162fccfa4a9a9020a18cc1d93904f38aed6aa1f52f526f601d90acea8bb9c7a207a1002ffd83cf80c1b5a39af0fbf7585faaa75b578c8ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b799d1ee4259c9a6e65b28ae4b1446a2177c5a7e7f947c8f25ea24d49b295abbbb9026ea2bf39724c1655646f57f0a9ecdfd4ef205f5f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0267fd02a5305aa9a60a5abdfca7f4edfe3934e161c3dd9f4671a524285f2e17c278b97b0bc825546889fa0dc669529cdec9d457b1fc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ce36136c98270e19ca42c1f88fe2b7e2890dcb874ff6209d3ae93c5e823e8d59907cffd032ff84bfe66216f97306f482bdf181531c929;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bec21c4618aca1a4e10dcf018605734400eb79d96c0648674875bd6aed9743288ddde11bf92d19b0e8c678225114332b5d6657b340965;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c1aaab87ce5be138dc202a6ef32b5a0adef1b5ff2e9dadd1489aa64682f01d970ae21258c7f276d24cdead8ed7843c75627b99a88d93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125c6d05676294d81b03f1e0c724a289fee81bf99d47aa90afb6665b0eb33c5e040f943dd13c4e8420c80a2ddbbde70442bea435b6059e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h443fceec47f03392845d161419ac3536a0263aeaf582e6dfcb3abecaad10e47fb44021f76f05d81506ea1db6377fdfe31ac7e00b33cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff1f6c9f15f7aeebba2e9228b010ffbd551618927c4f9c692d7080d8470135c9478d2361a981fdfb0d1ee3f6201fc52cf2d29f120bde6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a224f67abfed51cedca11a911ce729ad5d92c7a70dc75eec7ea91bfb7f983a76c5093b31dad830a277d70058a10a8c680bd46c0dc171a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b9c1dc82d59c3c8ac6f3d67970980a29871668aa8122c6784cbca052faa4932fc2ef125b3f860854d811378a44532ab3c334fd119eb64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99d49467d77f2b3fcb84068fbc24859cbf27ed07e52233152989f7be347785e07c9f1989efe3bb1e13d1b034dde37bb740476221bec85c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9fe3c5bffa3bcc9032fd7b8163e77a842f0d095abc4f46744fc91a428eae65c497f22ef2f8574b54afe0ce319b4a075894d415526825e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8e544b0b18db1bfff5509a57d76cf50c4143d22c92d0ec7bf0f61e6ea354dce6e81116c2a1ed37a137bb7db81cc5ec08d3e7c45d7f01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9329c9bad71bcf5138f5482daa2049f89a26496104e0a3dafcf2f7dddaee5f330d71afed8e0d171aea971d18c89f52901e950c8dd24d7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9229527b3fdec58176803d50b4f7410087bc47651647f0738a42b22d1e13a2a876846b737b3b53d554d404472e692693c3dae474bf30c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc2d35101b56100a989e4e449c606fc4038a0eb0f8acf54d130deb3ca4dbd2d3b0c01d2eadc533dd59e0b37708d9e00267f9a8f76c31e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137b362bff43d454691c065d35eaf825e76b063b61cf16f3eeb594d173ee51adbd3fafc8be3adea8dbb6f86464996c7cd3719744ae73dde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h570d29a8dc0acd089cd5cbebb425ecd8e918b2dcd7a218c537d25af1278538524d90aa4bad619ca1c22ec314dbb9f71ad2a9da6599de3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba10699e2abec94a1f3abb095d27cbf6c3158e690fb1020a3d594afa2f063715df5f33b4829926359f442c812802d02dd67cd2eb52b6e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17513789e052e4db1d79af127e3441a06f96b24eaec6db1af56fddfd99606fd44b6e0586f613f73d41222c337e579fcdab40ac92fa1d517;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78eb6261243bea782fc39869b73d22da46c0238ac9ac776a1a40c30e5c38ce22e786cca7515d20798f6ffe17ce0117d8fdf904c786c600;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hede6683024e72a7254442802a0d3006ef31a2a10aa84495728f3d83c08880acd52212364c1774cd9610a3d1a552ddd1cfe90178de9b82a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca48b3799d4e2562683d69200cf47e9abc8849121653ef2d268f43a1299d51318b120c9299906c86bd9fe4feaf29dcb03db8f48abfd191;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h939bc9255e5d14630229beb41cf960bb61343b4519ec3cc4225fac070d40c69a18a204a602afcf685fa10e6b9469b3e35e8c898783679d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38da6ca891e513f06ea29121fc69aa7997c95a17a2586437b96c572c43a06a20e7a1c014c57757644ff5017c2f10b6d738d135e44bf4f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e5ddaaea9842011c4e7533e71e79700f7c5078e8613c9e258a219bed631c4ae65656670440fee656ecbafbad70a4aa9129a2fe317d4eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98b146d998c9feaa4dc52f56c72666f33b9b5dd3bb34a0e964e5086040d1cda66417d7882f159f11d2e5ada091b00b2189c6b85be43ea4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcee8d738215731c512d242b19bdc70a77eb2dc3072943b4cfc92012fdc4120348722db46a2979df22ff865c4bd8da6f248285e973da82c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4ed7c7753e1e51abd81f8424fbdf49810cb75e76a17070258117f94cf92bc54756a8cbf517807b88f354d1c675e3e29256a7beb9edaac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbf493b553f2ac55fa9befabef91f6e8a20b3075c674979bf39ff8bce1df30bb860059b9061830f901eb9168555a51f8f59336acd45cd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccfae9de598972f823b0e764808cb3343a84143554322655978707e75afb4539632ff5ef2631b483f19df8fb63a7234980b09842ff1a65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd15f0d5052d838ae1e3229f610226aef67f649f8c85a70e962ef2834bf07daea4ea8d4a48ed95c9c577e363d5ed120e36f38be79765f23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb08c1f3f711ae31bbd1fc30f0115965e5957e3b8518efe70816f6c21101e0407e5908db42bd239dc89dba116e263dd72704d0c9a921145;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a09deb6d3e52186b9353b832fa4028ac42ae0d6d945cd4cc4d0173bff480acbafc6312729129e385ba89c70d6d34a9dab6e117875523d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b243bd7790675e53e882c3a68ed83e5a074d11c52b346d163baf0204bfaee7b7bcc515f4853b6895d7767e87f974779f85ed51c8ad8e88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191634e02f360652ccc9b9df4d0047f791531beda35c453b58b836612eede8e0c38bec608f180ec8fbc375509becbae7d9d564ae56b0155;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbdcc4d0d53a2fdafa791d29d49952773e727091272dd10557e61ea93ddafab9f57610dec388f0af0022b981f85a9744dae9f2fb9d17a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ef351a338ec8781e9a99dd9d689dae514fc749e7c84b2c7e7198d46eafd1ffa04c05779a34a3df918536eed22e20163777f3f313b68d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0699346343a190ad7e5fee71572c1afae97f405432a4b09b1c9293ce9c2defaf13ff03c57d5a8e42a890440be19afec1255e20cb292a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc16737a613eea0e588ad55ed349982a318170d55c345cab372dcd4d5519c5fd6e13fcf9dbec3fe5686d89234928e75dd14bc8adf760417;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b901587bf1ac15835bc4b7365324e7c876bea631662c14ca49e295d9bd766513da9f418e763ba98dbf0ae264d0353f9a9a4ed4cd6c08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162b4f87cb2c5105818f7636277942bad53dc1b8e671b7b196389696f35e5678e020078a084afa591083a2e32e8c5964525086492bfc850;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h355b7281f909becb09ab421bc5692624fb7246f588e7d8a85a10f084abe7d3f63084f89374b28a3d3d656103a15f1c7bc4e8ba0a9ed93b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5c474fa986689c1f9b2f2ef50df099931210a13a034bf0b6866679b5b528f25fdac596c5c1b6e890a48c0003a046d0d73738e90ff0966;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3f0d712c9fabb311974207661d6f06c041be586856a53efc2932680b9eebd679469c2e041a74461805ee8c20e3b5fac30b5c241bad04f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f1abb00d7728c3e130b07b6e169494675911327d16dc4d970293efefa7bf102766ecfb79e1b8023da0d670b2ec9f3d80301f39cec7e38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a147d0ca617a8088d8b596ada0e7ef15500844e805ed1979ccfba53e381421fd914977e56344cf74a2ae5c36e75ff8b5d91ea685b8da3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f350fe9f0a771e49c3f8c9bbcd616dcdc80d95e3ec157f70d64a3647af6329c836efdb87f1406eefdacdd66a62d871edaa8a434c70922a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c8d17ace31541bb2b89262d542c610fbae107492a4474dd9c937d3b384d7215d5e1de26d105d1a700c10de19ddddf0839e3e1a6b564e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c0e6a636129b450f66f04b2982d4b416a5c860a6bdb005dc407c7ced853af5d94237140117793f2bb0ee861ee323ea6dddcafb0eb7b12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd42de15de3e044dcb48aa41fcaaa5e6539ca7398af8fb140d67489e4fd25ffed48d145f543881cc8656c17ecb6626414e9e6f7ea0ae09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e56a941419bff986bd647ca6fa8de6e87b9e986697509cf432adda7be183a2e40f54da62189d488156b9d23e88ce8b11c211f09f12d1d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99bcec2b10541c75bc8b2cae62cfffb99fa87a40b2bb5771ac4f2b880b93610b4d8bdcb3fe9148e8436e48431eca71a566d43f48e92ac5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d66dcdd1604c710e553096914b5486374233d74a662777f26cd131e7891cae850b58d6a5640b08064a5691240c635d0c287d73e2e5791;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dfb02c479d2dec8577b500a789913191ec0a6cffc675e34a0b071f1be06e317164494f68e33837c9d08d66366d0b3963e0df2101614ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7c1284daf18b4981d361b8e059ea2a38f3349514b230b0b492b2a4b1544d6dcd21693db6dd85f5a0607a5f27289361f52275cb99be805;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc743ce1f79406b745bbe1854e9524f92ab5a81e8e9d3d495bd66a6235864f4eaa851dfed8f2ee6138c5fcdf4056cdaa395784ba3ff3716;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6ec7f885db8eef9f5bbc33fc6e80d9e3eafb3e064bb7610aa24356d2fee187d80bc40d72bba503f38bdb5517c9a8fce945ce0a958799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85a35508ed016472c78715d67171fc5c24643ebba971af2e0a5f63b2c05850feb22907a64805d123eaa6a0665bf3df31e0cf29174fde9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82bde7a87816c50ca71a3e505e581bf0ffdb97e17d6610828f3d8acde4cf6f7f441edacbee4ed23f9e0c198de55287d75f0a081e6f290d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162665bd7229fdc05ef316875b77032b36b50abde111a77225a072b0d5f316bf569a2191b79bf6e841b2c438f3ed0a5660425e9e3236045;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96499f0831172688e7482433ce6a26ad0b137d58b769dec6c10c2b8474de1b595231d7d438025a712efff11478880bf0a114e23b0776b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2970e6d6b938c46593fff258384c3cc12356c4338b77865d9db565e5d6241c098478eabe71cf75788f75dcce546c669a3d4c01ded3b2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba514cfa499f95c2cccb26f8d568f9daa7e3d2c2729547cf0ace70451152cf275a60b56a7e4a0bb1915f357af2c714c62411ab2b41dd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15fb7891d69181f5cffc07870b56c52ddf005af6d303418eeb5dcaf50cd681d06593311b6ed90003cb3df58d1bbf9f738ceca6174304fef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9c6af2e3ec2d3ae4a214d2233608cddf18d5fa3a34036aace86171caf921e4d8d8d36b115e9527273afe135e1f1b68af419577fde1b0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9c54a93aa37caa9508dab6b0222798c3ccd0fa5737ca06171743803d65af2387714885b5290e54e13b2538566d72fe3185d02a8bbdd1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6cda6d9ff2e43b80d0dc3da780a4df1a57aa005e769289c2b454d0bc864ae10bdeb299c8493516a0fbce112937cfea706b88ae26d90e1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8272c9d491ba65e264431d3ab3b2a244cb359344d9a3aa7ea8f96d33614cb11b4403bb93d4c27a678f7e32a3bb72c241eafc10ef7ccca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e5db6f4f0375735db5d72c3b11d1c78ecb548615a764a78aeed83f59d39866372cd8be025e0cc733ff2b499084f50d7f49e13d5e65fb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1f8ea8b6dac84aeb9cdbe6b4dd468ba1cd5b68ed2e7382adc012ea98df4b93c2b29ac9ef04513993b98d4ab615768072f4476021697ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1433ec07b770a23e4f3246bb9a57756c77f071b5ce4938752a5c9debf80f584e0d148b0071ad2f488cc529fc4dcfadf96c413ca429ccd5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180d01a189f52dea8d9b4a099d2f5cd0723182041cea5d1decfe73303af358220c37063ce2eadf236c9c7bd93cf31b9c3fcb3a94da32d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a01225acfd570ec8240bc37a3789e8d9c949881e138ab720f19b01e6cb87b1059154a0633977910d87e753569c70683afe6cf25596b39c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa72e06112c1a1d5b186be431971a157259253562e65def3e131cee4d426b1467fd9d51e78233e48214810c61653dd785c8a31c5556e8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1965ee13dbf42e889547cc7a94bac9bd00beec4cc38b68c476da6afb5d3766803d789cf4e47fc994f4be21f90959ec3916fffa77103131d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67c94c9a5b1086396f9a792f68ec2447d703a653ad60f947877d31d1bde1166843adb9deaaa8c0baf21328caa3d32f3e3dd3cb30af3053;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h493834af0429e2d2e6fdc7f5bef2e1fa95778978ffeb05e6febbefb2f2c0736126b510c3e52705784bf10676334959320243b320fbe7bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1702d175ee860fde30301d7571bff359120de1746bf19363a71dc46df987f9534a9d0d24483d3499a9de3ad55062648cd33ef5ec0867ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187702d6aa4997f4c0db6f335203c54f1ae35be0e2e98ebc928a25d8f52408b96090883aeca6d7e1a417d2dbdc962d75f865a37e40e92d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h882ca9439e1ed0f3f1919f1302c1630f65fb0125ebd0967642b741ad67213ef7c49a2b8f9d04ade7536c4e1c59f70611b3ef53e58b4286;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e1cdb3338997d19444bccdb9f825031ef3d2db6edc55a456492416eeba14c6a7784d86b25d05a8e55f5e09bdfb4834859dbe2cc8098f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d42153a1f87425399dc42b23f4c3161f436eba358c4b0d16f6611e0778db9c1b247e2b498012f3d106451dedc53fa8bfe5ed0b8fd29b84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bf1c118ba2ede8d079a9c9c5ac7a04f061795e844265bc4c5f996d7b37bdfed37c2d7802703f751e36b22dcc3187bede106d6ec077d32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31754df60d621a619dfe68036399322369aa66c3472498a8c284eb9b5a92a8f150604d7968743968d0f7051edf0f4c577317c65d55ac62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd4c4aa663d8aca73e7fcdca85d28a7cdacbe05c7d3d23e491fe9f15832d00d9043f1001ee490053ab2a5189f1afdc315bada573453bf2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20b0c000a5441370ba7831a82950497df9a8b750ce25f61e512772bb853c4698329b825a5e92baf13970f3995a5439d82e626b4b1952c3;
        #1
        $finish();
    end
endmodule
