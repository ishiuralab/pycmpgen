module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    compressor_CLA512_64 compressor_CLA512_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
        src32 <= 512'h0;
        src33 <= 512'h0;
        src34 <= 512'h0;
        src35 <= 512'h0;
        src36 <= 512'h0;
        src37 <= 512'h0;
        src38 <= 512'h0;
        src39 <= 512'h0;
        src40 <= 512'h0;
        src41 <= 512'h0;
        src42 <= 512'h0;
        src43 <= 512'h0;
        src44 <= 512'h0;
        src45 <= 512'h0;
        src46 <= 512'h0;
        src47 <= 512'h0;
        src48 <= 512'h0;
        src49 <= 512'h0;
        src50 <= 512'h0;
        src51 <= 512'h0;
        src52 <= 512'h0;
        src53 <= 512'h0;
        src54 <= 512'h0;
        src55 <= 512'h0;
        src56 <= 512'h0;
        src57 <= 512'h0;
        src58 <= 512'h0;
        src59 <= 512'h0;
        src60 <= 512'h0;
        src61 <= 512'h0;
        src62 <= 512'h0;
        src63 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA512_64(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    input [511:0]src32,
    input [511:0]src33,
    input [511:0]src34,
    input [511:0]src35,
    input [511:0]src36,
    input [511:0]src37,
    input [511:0]src38,
    input [511:0]src39,
    input [511:0]src40,
    input [511:0]src41,
    input [511:0]src42,
    input [511:0]src43,
    input [511:0]src44,
    input [511:0]src45,
    input [511:0]src46,
    input [511:0]src47,
    input [511:0]src48,
    input [511:0]src49,
    input [511:0]src50,
    input [511:0]src51,
    input [511:0]src52,
    input [511:0]src53,
    input [511:0]src54,
    input [511:0]src55,
    input [511:0]src56,
    input [511:0]src57,
    input [511:0]src58,
    input [511:0]src59,
    input [511:0]src60,
    input [511:0]src61,
    input [511:0]src62,
    input [511:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [0:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], 1'h0, comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      input wire [511:0] src32,
      input wire [511:0] src33,
      input wire [511:0] src34,
      input wire [511:0] src35,
      input wire [511:0] src36,
      input wire [511:0] src37,
      input wire [511:0] src38,
      input wire [511:0] src39,
      input wire [511:0] src40,
      input wire [511:0] src41,
      input wire [511:0] src42,
      input wire [511:0] src43,
      input wire [511:0] src44,
      input wire [511:0] src45,
      input wire [511:0] src46,
      input wire [511:0] src47,
      input wire [511:0] src48,
      input wire [511:0] src49,
      input wire [511:0] src50,
      input wire [511:0] src51,
      input wire [511:0] src52,
      input wire [511:0] src53,
      input wire [511:0] src54,
      input wire [511:0] src55,
      input wire [511:0] src56,
      input wire [511:0] src57,
      input wire [511:0] src58,
      input wire [511:0] src59,
      input wire [511:0] src60,
      input wire [511:0] src61,
      input wire [511:0] src62,
      input wire [511:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [0:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [511:0] stage0_32;
   wire [511:0] stage0_33;
   wire [511:0] stage0_34;
   wire [511:0] stage0_35;
   wire [511:0] stage0_36;
   wire [511:0] stage0_37;
   wire [511:0] stage0_38;
   wire [511:0] stage0_39;
   wire [511:0] stage0_40;
   wire [511:0] stage0_41;
   wire [511:0] stage0_42;
   wire [511:0] stage0_43;
   wire [511:0] stage0_44;
   wire [511:0] stage0_45;
   wire [511:0] stage0_46;
   wire [511:0] stage0_47;
   wire [511:0] stage0_48;
   wire [511:0] stage0_49;
   wire [511:0] stage0_50;
   wire [511:0] stage0_51;
   wire [511:0] stage0_52;
   wire [511:0] stage0_53;
   wire [511:0] stage0_54;
   wire [511:0] stage0_55;
   wire [511:0] stage0_56;
   wire [511:0] stage0_57;
   wire [511:0] stage0_58;
   wire [511:0] stage0_59;
   wire [511:0] stage0_60;
   wire [511:0] stage0_61;
   wire [511:0] stage0_62;
   wire [511:0] stage0_63;
   wire [118:0] stage1_0;
   wire [168:0] stage1_1;
   wire [220:0] stage1_2;
   wire [321:0] stage1_3;
   wire [250:0] stage1_4;
   wire [216:0] stage1_5;
   wire [179:0] stage1_6;
   wire [339:0] stage1_7;
   wire [238:0] stage1_8;
   wire [362:0] stage1_9;
   wire [152:0] stage1_10;
   wire [317:0] stage1_11;
   wire [218:0] stage1_12;
   wire [184:0] stage1_13;
   wire [255:0] stage1_14;
   wire [257:0] stage1_15;
   wire [223:0] stage1_16;
   wire [217:0] stage1_17;
   wire [241:0] stage1_18;
   wire [218:0] stage1_19;
   wire [243:0] stage1_20;
   wire [204:0] stage1_21;
   wire [200:0] stage1_22;
   wire [298:0] stage1_23;
   wire [234:0] stage1_24;
   wire [210:0] stage1_25;
   wire [188:0] stage1_26;
   wire [211:0] stage1_27;
   wire [248:0] stage1_28;
   wire [220:0] stage1_29;
   wire [232:0] stage1_30;
   wire [211:0] stage1_31;
   wire [414:0] stage1_32;
   wire [209:0] stage1_33;
   wire [267:0] stage1_34;
   wire [190:0] stage1_35;
   wire [330:0] stage1_36;
   wire [302:0] stage1_37;
   wire [276:0] stage1_38;
   wire [196:0] stage1_39;
   wire [229:0] stage1_40;
   wire [276:0] stage1_41;
   wire [228:0] stage1_42;
   wire [243:0] stage1_43;
   wire [268:0] stage1_44;
   wire [188:0] stage1_45;
   wire [299:0] stage1_46;
   wire [277:0] stage1_47;
   wire [210:0] stage1_48;
   wire [241:0] stage1_49;
   wire [216:0] stage1_50;
   wire [226:0] stage1_51;
   wire [303:0] stage1_52;
   wire [186:0] stage1_53;
   wire [262:0] stage1_54;
   wire [225:0] stage1_55;
   wire [256:0] stage1_56;
   wire [179:0] stage1_57;
   wire [242:0] stage1_58;
   wire [293:0] stage1_59;
   wire [199:0] stage1_60;
   wire [216:0] stage1_61;
   wire [372:0] stage1_62;
   wire [294:0] stage1_63;
   wire [111:0] stage1_64;
   wire [56:0] stage1_65;
   wire [33:0] stage2_0;
   wire [38:0] stage2_1;
   wire [72:0] stage2_2;
   wire [253:0] stage2_3;
   wire [92:0] stage2_4;
   wire [111:0] stage2_5;
   wire [120:0] stage2_6;
   wire [96:0] stage2_7;
   wire [172:0] stage2_8;
   wire [104:0] stage2_9;
   wire [133:0] stage2_10;
   wire [135:0] stage2_11;
   wire [127:0] stage2_12;
   wire [71:0] stage2_13;
   wire [114:0] stage2_14;
   wire [114:0] stage2_15;
   wire [109:0] stage2_16;
   wire [89:0] stage2_17;
   wire [161:0] stage2_18;
   wire [93:0] stage2_19;
   wire [87:0] stage2_20;
   wire [111:0] stage2_21;
   wire [109:0] stage2_22;
   wire [97:0] stage2_23;
   wire [84:0] stage2_24;
   wire [122:0] stage2_25;
   wire [130:0] stage2_26;
   wire [85:0] stage2_27;
   wire [79:0] stage2_28;
   wire [111:0] stage2_29;
   wire [99:0] stage2_30;
   wire [127:0] stage2_31;
   wire [117:0] stage2_32;
   wire [108:0] stage2_33;
   wire [127:0] stage2_34;
   wire [117:0] stage2_35;
   wire [119:0] stage2_36;
   wire [113:0] stage2_37;
   wire [99:0] stage2_38;
   wire [107:0] stage2_39;
   wire [139:0] stage2_40;
   wire [122:0] stage2_41;
   wire [81:0] stage2_42;
   wire [110:0] stage2_43;
   wire [137:0] stage2_44;
   wire [131:0] stage2_45;
   wire [92:0] stage2_46;
   wire [107:0] stage2_47;
   wire [153:0] stage2_48;
   wire [115:0] stage2_49;
   wire [152:0] stage2_50;
   wire [87:0] stage2_51;
   wire [127:0] stage2_52;
   wire [96:0] stage2_53;
   wire [123:0] stage2_54;
   wire [110:0] stage2_55;
   wire [131:0] stage2_56;
   wire [78:0] stage2_57;
   wire [84:0] stage2_58;
   wire [139:0] stage2_59;
   wire [110:0] stage2_60;
   wire [101:0] stage2_61;
   wire [144:0] stage2_62;
   wire [112:0] stage2_63;
   wire [101:0] stage2_64;
   wire [67:0] stage2_65;
   wire [53:0] stage2_66;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [14:0] stage3_2;
   wire [51:0] stage3_3;
   wire [59:0] stage3_4;
   wire [54:0] stage3_5;
   wire [66:0] stage3_6;
   wire [54:0] stage3_7;
   wire [46:0] stage3_8;
   wire [52:0] stage3_9;
   wire [67:0] stage3_10;
   wire [60:0] stage3_11;
   wire [80:0] stage3_12;
   wire [46:0] stage3_13;
   wire [34:0] stage3_14;
   wire [50:0] stage3_15;
   wire [58:0] stage3_16;
   wire [43:0] stage3_17;
   wire [63:0] stage3_18;
   wire [45:0] stage3_19;
   wire [57:0] stage3_20;
   wire [62:0] stage3_21;
   wire [49:0] stage3_22;
   wire [48:0] stage3_23;
   wire [34:0] stage3_24;
   wire [51:0] stage3_25;
   wire [51:0] stage3_26;
   wire [41:0] stage3_27;
   wire [69:0] stage3_28;
   wire [58:0] stage3_29;
   wire [38:0] stage3_30;
   wire [41:0] stage3_31;
   wire [55:0] stage3_32;
   wire [62:0] stage3_33;
   wire [44:0] stage3_34;
   wire [56:0] stage3_35;
   wire [55:0] stage3_36;
   wire [34:0] stage3_37;
   wire [68:0] stage3_38;
   wire [59:0] stage3_39;
   wire [45:0] stage3_40;
   wire [56:0] stage3_41;
   wire [53:0] stage3_42;
   wire [59:0] stage3_43;
   wire [84:0] stage3_44;
   wire [39:0] stage3_45;
   wire [48:0] stage3_46;
   wire [73:0] stage3_47;
   wire [36:0] stage3_48;
   wire [64:0] stage3_49;
   wire [63:0] stage3_50;
   wire [53:0] stage3_51;
   wire [55:0] stage3_52;
   wire [52:0] stage3_53;
   wire [62:0] stage3_54;
   wire [46:0] stage3_55;
   wire [38:0] stage3_56;
   wire [52:0] stage3_57;
   wire [48:0] stage3_58;
   wire [45:0] stage3_59;
   wire [52:0] stage3_60;
   wire [56:0] stage3_61;
   wire [40:0] stage3_62;
   wire [71:0] stage3_63;
   wire [50:0] stage3_64;
   wire [32:0] stage3_65;
   wire [53:0] stage3_66;
   wire [14:0] stage3_67;
   wire [4:0] stage3_68;
   wire [5:0] stage4_0;
   wire [6:0] stage4_1;
   wire [8:0] stage4_2;
   wire [21:0] stage4_3;
   wire [24:0] stage4_4;
   wire [46:0] stage4_5;
   wire [20:0] stage4_6;
   wire [39:0] stage4_7;
   wire [34:0] stage4_8;
   wire [13:0] stage4_9;
   wire [28:0] stage4_10;
   wire [33:0] stage4_11;
   wire [19:0] stage4_12;
   wire [27:0] stage4_13;
   wire [29:0] stage4_14;
   wire [22:0] stage4_15;
   wire [32:0] stage4_16;
   wire [22:0] stage4_17;
   wire [31:0] stage4_18;
   wire [19:0] stage4_19;
   wire [21:0] stage4_20;
   wire [26:0] stage4_21;
   wire [20:0] stage4_22;
   wire [23:0] stage4_23;
   wire [23:0] stage4_24;
   wire [19:0] stage4_25;
   wire [20:0] stage4_26;
   wire [20:0] stage4_27;
   wire [31:0] stage4_28;
   wire [23:0] stage4_29;
   wire [25:0] stage4_30;
   wire [16:0] stage4_31;
   wire [23:0] stage4_32;
   wire [33:0] stage4_33;
   wire [29:0] stage4_34;
   wire [23:0] stage4_35;
   wire [37:0] stage4_36;
   wire [15:0] stage4_37;
   wire [26:0] stage4_38;
   wire [22:0] stage4_39;
   wire [28:0] stage4_40;
   wire [23:0] stage4_41;
   wire [28:0] stage4_42;
   wire [22:0] stage4_43;
   wire [39:0] stage4_44;
   wire [25:0] stage4_45;
   wire [24:0] stage4_46;
   wire [25:0] stage4_47;
   wire [21:0] stage4_48;
   wire [27:0] stage4_49;
   wire [23:0] stage4_50;
   wire [26:0] stage4_51;
   wire [22:0] stage4_52;
   wire [28:0] stage4_53;
   wire [30:0] stage4_54;
   wire [28:0] stage4_55;
   wire [28:0] stage4_56;
   wire [24:0] stage4_57;
   wire [15:0] stage4_58;
   wire [15:0] stage4_59;
   wire [24:0] stage4_60;
   wire [28:0] stage4_61;
   wire [23:0] stage4_62;
   wire [17:0] stage4_63;
   wire [26:0] stage4_64;
   wire [22:0] stage4_65;
   wire [14:0] stage4_66;
   wire [16:0] stage4_67;
   wire [11:0] stage4_68;
   wire [2:0] stage4_69;
   wire [0:0] stage4_70;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [2:0] stage5_2;
   wire [7:0] stage5_3;
   wire [8:0] stage5_4;
   wire [20:0] stage5_5;
   wire [13:0] stage5_6;
   wire [10:0] stage5_7;
   wire [15:0] stage5_8;
   wire [12:0] stage5_9;
   wire [9:0] stage5_10;
   wire [19:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [14:0] stage5_14;
   wire [15:0] stage5_15;
   wire [13:0] stage5_16;
   wire [7:0] stage5_17;
   wire [13:0] stage5_18;
   wire [13:0] stage5_19;
   wire [7:0] stage5_20;
   wire [10:0] stage5_21;
   wire [14:0] stage5_22;
   wire [11:0] stage5_23;
   wire [8:0] stage5_24;
   wire [12:0] stage5_25;
   wire [16:0] stage5_26;
   wire [8:0] stage5_27;
   wire [11:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [11:0] stage5_31;
   wire [14:0] stage5_32;
   wire [8:0] stage5_33;
   wire [20:0] stage5_34;
   wire [8:0] stage5_35;
   wire [18:0] stage5_36;
   wire [10:0] stage5_37;
   wire [6:0] stage5_38;
   wire [10:0] stage5_39;
   wire [19:0] stage5_40;
   wire [8:0] stage5_41;
   wire [19:0] stage5_42;
   wire [7:0] stage5_43;
   wire [25:0] stage5_44;
   wire [9:0] stage5_45;
   wire [10:0] stage5_46;
   wire [12:0] stage5_47;
   wire [17:0] stage5_48;
   wire [16:0] stage5_49;
   wire [9:0] stage5_50;
   wire [9:0] stage5_51;
   wire [12:0] stage5_52;
   wire [11:0] stage5_53;
   wire [16:0] stage5_54;
   wire [17:0] stage5_55;
   wire [12:0] stage5_56;
   wire [8:0] stage5_57;
   wire [23:0] stage5_58;
   wire [5:0] stage5_59;
   wire [13:0] stage5_60;
   wire [9:0] stage5_61;
   wire [7:0] stage5_62;
   wire [10:0] stage5_63;
   wire [19:0] stage5_64;
   wire [5:0] stage5_65;
   wire [12:0] stage5_66;
   wire [7:0] stage5_67;
   wire [11:0] stage5_68;
   wire [2:0] stage5_69;
   wire [3:0] stage5_70;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [2:0] stage6_2;
   wire [3:0] stage6_3;
   wire [2:0] stage6_4;
   wire [6:0] stage6_5;
   wire [5:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [7:0] stage6_9;
   wire [4:0] stage6_10;
   wire [5:0] stage6_11;
   wire [7:0] stage6_12;
   wire [4:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [11:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [8:0] stage6_25;
   wire [4:0] stage6_26;
   wire [4:0] stage6_27;
   wire [3:0] stage6_28;
   wire [5:0] stage6_29;
   wire [7:0] stage6_30;
   wire [2:0] stage6_31;
   wire [5:0] stage6_32;
   wire [7:0] stage6_33;
   wire [5:0] stage6_34;
   wire [4:0] stage6_35;
   wire [7:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [4:0] stage6_39;
   wire [9:0] stage6_40;
   wire [10:0] stage6_41;
   wire [3:0] stage6_42;
   wire [4:0] stage6_43;
   wire [7:0] stage6_44;
   wire [6:0] stage6_45;
   wire [6:0] stage6_46;
   wire [3:0] stage6_47;
   wire [5:0] stage6_48;
   wire [9:0] stage6_49;
   wire [4:0] stage6_50;
   wire [4:0] stage6_51;
   wire [7:0] stage6_52;
   wire [3:0] stage6_53;
   wire [5:0] stage6_54;
   wire [5:0] stage6_55;
   wire [6:0] stage6_56;
   wire [6:0] stage6_57;
   wire [6:0] stage6_58;
   wire [4:0] stage6_59;
   wire [6:0] stage6_60;
   wire [5:0] stage6_61;
   wire [4:0] stage6_62;
   wire [2:0] stage6_63;
   wire [5:0] stage6_64;
   wire [9:0] stage6_65;
   wire [2:0] stage6_66;
   wire [4:0] stage6_67;
   wire [9:0] stage6_68;
   wire [2:0] stage6_69;
   wire [1:0] stage6_70;
   wire [1:0] stage6_71;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [2:0] stage7_2;
   wire [3:0] stage7_3;
   wire [0:0] stage7_4;
   wire [4:0] stage7_5;
   wire [1:0] stage7_6;
   wire [6:0] stage7_7;
   wire [0:0] stage7_8;
   wire [4:0] stage7_9;
   wire [3:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [6:0] stage7_13;
   wire [2:0] stage7_14;
   wire [1:0] stage7_15;
   wire [6:0] stage7_16;
   wire [2:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [0:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [6:0] stage7_23;
   wire [2:0] stage7_24;
   wire [5:0] stage7_25;
   wire [6:0] stage7_26;
   wire [0:0] stage7_27;
   wire [1:0] stage7_28;
   wire [2:0] stage7_29;
   wire [3:0] stage7_30;
   wire [1:0] stage7_31;
   wire [2:0] stage7_32;
   wire [2:0] stage7_33;
   wire [5:0] stage7_34;
   wire [6:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [2:0] stage7_38;
   wire [3:0] stage7_39;
   wire [1:0] stage7_40;
   wire [5:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [6:0] stage7_45;
   wire [6:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [5:0] stage7_49;
   wire [2:0] stage7_50;
   wire [5:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [4:0] stage7_54;
   wire [1:0] stage7_55;
   wire [5:0] stage7_56;
   wire [2:0] stage7_57;
   wire [1:0] stage7_58;
   wire [2:0] stage7_59;
   wire [4:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [4:0] stage7_63;
   wire [2:0] stage7_64;
   wire [11:0] stage7_65;
   wire [0:0] stage7_66;
   wire [0:0] stage7_67;
   wire [3:0] stage7_68;
   wire [2:0] stage7_69;
   wire [2:0] stage7_70;
   wire [2:0] stage7_71;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [1:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [0:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_2[7]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[8]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[9]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[10]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[11]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[12]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[13]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[14]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[15]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[16]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[17]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[18]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[19]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[20]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[21]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[22]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[23]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[24]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[25]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[26]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[27]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[28]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[29]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[30]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[31]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[32]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[33]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[34]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[35]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[36]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_2[37]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_2[38]},
      {stage0_3[31]},
      {stage1_4[31],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_2[39]},
      {stage0_3[32]},
      {stage1_4[32],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_2[40]},
      {stage0_3[33]},
      {stage1_4[33],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_2[41]},
      {stage0_3[34]},
      {stage1_4[34],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_2[42]},
      {stage0_3[35]},
      {stage1_4[35],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_2[43]},
      {stage0_3[36]},
      {stage1_4[36],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_2[44]},
      {stage0_3[37]},
      {stage1_4[37],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc1163_5 gpc45 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_2[45]},
      {stage0_3[38]},
      {stage1_4[38],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc1163_5 gpc46 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_2[46]},
      {stage0_3[39]},
      {stage1_4[39],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc1163_5 gpc47 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_2[47]},
      {stage0_3[40]},
      {stage1_4[40],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc1163_5 gpc48 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_2[48]},
      {stage0_3[41]},
      {stage1_4[41],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc1163_5 gpc49 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_2[49]},
      {stage0_3[42]},
      {stage1_4[42],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc1163_5 gpc50 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_2[50]},
      {stage0_3[43]},
      {stage1_4[43],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc1163_5 gpc51 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_2[51]},
      {stage0_3[44]},
      {stage1_4[44],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc1163_5 gpc52 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_2[52]},
      {stage0_3[45]},
      {stage1_4[45],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc1163_5 gpc53 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_2[53]},
      {stage0_3[46]},
      {stage1_4[46],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc1163_5 gpc54 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_2[54]},
      {stage0_3[47]},
      {stage1_4[47],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc1163_5 gpc55 (
      {stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_2[55]},
      {stage0_3[48]},
      {stage1_4[48],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc1163_5 gpc56 (
      {stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_2[56]},
      {stage0_3[49]},
      {stage1_4[49],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[50],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[51],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[52],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[53],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc615_5 gpc61 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_1[307]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[54],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc615_5 gpc62 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_1[308]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[55],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc615_5 gpc63 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_1[309]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[56],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc615_5 gpc64 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_1[310]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[57],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc615_5 gpc65 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247]},
      {stage0_1[311]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[58],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc615_5 gpc66 (
      {stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_1[312]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[59],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc615_5 gpc67 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_1[313]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[60],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc615_5 gpc68 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_1[314]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[61],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc615_5 gpc69 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_1[315]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[62],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc615_5 gpc70 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_1[316]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[63],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc615_5 gpc71 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277]},
      {stage0_1[317]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[64],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc615_5 gpc72 (
      {stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_1[318]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[65],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc615_5 gpc73 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_1[319]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[66],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc615_5 gpc74 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_1[320]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[67],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc615_5 gpc75 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_1[321]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[68],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc615_5 gpc76 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_1[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[69],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc615_5 gpc77 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307]},
      {stage0_1[323]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[70],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc615_5 gpc78 (
      {stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_1[324]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[71],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc615_5 gpc79 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_1[325]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[72],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc615_5 gpc80 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_1[326]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[73],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc615_5 gpc81 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_1[327]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[74],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc615_5 gpc82 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_1[328]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[75],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc615_5 gpc83 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337]},
      {stage0_1[329]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[76],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc615_5 gpc84 (
      {stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_1[330]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[77],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc615_5 gpc85 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_1[331]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[78],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc615_5 gpc86 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_1[332]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[79],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc615_5 gpc87 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_1[333]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[80],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc615_5 gpc88 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_1[334]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[81],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc615_5 gpc89 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367]},
      {stage0_1[335]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[82],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc615_5 gpc90 (
      {stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_1[336]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[83],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc615_5 gpc91 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_1[337]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[84],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc615_5 gpc92 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_1[338]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[85],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc615_5 gpc93 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_1[339]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[86],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc615_5 gpc94 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_1[340]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[87],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc615_5 gpc95 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397]},
      {stage0_1[341]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[88],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc615_5 gpc96 (
      {stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_1[342]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[89],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc615_5 gpc97 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_1[343]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[90],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc615_5 gpc98 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_1[344]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[91],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc615_5 gpc99 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_1[345]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[92],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc615_5 gpc100 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_1[346]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[93],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc615_5 gpc101 (
      {stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427]},
      {stage0_1[347]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[94],stage1_3[101],stage1_2[101],stage1_1[101],stage1_0[101]}
   );
   gpc615_5 gpc102 (
      {stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_1[348]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[95],stage1_3[102],stage1_2[102],stage1_1[102],stage1_0[102]}
   );
   gpc615_5 gpc103 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_1[349]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[96],stage1_3[103],stage1_2[103],stage1_1[103],stage1_0[103]}
   );
   gpc615_5 gpc104 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_1[350]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[97],stage1_3[104],stage1_2[104],stage1_1[104],stage1_0[104]}
   );
   gpc615_5 gpc105 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_1[351]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[98],stage1_3[105],stage1_2[105],stage1_1[105],stage1_0[105]}
   );
   gpc615_5 gpc106 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452]},
      {stage0_1[352]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[99],stage1_3[106],stage1_2[106],stage1_1[106],stage1_0[106]}
   );
   gpc615_5 gpc107 (
      {stage0_0[453], stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457]},
      {stage0_1[353]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[100],stage1_3[107],stage1_2[107],stage1_1[107],stage1_0[107]}
   );
   gpc615_5 gpc108 (
      {stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461], stage0_0[462]},
      {stage0_1[354]},
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage1_4[101],stage1_3[108],stage1_2[108],stage1_1[108],stage1_0[108]}
   );
   gpc615_5 gpc109 (
      {stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_1[355]},
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage1_4[102],stage1_3[109],stage1_2[109],stage1_1[109],stage1_0[109]}
   );
   gpc615_5 gpc110 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_1[356]},
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage1_4[103],stage1_3[110],stage1_2[110],stage1_1[110],stage1_0[110]}
   );
   gpc615_5 gpc111 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_1[357]},
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage1_4[104],stage1_3[111],stage1_2[111],stage1_1[111],stage1_0[111]}
   );
   gpc615_5 gpc112 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482]},
      {stage0_1[358]},
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage1_4[105],stage1_3[112],stage1_2[112],stage1_1[112],stage1_0[112]}
   );
   gpc615_5 gpc113 (
      {stage0_0[483], stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487]},
      {stage0_1[359]},
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage1_4[106],stage1_3[113],stage1_2[113],stage1_1[113],stage1_0[113]}
   );
   gpc615_5 gpc114 (
      {stage0_0[488], stage0_0[489], stage0_0[490], stage0_0[491], stage0_0[492]},
      {stage0_1[360]},
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage1_4[107],stage1_3[114],stage1_2[114],stage1_1[114],stage1_0[114]}
   );
   gpc615_5 gpc115 (
      {stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496], stage0_0[497]},
      {stage0_1[361]},
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage1_4[108],stage1_3[115],stage1_2[115],stage1_1[115],stage1_0[115]}
   );
   gpc615_5 gpc116 (
      {stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_1[362]},
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416]},
      {stage1_4[109],stage1_3[116],stage1_2[116],stage1_1[116],stage1_0[116]}
   );
   gpc615_5 gpc117 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507]},
      {stage0_1[363]},
      {stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage1_4[110],stage1_3[117],stage1_2[117],stage1_1[117],stage1_0[117]}
   );
   gpc615_5 gpc118 (
      {stage0_0[508], stage0_0[509], stage0_0[510], stage0_0[511], 1'b0},
      {stage0_1[364]},
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage1_4[111],stage1_3[118],stage1_2[118],stage1_1[118],stage1_0[118]}
   );
   gpc7_3 gpc119 (
      {stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc7_3 gpc120 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[0],stage1_4[112],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[1],stage1_4[113],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[2],stage1_4[114],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[3],stage1_4[115],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[4],stage1_4[116],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[5],stage1_4[117],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[6],stage1_4[118],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[7],stage1_4[119],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[8],stage1_4[120],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[9],stage1_4[121],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[10],stage1_4[122],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[11],stage1_4[123],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[12],stage1_4[124],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[13],stage1_4[125],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[14],stage1_4[126],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[15],stage1_4[127],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479], stage0_1[480]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[16],stage1_4[128],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc615_5 gpc138 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[17],stage1_4[129],stage1_3[138]}
   );
   gpc615_5 gpc139 (
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[18],stage1_4[130],stage1_3[139]}
   );
   gpc615_5 gpc140 (
      {stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[19],stage1_4[131],stage1_3[140]}
   );
   gpc615_5 gpc141 (
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[20],stage1_4[132],stage1_3[141]}
   );
   gpc615_5 gpc142 (
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[21],stage1_4[133],stage1_3[142]}
   );
   gpc615_5 gpc143 (
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181]},
      {stage0_4[5]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[5],stage1_5[22],stage1_4[134],stage1_3[143]}
   );
   gpc615_5 gpc144 (
      {stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage0_4[6]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[6],stage1_5[23],stage1_4[135],stage1_3[144]}
   );
   gpc615_5 gpc145 (
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191]},
      {stage0_4[7]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[7],stage1_5[24],stage1_4[136],stage1_3[145]}
   );
   gpc615_5 gpc146 (
      {stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage0_4[8]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[8],stage1_5[25],stage1_4[137],stage1_3[146]}
   );
   gpc615_5 gpc147 (
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage0_4[9]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[9],stage1_5[26],stage1_4[138],stage1_3[147]}
   );
   gpc615_5 gpc148 (
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage0_4[10]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[10],stage1_5[27],stage1_4[139],stage1_3[148]}
   );
   gpc615_5 gpc149 (
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211]},
      {stage0_4[11]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[11],stage1_5[28],stage1_4[140],stage1_3[149]}
   );
   gpc615_5 gpc150 (
      {stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage0_4[12]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[12],stage1_5[29],stage1_4[141],stage1_3[150]}
   );
   gpc615_5 gpc151 (
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221]},
      {stage0_4[13]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[13],stage1_5[30],stage1_4[142],stage1_3[151]}
   );
   gpc615_5 gpc152 (
      {stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage0_4[14]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[14],stage1_5[31],stage1_4[143],stage1_3[152]}
   );
   gpc615_5 gpc153 (
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage0_4[15]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[15],stage1_5[32],stage1_4[144],stage1_3[153]}
   );
   gpc615_5 gpc154 (
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage0_4[16]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[16],stage1_5[33],stage1_4[145],stage1_3[154]}
   );
   gpc615_5 gpc155 (
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241]},
      {stage0_4[17]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[17],stage1_5[34],stage1_4[146],stage1_3[155]}
   );
   gpc615_5 gpc156 (
      {stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage0_4[18]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[18],stage1_5[35],stage1_4[147],stage1_3[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251]},
      {stage0_4[19]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[19],stage1_5[36],stage1_4[148],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage0_4[20]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[20],stage1_5[37],stage1_4[149],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage0_4[21]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[21],stage1_5[38],stage1_4[150],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage0_4[22]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[22],stage1_5[39],stage1_4[151],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271]},
      {stage0_4[23]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[23],stage1_5[40],stage1_4[152],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage0_4[24]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[24],stage1_5[41],stage1_4[153],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281]},
      {stage0_4[25]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[25],stage1_5[42],stage1_4[154],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage0_4[26]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[26],stage1_5[43],stage1_4[155],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage0_4[27]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[27],stage1_5[44],stage1_4[156],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage0_4[28]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[28],stage1_5[45],stage1_4[157],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301]},
      {stage0_4[29]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[29],stage1_5[46],stage1_4[158],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage0_4[30]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[30],stage1_5[47],stage1_4[159],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311]},
      {stage0_4[31]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[31],stage1_5[48],stage1_4[160],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316]},
      {stage0_4[32]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[32],stage1_5[49],stage1_4[161],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage0_4[33]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[33],stage1_5[50],stage1_4[162],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage0_4[34]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[34],stage1_5[51],stage1_4[163],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331]},
      {stage0_4[35]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[35],stage1_5[52],stage1_4[164],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage0_4[36]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[36],stage1_5[53],stage1_4[165],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341]},
      {stage0_4[37]},
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage1_7[37],stage1_6[37],stage1_5[54],stage1_4[166],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346]},
      {stage0_4[38]},
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage1_7[38],stage1_6[38],stage1_5[55],stage1_4[167],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350], stage0_3[351]},
      {stage0_4[39]},
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage1_7[39],stage1_6[39],stage1_5[56],stage1_4[168],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage0_4[40]},
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage1_7[40],stage1_6[40],stage1_5[57],stage1_4[169],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361]},
      {stage0_4[41]},
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage1_7[41],stage1_6[41],stage1_5[58],stage1_4[170],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366]},
      {stage0_4[42]},
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage1_7[42],stage1_6[42],stage1_5[59],stage1_4[171],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370], stage0_3[371]},
      {stage0_4[43]},
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage1_7[43],stage1_6[43],stage1_5[60],stage1_4[172],stage1_3[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[44],stage1_6[44],stage1_5[61],stage1_4[173]}
   );
   gpc606_5 gpc183 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[45],stage1_6[45],stage1_5[62],stage1_4[174]}
   );
   gpc606_5 gpc184 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[46],stage1_6[46],stage1_5[63],stage1_4[175]}
   );
   gpc606_5 gpc185 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[47],stage1_6[47],stage1_5[64],stage1_4[176]}
   );
   gpc606_5 gpc186 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[48],stage1_6[48],stage1_5[65],stage1_4[177]}
   );
   gpc606_5 gpc187 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[49],stage1_6[49],stage1_5[66],stage1_4[178]}
   );
   gpc606_5 gpc188 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[50],stage1_6[50],stage1_5[67],stage1_4[179]}
   );
   gpc606_5 gpc189 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[51],stage1_6[51],stage1_5[68],stage1_4[180]}
   );
   gpc606_5 gpc190 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[52],stage1_6[52],stage1_5[69],stage1_4[181]}
   );
   gpc606_5 gpc191 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[53],stage1_6[53],stage1_5[70],stage1_4[182]}
   );
   gpc606_5 gpc192 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[54],stage1_6[54],stage1_5[71],stage1_4[183]}
   );
   gpc606_5 gpc193 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[55],stage1_6[55],stage1_5[72],stage1_4[184]}
   );
   gpc606_5 gpc194 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[56],stage1_6[56],stage1_5[73],stage1_4[185]}
   );
   gpc606_5 gpc195 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[57],stage1_6[57],stage1_5[74],stage1_4[186]}
   );
   gpc606_5 gpc196 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[58],stage1_6[58],stage1_5[75],stage1_4[187]}
   );
   gpc606_5 gpc197 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[59],stage1_6[59],stage1_5[76],stage1_4[188]}
   );
   gpc606_5 gpc198 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[60],stage1_6[60],stage1_5[77],stage1_4[189]}
   );
   gpc606_5 gpc199 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[61],stage1_6[61],stage1_5[78],stage1_4[190]}
   );
   gpc606_5 gpc200 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[62],stage1_6[62],stage1_5[79],stage1_4[191]}
   );
   gpc606_5 gpc201 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[63],stage1_6[63],stage1_5[80],stage1_4[192]}
   );
   gpc606_5 gpc202 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[64],stage1_6[64],stage1_5[81],stage1_4[193]}
   );
   gpc606_5 gpc203 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[65],stage1_6[65],stage1_5[82],stage1_4[194]}
   );
   gpc606_5 gpc204 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[66],stage1_6[66],stage1_5[83],stage1_4[195]}
   );
   gpc606_5 gpc205 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[67],stage1_6[67],stage1_5[84],stage1_4[196]}
   );
   gpc606_5 gpc206 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[68],stage1_6[68],stage1_5[85],stage1_4[197]}
   );
   gpc606_5 gpc207 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[69],stage1_6[69],stage1_5[86],stage1_4[198]}
   );
   gpc606_5 gpc208 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[70],stage1_6[70],stage1_5[87],stage1_4[199]}
   );
   gpc606_5 gpc209 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[71],stage1_6[71],stage1_5[88],stage1_4[200]}
   );
   gpc606_5 gpc210 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[72],stage1_6[72],stage1_5[89],stage1_4[201]}
   );
   gpc606_5 gpc211 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[73],stage1_6[73],stage1_5[90],stage1_4[202]}
   );
   gpc606_5 gpc212 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[74],stage1_6[74],stage1_5[91],stage1_4[203]}
   );
   gpc606_5 gpc213 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[75],stage1_6[75],stage1_5[92],stage1_4[204]}
   );
   gpc606_5 gpc214 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[76],stage1_6[76],stage1_5[93],stage1_4[205]}
   );
   gpc606_5 gpc215 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[77],stage1_6[77],stage1_5[94],stage1_4[206]}
   );
   gpc606_5 gpc216 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[78],stage1_6[78],stage1_5[95],stage1_4[207]}
   );
   gpc606_5 gpc217 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[79],stage1_6[79],stage1_5[96],stage1_4[208]}
   );
   gpc606_5 gpc218 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[80],stage1_6[80],stage1_5[97],stage1_4[209]}
   );
   gpc606_5 gpc219 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[81],stage1_6[81],stage1_5[98],stage1_4[210]}
   );
   gpc606_5 gpc220 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[82],stage1_6[82],stage1_5[99],stage1_4[211]}
   );
   gpc606_5 gpc221 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[83],stage1_6[83],stage1_5[100],stage1_4[212]}
   );
   gpc606_5 gpc222 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[84],stage1_6[84],stage1_5[101],stage1_4[213]}
   );
   gpc606_5 gpc223 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[85],stage1_6[85],stage1_5[102],stage1_4[214]}
   );
   gpc606_5 gpc224 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[86],stage1_6[86],stage1_5[103],stage1_4[215]}
   );
   gpc606_5 gpc225 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[87],stage1_6[87],stage1_5[104],stage1_4[216]}
   );
   gpc606_5 gpc226 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[88],stage1_6[88],stage1_5[105],stage1_4[217]}
   );
   gpc606_5 gpc227 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[89],stage1_6[89],stage1_5[106],stage1_4[218]}
   );
   gpc606_5 gpc228 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[90],stage1_6[90],stage1_5[107],stage1_4[219]}
   );
   gpc606_5 gpc229 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[91],stage1_6[91],stage1_5[108],stage1_4[220]}
   );
   gpc606_5 gpc230 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[92],stage1_6[92],stage1_5[109],stage1_4[221]}
   );
   gpc606_5 gpc231 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[93],stage1_6[93],stage1_5[110],stage1_4[222]}
   );
   gpc606_5 gpc232 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[94],stage1_6[94],stage1_5[111],stage1_4[223]}
   );
   gpc606_5 gpc233 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[95],stage1_6[95],stage1_5[112],stage1_4[224]}
   );
   gpc606_5 gpc234 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[96],stage1_6[96],stage1_5[113],stage1_4[225]}
   );
   gpc606_5 gpc235 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[97],stage1_6[97],stage1_5[114],stage1_4[226]}
   );
   gpc606_5 gpc236 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[98],stage1_6[98],stage1_5[115],stage1_4[227]}
   );
   gpc606_5 gpc237 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[99],stage1_6[99],stage1_5[116],stage1_4[228]}
   );
   gpc606_5 gpc238 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[100],stage1_6[100],stage1_5[117],stage1_4[229]}
   );
   gpc606_5 gpc239 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[101],stage1_6[101],stage1_5[118],stage1_4[230]}
   );
   gpc606_5 gpc240 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[102],stage1_6[102],stage1_5[119],stage1_4[231]}
   );
   gpc606_5 gpc241 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[103],stage1_6[103],stage1_5[120],stage1_4[232]}
   );
   gpc606_5 gpc242 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[104],stage1_6[104],stage1_5[121],stage1_4[233]}
   );
   gpc606_5 gpc243 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[105],stage1_6[105],stage1_5[122],stage1_4[234]}
   );
   gpc606_5 gpc244 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[106],stage1_6[106],stage1_5[123],stage1_4[235]}
   );
   gpc606_5 gpc245 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[107],stage1_6[107],stage1_5[124],stage1_4[236]}
   );
   gpc606_5 gpc246 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[108],stage1_6[108],stage1_5[125],stage1_4[237]}
   );
   gpc606_5 gpc247 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[109],stage1_6[109],stage1_5[126],stage1_4[238]}
   );
   gpc606_5 gpc248 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[110],stage1_6[110],stage1_5[127],stage1_4[239]}
   );
   gpc606_5 gpc249 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[111],stage1_6[111],stage1_5[128],stage1_4[240]}
   );
   gpc606_5 gpc250 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[112],stage1_6[112],stage1_5[129],stage1_4[241]}
   );
   gpc606_5 gpc251 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[113],stage1_6[113],stage1_5[130],stage1_4[242]}
   );
   gpc606_5 gpc252 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[114],stage1_6[114],stage1_5[131],stage1_4[243]}
   );
   gpc606_5 gpc253 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[115],stage1_6[115],stage1_5[132],stage1_4[244]}
   );
   gpc606_5 gpc254 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[116],stage1_6[116],stage1_5[133],stage1_4[245]}
   );
   gpc606_5 gpc255 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486], stage0_4[487]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[117],stage1_6[117],stage1_5[134],stage1_4[246]}
   );
   gpc606_5 gpc256 (
      {stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491], stage0_4[492], stage0_4[493]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[118],stage1_6[118],stage1_5[135],stage1_4[247]}
   );
   gpc606_5 gpc257 (
      {stage0_4[494], stage0_4[495], stage0_4[496], stage0_4[497], stage0_4[498], stage0_4[499]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[119],stage1_6[119],stage1_5[136],stage1_4[248]}
   );
   gpc606_5 gpc258 (
      {stage0_4[500], stage0_4[501], stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[120],stage1_6[120],stage1_5[137],stage1_4[249]}
   );
   gpc606_5 gpc259 (
      {stage0_4[506], stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage1_8[77],stage1_7[121],stage1_6[121],stage1_5[138],stage1_4[250]}
   );
   gpc606_5 gpc260 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[78],stage1_7[122],stage1_6[122],stage1_5[139]}
   );
   gpc606_5 gpc261 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[79],stage1_7[123],stage1_6[123],stage1_5[140]}
   );
   gpc606_5 gpc262 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[80],stage1_7[124],stage1_6[124],stage1_5[141]}
   );
   gpc606_5 gpc263 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[81],stage1_7[125],stage1_6[125],stage1_5[142]}
   );
   gpc606_5 gpc264 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[82],stage1_7[126],stage1_6[126],stage1_5[143]}
   );
   gpc606_5 gpc265 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[83],stage1_7[127],stage1_6[127],stage1_5[144]}
   );
   gpc606_5 gpc266 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[84],stage1_7[128],stage1_6[128],stage1_5[145]}
   );
   gpc606_5 gpc267 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[85],stage1_7[129],stage1_6[129],stage1_5[146]}
   );
   gpc606_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[86],stage1_7[130],stage1_6[130],stage1_5[147]}
   );
   gpc606_5 gpc269 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[87],stage1_7[131],stage1_6[131],stage1_5[148]}
   );
   gpc606_5 gpc270 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[88],stage1_7[132],stage1_6[132],stage1_5[149]}
   );
   gpc606_5 gpc271 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[89],stage1_7[133],stage1_6[133],stage1_5[150]}
   );
   gpc606_5 gpc272 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[90],stage1_7[134],stage1_6[134],stage1_5[151]}
   );
   gpc606_5 gpc273 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[91],stage1_7[135],stage1_6[135],stage1_5[152]}
   );
   gpc606_5 gpc274 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[92],stage1_7[136],stage1_6[136],stage1_5[153]}
   );
   gpc606_5 gpc275 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[93],stage1_7[137],stage1_6[137],stage1_5[154]}
   );
   gpc606_5 gpc276 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[94],stage1_7[138],stage1_6[138],stage1_5[155]}
   );
   gpc606_5 gpc277 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[95],stage1_7[139],stage1_6[139],stage1_5[156]}
   );
   gpc606_5 gpc278 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[96],stage1_7[140],stage1_6[140],stage1_5[157]}
   );
   gpc606_5 gpc279 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[97],stage1_7[141],stage1_6[141],stage1_5[158]}
   );
   gpc606_5 gpc280 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[98],stage1_7[142],stage1_6[142],stage1_5[159]}
   );
   gpc606_5 gpc281 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[99],stage1_7[143],stage1_6[143],stage1_5[160]}
   );
   gpc606_5 gpc282 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[100],stage1_7[144],stage1_6[144],stage1_5[161]}
   );
   gpc606_5 gpc283 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[101],stage1_7[145],stage1_6[145],stage1_5[162]}
   );
   gpc606_5 gpc284 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[102],stage1_7[146],stage1_6[146],stage1_5[163]}
   );
   gpc606_5 gpc285 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[103],stage1_7[147],stage1_6[147],stage1_5[164]}
   );
   gpc606_5 gpc286 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[104],stage1_7[148],stage1_6[148],stage1_5[165]}
   );
   gpc606_5 gpc287 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[105],stage1_7[149],stage1_6[149],stage1_5[166]}
   );
   gpc606_5 gpc288 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[106],stage1_7[150],stage1_6[150],stage1_5[167]}
   );
   gpc606_5 gpc289 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[107],stage1_7[151],stage1_6[151],stage1_5[168]}
   );
   gpc606_5 gpc290 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[108],stage1_7[152],stage1_6[152],stage1_5[169]}
   );
   gpc606_5 gpc291 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[109],stage1_7[153],stage1_6[153],stage1_5[170]}
   );
   gpc606_5 gpc292 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[110],stage1_7[154],stage1_6[154],stage1_5[171]}
   );
   gpc606_5 gpc293 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[111],stage1_7[155],stage1_6[155],stage1_5[172]}
   );
   gpc615_5 gpc294 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472]},
      {stage0_7[204]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[34],stage1_8[112],stage1_7[156],stage1_6[156]}
   );
   gpc615_5 gpc295 (
      {stage0_6[473], stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477]},
      {stage0_7[205]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[35],stage1_8[113],stage1_7[157],stage1_6[157]}
   );
   gpc615_5 gpc296 (
      {stage0_6[478], stage0_6[479], stage0_6[480], stage0_6[481], stage0_6[482]},
      {stage0_7[206]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[36],stage1_8[114],stage1_7[158],stage1_6[158]}
   );
   gpc615_5 gpc297 (
      {stage0_6[483], stage0_6[484], stage0_6[485], stage0_6[486], stage0_6[487]},
      {stage0_7[207]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[37],stage1_8[115],stage1_7[159],stage1_6[159]}
   );
   gpc615_5 gpc298 (
      {stage0_6[488], stage0_6[489], stage0_6[490], stage0_6[491], stage0_6[492]},
      {stage0_7[208]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[38],stage1_8[116],stage1_7[160],stage1_6[160]}
   );
   gpc615_5 gpc299 (
      {stage0_7[209], stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[39],stage1_8[117],stage1_7[161]}
   );
   gpc615_5 gpc300 (
      {stage0_7[214], stage0_7[215], stage0_7[216], stage0_7[217], stage0_7[218]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[40],stage1_8[118],stage1_7[162]}
   );
   gpc615_5 gpc301 (
      {stage0_7[219], stage0_7[220], stage0_7[221], stage0_7[222], stage0_7[223]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[41],stage1_8[119],stage1_7[163]}
   );
   gpc615_5 gpc302 (
      {stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227], stage0_7[228]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[42],stage1_8[120],stage1_7[164]}
   );
   gpc615_5 gpc303 (
      {stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[43],stage1_8[121],stage1_7[165]}
   );
   gpc615_5 gpc304 (
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[44],stage1_8[122],stage1_7[166]}
   );
   gpc615_5 gpc305 (
      {stage0_7[239], stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[45],stage1_8[123],stage1_7[167]}
   );
   gpc615_5 gpc306 (
      {stage0_7[244], stage0_7[245], stage0_7[246], stage0_7[247], stage0_7[248]},
      {stage0_8[37]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[12],stage1_9[46],stage1_8[124],stage1_7[168]}
   );
   gpc615_5 gpc307 (
      {stage0_7[249], stage0_7[250], stage0_7[251], stage0_7[252], stage0_7[253]},
      {stage0_8[38]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[13],stage1_9[47],stage1_8[125],stage1_7[169]}
   );
   gpc615_5 gpc308 (
      {stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257], stage0_7[258]},
      {stage0_8[39]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[14],stage1_9[48],stage1_8[126],stage1_7[170]}
   );
   gpc615_5 gpc309 (
      {stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage0_8[40]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[15],stage1_9[49],stage1_8[127],stage1_7[171]}
   );
   gpc615_5 gpc310 (
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268]},
      {stage0_8[41]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[16],stage1_9[50],stage1_8[128],stage1_7[172]}
   );
   gpc615_5 gpc311 (
      {stage0_7[269], stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273]},
      {stage0_8[42]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[17],stage1_9[51],stage1_8[129],stage1_7[173]}
   );
   gpc615_5 gpc312 (
      {stage0_7[274], stage0_7[275], stage0_7[276], stage0_7[277], stage0_7[278]},
      {stage0_8[43]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[18],stage1_9[52],stage1_8[130],stage1_7[174]}
   );
   gpc615_5 gpc313 (
      {stage0_7[279], stage0_7[280], stage0_7[281], stage0_7[282], stage0_7[283]},
      {stage0_8[44]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[19],stage1_9[53],stage1_8[131],stage1_7[175]}
   );
   gpc615_5 gpc314 (
      {stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287], stage0_7[288]},
      {stage0_8[45]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[20],stage1_9[54],stage1_8[132],stage1_7[176]}
   );
   gpc615_5 gpc315 (
      {stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage0_8[46]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[21],stage1_9[55],stage1_8[133],stage1_7[177]}
   );
   gpc615_5 gpc316 (
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298]},
      {stage0_8[47]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[22],stage1_9[56],stage1_8[134],stage1_7[178]}
   );
   gpc615_5 gpc317 (
      {stage0_7[299], stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303]},
      {stage0_8[48]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[23],stage1_9[57],stage1_8[135],stage1_7[179]}
   );
   gpc615_5 gpc318 (
      {stage0_7[304], stage0_7[305], stage0_7[306], stage0_7[307], stage0_7[308]},
      {stage0_8[49]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[24],stage1_9[58],stage1_8[136],stage1_7[180]}
   );
   gpc615_5 gpc319 (
      {stage0_7[309], stage0_7[310], stage0_7[311], stage0_7[312], stage0_7[313]},
      {stage0_8[50]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[25],stage1_9[59],stage1_8[137],stage1_7[181]}
   );
   gpc615_5 gpc320 (
      {stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317], stage0_7[318]},
      {stage0_8[51]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[26],stage1_9[60],stage1_8[138],stage1_7[182]}
   );
   gpc615_5 gpc321 (
      {stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage0_8[52]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[27],stage1_9[61],stage1_8[139],stage1_7[183]}
   );
   gpc615_5 gpc322 (
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328]},
      {stage0_8[53]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[28],stage1_9[62],stage1_8[140],stage1_7[184]}
   );
   gpc615_5 gpc323 (
      {stage0_7[329], stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333]},
      {stage0_8[54]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[29],stage1_9[63],stage1_8[141],stage1_7[185]}
   );
   gpc615_5 gpc324 (
      {stage0_7[334], stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338]},
      {stage0_8[55]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[30],stage1_9[64],stage1_8[142],stage1_7[186]}
   );
   gpc615_5 gpc325 (
      {stage0_7[339], stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343]},
      {stage0_8[56]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[31],stage1_9[65],stage1_8[143],stage1_7[187]}
   );
   gpc615_5 gpc326 (
      {stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348]},
      {stage0_8[57]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[32],stage1_9[66],stage1_8[144],stage1_7[188]}
   );
   gpc615_5 gpc327 (
      {stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage0_8[58]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[33],stage1_9[67],stage1_8[145],stage1_7[189]}
   );
   gpc615_5 gpc328 (
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358]},
      {stage0_8[59]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[34],stage1_9[68],stage1_8[146],stage1_7[190]}
   );
   gpc615_5 gpc329 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363]},
      {stage0_8[60]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[35],stage1_9[69],stage1_8[147],stage1_7[191]}
   );
   gpc606_5 gpc330 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[31],stage1_10[36],stage1_9[70],stage1_8[148]}
   );
   gpc606_5 gpc331 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[32],stage1_10[37],stage1_9[71],stage1_8[149]}
   );
   gpc606_5 gpc332 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[33],stage1_10[38],stage1_9[72],stage1_8[150]}
   );
   gpc606_5 gpc333 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[34],stage1_10[39],stage1_9[73],stage1_8[151]}
   );
   gpc606_5 gpc334 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[35],stage1_10[40],stage1_9[74],stage1_8[152]}
   );
   gpc606_5 gpc335 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[36],stage1_10[41],stage1_9[75],stage1_8[153]}
   );
   gpc606_5 gpc336 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[37],stage1_10[42],stage1_9[76],stage1_8[154]}
   );
   gpc606_5 gpc337 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[38],stage1_10[43],stage1_9[77],stage1_8[155]}
   );
   gpc606_5 gpc338 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[39],stage1_10[44],stage1_9[78],stage1_8[156]}
   );
   gpc606_5 gpc339 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[40],stage1_10[45],stage1_9[79],stage1_8[157]}
   );
   gpc606_5 gpc340 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[41],stage1_10[46],stage1_9[80],stage1_8[158]}
   );
   gpc606_5 gpc341 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[42],stage1_10[47],stage1_9[81],stage1_8[159]}
   );
   gpc606_5 gpc342 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[43],stage1_10[48],stage1_9[82],stage1_8[160]}
   );
   gpc606_5 gpc343 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[44],stage1_10[49],stage1_9[83],stage1_8[161]}
   );
   gpc606_5 gpc344 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[45],stage1_10[50],stage1_9[84],stage1_8[162]}
   );
   gpc606_5 gpc345 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[46],stage1_10[51],stage1_9[85],stage1_8[163]}
   );
   gpc606_5 gpc346 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[47],stage1_10[52],stage1_9[86],stage1_8[164]}
   );
   gpc606_5 gpc347 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[48],stage1_10[53],stage1_9[87],stage1_8[165]}
   );
   gpc606_5 gpc348 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[49],stage1_10[54],stage1_9[88],stage1_8[166]}
   );
   gpc606_5 gpc349 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[50],stage1_10[55],stage1_9[89],stage1_8[167]}
   );
   gpc606_5 gpc350 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[51],stage1_10[56],stage1_9[90],stage1_8[168]}
   );
   gpc606_5 gpc351 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[52],stage1_10[57],stage1_9[91],stage1_8[169]}
   );
   gpc606_5 gpc352 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[53],stage1_10[58],stage1_9[92],stage1_8[170]}
   );
   gpc606_5 gpc353 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[54],stage1_10[59],stage1_9[93],stage1_8[171]}
   );
   gpc606_5 gpc354 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[55],stage1_10[60],stage1_9[94],stage1_8[172]}
   );
   gpc606_5 gpc355 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[56],stage1_10[61],stage1_9[95],stage1_8[173]}
   );
   gpc606_5 gpc356 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[57],stage1_10[62],stage1_9[96],stage1_8[174]}
   );
   gpc606_5 gpc357 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[58],stage1_10[63],stage1_9[97],stage1_8[175]}
   );
   gpc606_5 gpc358 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[59],stage1_10[64],stage1_9[98],stage1_8[176]}
   );
   gpc606_5 gpc359 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[60],stage1_10[65],stage1_9[99],stage1_8[177]}
   );
   gpc606_5 gpc360 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[61],stage1_10[66],stage1_9[100],stage1_8[178]}
   );
   gpc606_5 gpc361 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[62],stage1_10[67],stage1_9[101],stage1_8[179]}
   );
   gpc606_5 gpc362 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[63],stage1_10[68],stage1_9[102],stage1_8[180]}
   );
   gpc606_5 gpc363 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[64],stage1_10[69],stage1_9[103],stage1_8[181]}
   );
   gpc606_5 gpc364 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[65],stage1_10[70],stage1_9[104],stage1_8[182]}
   );
   gpc606_5 gpc365 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[66],stage1_10[71],stage1_9[105],stage1_8[183]}
   );
   gpc606_5 gpc366 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[67],stage1_10[72],stage1_9[106],stage1_8[184]}
   );
   gpc606_5 gpc367 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[68],stage1_10[73],stage1_9[107],stage1_8[185]}
   );
   gpc606_5 gpc368 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[69],stage1_10[74],stage1_9[108],stage1_8[186]}
   );
   gpc606_5 gpc369 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[70],stage1_10[75],stage1_9[109],stage1_8[187]}
   );
   gpc606_5 gpc370 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[71],stage1_10[76],stage1_9[110],stage1_8[188]}
   );
   gpc606_5 gpc371 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[72],stage1_10[77],stage1_9[111],stage1_8[189]}
   );
   gpc606_5 gpc372 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[73],stage1_10[78],stage1_9[112],stage1_8[190]}
   );
   gpc606_5 gpc373 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[74],stage1_10[79],stage1_9[113],stage1_8[191]}
   );
   gpc606_5 gpc374 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[75],stage1_10[80],stage1_9[114],stage1_8[192]}
   );
   gpc606_5 gpc375 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[76],stage1_10[81],stage1_9[115],stage1_8[193]}
   );
   gpc606_5 gpc376 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[77],stage1_10[82],stage1_9[116],stage1_8[194]}
   );
   gpc606_5 gpc377 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[78],stage1_10[83],stage1_9[117],stage1_8[195]}
   );
   gpc606_5 gpc378 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[79],stage1_10[84],stage1_9[118],stage1_8[196]}
   );
   gpc606_5 gpc379 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[80],stage1_10[85],stage1_9[119],stage1_8[197]}
   );
   gpc606_5 gpc380 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[81],stage1_10[86],stage1_9[120],stage1_8[198]}
   );
   gpc606_5 gpc381 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[82],stage1_10[87],stage1_9[121],stage1_8[199]}
   );
   gpc606_5 gpc382 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[83],stage1_10[88],stage1_9[122],stage1_8[200]}
   );
   gpc606_5 gpc383 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[84],stage1_10[89],stage1_9[123],stage1_8[201]}
   );
   gpc606_5 gpc384 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[85],stage1_10[90],stage1_9[124],stage1_8[202]}
   );
   gpc606_5 gpc385 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[86],stage1_10[91],stage1_9[125],stage1_8[203]}
   );
   gpc606_5 gpc386 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[87],stage1_10[92],stage1_9[126],stage1_8[204]}
   );
   gpc606_5 gpc387 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[88],stage1_10[93],stage1_9[127],stage1_8[205]}
   );
   gpc606_5 gpc388 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[89],stage1_10[94],stage1_9[128],stage1_8[206]}
   );
   gpc606_5 gpc389 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[90],stage1_10[95],stage1_9[129],stage1_8[207]}
   );
   gpc606_5 gpc390 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[91],stage1_10[96],stage1_9[130],stage1_8[208]}
   );
   gpc606_5 gpc391 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[92],stage1_10[97],stage1_9[131],stage1_8[209]}
   );
   gpc606_5 gpc392 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[93],stage1_10[98],stage1_9[132],stage1_8[210]}
   );
   gpc606_5 gpc393 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[94],stage1_10[99],stage1_9[133],stage1_8[211]}
   );
   gpc606_5 gpc394 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[95],stage1_10[100],stage1_9[134],stage1_8[212]}
   );
   gpc606_5 gpc395 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[96],stage1_10[101],stage1_9[135],stage1_8[213]}
   );
   gpc606_5 gpc396 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[97],stage1_10[102],stage1_9[136],stage1_8[214]}
   );
   gpc606_5 gpc397 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[98],stage1_10[103],stage1_9[137],stage1_8[215]}
   );
   gpc606_5 gpc398 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[99],stage1_10[104],stage1_9[138],stage1_8[216]}
   );
   gpc606_5 gpc399 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[100],stage1_10[105],stage1_9[139],stage1_8[217]}
   );
   gpc606_5 gpc400 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[101],stage1_10[106],stage1_9[140],stage1_8[218]}
   );
   gpc606_5 gpc401 (
      {stage0_8[487], stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[102],stage1_10[107],stage1_9[141],stage1_8[219]}
   );
   gpc606_5 gpc402 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[72],stage1_11[103],stage1_10[108],stage1_9[142]}
   );
   gpc606_5 gpc403 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[73],stage1_11[104],stage1_10[109],stage1_9[143]}
   );
   gpc606_5 gpc404 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[74],stage1_11[105],stage1_10[110],stage1_9[144]}
   );
   gpc606_5 gpc405 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[75],stage1_11[106],stage1_10[111],stage1_9[145]}
   );
   gpc606_5 gpc406 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[76],stage1_11[107],stage1_10[112],stage1_9[146]}
   );
   gpc606_5 gpc407 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[77],stage1_11[108],stage1_10[113],stage1_9[147]}
   );
   gpc606_5 gpc408 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[78],stage1_11[109],stage1_10[114],stage1_9[148]}
   );
   gpc606_5 gpc409 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[79],stage1_11[110],stage1_10[115],stage1_9[149]}
   );
   gpc606_5 gpc410 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[80],stage1_11[111],stage1_10[116],stage1_9[150]}
   );
   gpc606_5 gpc411 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[81],stage1_11[112],stage1_10[117],stage1_9[151]}
   );
   gpc606_5 gpc412 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[82],stage1_11[113],stage1_10[118],stage1_9[152]}
   );
   gpc606_5 gpc413 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[83],stage1_11[114],stage1_10[119],stage1_9[153]}
   );
   gpc606_5 gpc414 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[84],stage1_11[115],stage1_10[120],stage1_9[154]}
   );
   gpc606_5 gpc415 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[85],stage1_11[116],stage1_10[121],stage1_9[155]}
   );
   gpc606_5 gpc416 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[86],stage1_11[117],stage1_10[122],stage1_9[156]}
   );
   gpc606_5 gpc417 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[87],stage1_11[118],stage1_10[123],stage1_9[157]}
   );
   gpc606_5 gpc418 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[88],stage1_11[119],stage1_10[124],stage1_9[158]}
   );
   gpc606_5 gpc419 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[89],stage1_11[120],stage1_10[125],stage1_9[159]}
   );
   gpc606_5 gpc420 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[90],stage1_11[121],stage1_10[126],stage1_9[160]}
   );
   gpc606_5 gpc421 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[91],stage1_11[122],stage1_10[127],stage1_9[161]}
   );
   gpc606_5 gpc422 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[92],stage1_11[123],stage1_10[128],stage1_9[162]}
   );
   gpc615_5 gpc423 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[126]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[21],stage1_12[93],stage1_11[124],stage1_10[129]}
   );
   gpc615_5 gpc424 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[127]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[22],stage1_12[94],stage1_11[125],stage1_10[130]}
   );
   gpc615_5 gpc425 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[128]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[23],stage1_12[95],stage1_11[126],stage1_10[131]}
   );
   gpc615_5 gpc426 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[129]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[24],stage1_12[96],stage1_11[127],stage1_10[132]}
   );
   gpc615_5 gpc427 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[130]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[25],stage1_12[97],stage1_11[128],stage1_10[133]}
   );
   gpc615_5 gpc428 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[131]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[26],stage1_12[98],stage1_11[129],stage1_10[134]}
   );
   gpc615_5 gpc429 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[132]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[27],stage1_12[99],stage1_11[130],stage1_10[135]}
   );
   gpc615_5 gpc430 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[133]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[28],stage1_12[100],stage1_11[131],stage1_10[136]}
   );
   gpc615_5 gpc431 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[134]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[29],stage1_12[101],stage1_11[132],stage1_10[137]}
   );
   gpc615_5 gpc432 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[135]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[30],stage1_12[102],stage1_11[133],stage1_10[138]}
   );
   gpc615_5 gpc433 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[136]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[31],stage1_12[103],stage1_11[134],stage1_10[139]}
   );
   gpc615_5 gpc434 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[137]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[32],stage1_12[104],stage1_11[135],stage1_10[140]}
   );
   gpc615_5 gpc435 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[138]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[33],stage1_12[105],stage1_11[136],stage1_10[141]}
   );
   gpc615_5 gpc436 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[139]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[34],stage1_12[106],stage1_11[137],stage1_10[142]}
   );
   gpc615_5 gpc437 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[84]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[14],stage1_13[35],stage1_12[107],stage1_11[138]}
   );
   gpc615_5 gpc438 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[85]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[15],stage1_13[36],stage1_12[108],stage1_11[139]}
   );
   gpc615_5 gpc439 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[86]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[16],stage1_13[37],stage1_12[109],stage1_11[140]}
   );
   gpc615_5 gpc440 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[87]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[17],stage1_13[38],stage1_12[110],stage1_11[141]}
   );
   gpc615_5 gpc441 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[88]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[18],stage1_13[39],stage1_12[111],stage1_11[142]}
   );
   gpc615_5 gpc442 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[89]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[19],stage1_13[40],stage1_12[112],stage1_11[143]}
   );
   gpc615_5 gpc443 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[90]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[20],stage1_13[41],stage1_12[113],stage1_11[144]}
   );
   gpc615_5 gpc444 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[91]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[21],stage1_13[42],stage1_12[114],stage1_11[145]}
   );
   gpc615_5 gpc445 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[92]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[22],stage1_13[43],stage1_12[115],stage1_11[146]}
   );
   gpc615_5 gpc446 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[93]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[23],stage1_13[44],stage1_12[116],stage1_11[147]}
   );
   gpc615_5 gpc447 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[94]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[24],stage1_13[45],stage1_12[117],stage1_11[148]}
   );
   gpc615_5 gpc448 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[95]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[25],stage1_13[46],stage1_12[118],stage1_11[149]}
   );
   gpc615_5 gpc449 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[96]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[26],stage1_13[47],stage1_12[119],stage1_11[150]}
   );
   gpc615_5 gpc450 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[97]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[27],stage1_13[48],stage1_12[120],stage1_11[151]}
   );
   gpc615_5 gpc451 (
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214]},
      {stage0_12[98]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[28],stage1_13[49],stage1_12[121],stage1_11[152]}
   );
   gpc615_5 gpc452 (
      {stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage0_12[99]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[29],stage1_13[50],stage1_12[122],stage1_11[153]}
   );
   gpc615_5 gpc453 (
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224]},
      {stage0_12[100]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[30],stage1_13[51],stage1_12[123],stage1_11[154]}
   );
   gpc615_5 gpc454 (
      {stage0_11[225], stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229]},
      {stage0_12[101]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[31],stage1_13[52],stage1_12[124],stage1_11[155]}
   );
   gpc615_5 gpc455 (
      {stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233], stage0_11[234]},
      {stage0_12[102]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[32],stage1_13[53],stage1_12[125],stage1_11[156]}
   );
   gpc615_5 gpc456 (
      {stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage0_12[103]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[33],stage1_13[54],stage1_12[126],stage1_11[157]}
   );
   gpc615_5 gpc457 (
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244]},
      {stage0_12[104]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[34],stage1_13[55],stage1_12[127],stage1_11[158]}
   );
   gpc615_5 gpc458 (
      {stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage0_12[105]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[35],stage1_13[56],stage1_12[128],stage1_11[159]}
   );
   gpc615_5 gpc459 (
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254]},
      {stage0_12[106]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[36],stage1_13[57],stage1_12[129],stage1_11[160]}
   );
   gpc615_5 gpc460 (
      {stage0_11[255], stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259]},
      {stage0_12[107]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[37],stage1_13[58],stage1_12[130],stage1_11[161]}
   );
   gpc615_5 gpc461 (
      {stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263], stage0_11[264]},
      {stage0_12[108]},
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage1_15[24],stage1_14[38],stage1_13[59],stage1_12[131],stage1_11[162]}
   );
   gpc615_5 gpc462 (
      {stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage0_12[109]},
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage1_15[25],stage1_14[39],stage1_13[60],stage1_12[132],stage1_11[163]}
   );
   gpc615_5 gpc463 (
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274]},
      {stage0_12[110]},
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage1_15[26],stage1_14[40],stage1_13[61],stage1_12[133],stage1_11[164]}
   );
   gpc615_5 gpc464 (
      {stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage0_12[111]},
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage1_15[27],stage1_14[41],stage1_13[62],stage1_12[134],stage1_11[165]}
   );
   gpc615_5 gpc465 (
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[112]},
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage1_15[28],stage1_14[42],stage1_13[63],stage1_12[135],stage1_11[166]}
   );
   gpc615_5 gpc466 (
      {stage0_11[285], stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289]},
      {stage0_12[113]},
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage1_15[29],stage1_14[43],stage1_13[64],stage1_12[136],stage1_11[167]}
   );
   gpc615_5 gpc467 (
      {stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293], stage0_11[294]},
      {stage0_12[114]},
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage1_15[30],stage1_14[44],stage1_13[65],stage1_12[137],stage1_11[168]}
   );
   gpc615_5 gpc468 (
      {stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage0_12[115]},
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage1_15[31],stage1_14[45],stage1_13[66],stage1_12[138],stage1_11[169]}
   );
   gpc615_5 gpc469 (
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304]},
      {stage0_12[116]},
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage1_15[32],stage1_14[46],stage1_13[67],stage1_12[139],stage1_11[170]}
   );
   gpc615_5 gpc470 (
      {stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage0_12[117]},
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage1_15[33],stage1_14[47],stage1_13[68],stage1_12[140],stage1_11[171]}
   );
   gpc615_5 gpc471 (
      {stage0_11[310], stage0_11[311], stage0_11[312], stage0_11[313], stage0_11[314]},
      {stage0_12[118]},
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage1_15[34],stage1_14[48],stage1_13[69],stage1_12[141],stage1_11[172]}
   );
   gpc615_5 gpc472 (
      {stage0_11[315], stage0_11[316], stage0_11[317], stage0_11[318], stage0_11[319]},
      {stage0_12[119]},
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage1_15[35],stage1_14[49],stage1_13[70],stage1_12[142],stage1_11[173]}
   );
   gpc615_5 gpc473 (
      {stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323], stage0_11[324]},
      {stage0_12[120]},
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage1_15[36],stage1_14[50],stage1_13[71],stage1_12[143],stage1_11[174]}
   );
   gpc615_5 gpc474 (
      {stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage0_12[121]},
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage1_15[37],stage1_14[51],stage1_13[72],stage1_12[144],stage1_11[175]}
   );
   gpc615_5 gpc475 (
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334]},
      {stage0_12[122]},
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage1_15[38],stage1_14[52],stage1_13[73],stage1_12[145],stage1_11[176]}
   );
   gpc615_5 gpc476 (
      {stage0_11[335], stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339]},
      {stage0_12[123]},
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage1_15[39],stage1_14[53],stage1_13[74],stage1_12[146],stage1_11[177]}
   );
   gpc615_5 gpc477 (
      {stage0_11[340], stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344]},
      {stage0_12[124]},
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage1_15[40],stage1_14[54],stage1_13[75],stage1_12[147],stage1_11[178]}
   );
   gpc615_5 gpc478 (
      {stage0_11[345], stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349]},
      {stage0_12[125]},
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage1_15[41],stage1_14[55],stage1_13[76],stage1_12[148],stage1_11[179]}
   );
   gpc615_5 gpc479 (
      {stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354]},
      {stage0_12[126]},
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage1_15[42],stage1_14[56],stage1_13[77],stage1_12[149],stage1_11[180]}
   );
   gpc615_5 gpc480 (
      {stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage0_12[127]},
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage1_15[43],stage1_14[57],stage1_13[78],stage1_12[150],stage1_11[181]}
   );
   gpc615_5 gpc481 (
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364]},
      {stage0_12[128]},
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage1_15[44],stage1_14[58],stage1_13[79],stage1_12[151],stage1_11[182]}
   );
   gpc615_5 gpc482 (
      {stage0_11[365], stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369]},
      {stage0_12[129]},
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage1_15[45],stage1_14[59],stage1_13[80],stage1_12[152],stage1_11[183]}
   );
   gpc615_5 gpc483 (
      {stage0_11[370], stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374]},
      {stage0_12[130]},
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage1_15[46],stage1_14[60],stage1_13[81],stage1_12[153],stage1_11[184]}
   );
   gpc615_5 gpc484 (
      {stage0_11[375], stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379]},
      {stage0_12[131]},
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage1_15[47],stage1_14[61],stage1_13[82],stage1_12[154],stage1_11[185]}
   );
   gpc606_5 gpc485 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[48],stage1_14[62],stage1_13[83],stage1_12[155]}
   );
   gpc606_5 gpc486 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[49],stage1_14[63],stage1_13[84],stage1_12[156]}
   );
   gpc606_5 gpc487 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[50],stage1_14[64],stage1_13[85],stage1_12[157]}
   );
   gpc606_5 gpc488 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[51],stage1_14[65],stage1_13[86],stage1_12[158]}
   );
   gpc606_5 gpc489 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[52],stage1_14[66],stage1_13[87],stage1_12[159]}
   );
   gpc606_5 gpc490 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[53],stage1_14[67],stage1_13[88],stage1_12[160]}
   );
   gpc606_5 gpc491 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[54],stage1_14[68],stage1_13[89],stage1_12[161]}
   );
   gpc606_5 gpc492 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[55],stage1_14[69],stage1_13[90],stage1_12[162]}
   );
   gpc606_5 gpc493 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[56],stage1_14[70],stage1_13[91],stage1_12[163]}
   );
   gpc606_5 gpc494 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[57],stage1_14[71],stage1_13[92],stage1_12[164]}
   );
   gpc606_5 gpc495 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[58],stage1_14[72],stage1_13[93],stage1_12[165]}
   );
   gpc606_5 gpc496 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[59],stage1_14[73],stage1_13[94],stage1_12[166]}
   );
   gpc606_5 gpc497 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[60],stage1_14[74],stage1_13[95],stage1_12[167]}
   );
   gpc606_5 gpc498 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[61],stage1_14[75],stage1_13[96],stage1_12[168]}
   );
   gpc606_5 gpc499 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[62],stage1_14[76],stage1_13[97],stage1_12[169]}
   );
   gpc606_5 gpc500 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[63],stage1_14[77],stage1_13[98],stage1_12[170]}
   );
   gpc606_5 gpc501 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[64],stage1_14[78],stage1_13[99],stage1_12[171]}
   );
   gpc606_5 gpc502 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[65],stage1_14[79],stage1_13[100],stage1_12[172]}
   );
   gpc606_5 gpc503 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[66],stage1_14[80],stage1_13[101],stage1_12[173]}
   );
   gpc606_5 gpc504 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[67],stage1_14[81],stage1_13[102],stage1_12[174]}
   );
   gpc606_5 gpc505 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[68],stage1_14[82],stage1_13[103],stage1_12[175]}
   );
   gpc606_5 gpc506 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[69],stage1_14[83],stage1_13[104],stage1_12[176]}
   );
   gpc606_5 gpc507 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[70],stage1_14[84],stage1_13[105],stage1_12[177]}
   );
   gpc606_5 gpc508 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[71],stage1_14[85],stage1_13[106],stage1_12[178]}
   );
   gpc606_5 gpc509 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[72],stage1_14[86],stage1_13[107],stage1_12[179]}
   );
   gpc606_5 gpc510 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[73],stage1_14[87],stage1_13[108],stage1_12[180]}
   );
   gpc606_5 gpc511 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[74],stage1_14[88],stage1_13[109],stage1_12[181]}
   );
   gpc606_5 gpc512 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[75],stage1_14[89],stage1_13[110],stage1_12[182]}
   );
   gpc606_5 gpc513 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[76],stage1_14[90],stage1_13[111],stage1_12[183]}
   );
   gpc606_5 gpc514 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[77],stage1_14[91],stage1_13[112],stage1_12[184]}
   );
   gpc606_5 gpc515 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[78],stage1_14[92],stage1_13[113],stage1_12[185]}
   );
   gpc606_5 gpc516 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[79],stage1_14[93],stage1_13[114],stage1_12[186]}
   );
   gpc606_5 gpc517 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[80],stage1_14[94],stage1_13[115],stage1_12[187]}
   );
   gpc606_5 gpc518 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[81],stage1_14[95],stage1_13[116],stage1_12[188]}
   );
   gpc606_5 gpc519 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[82],stage1_14[96],stage1_13[117],stage1_12[189]}
   );
   gpc606_5 gpc520 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[83],stage1_14[97],stage1_13[118],stage1_12[190]}
   );
   gpc606_5 gpc521 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[84],stage1_14[98],stage1_13[119],stage1_12[191]}
   );
   gpc606_5 gpc522 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[85],stage1_14[99],stage1_13[120],stage1_12[192]}
   );
   gpc606_5 gpc523 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[86],stage1_14[100],stage1_13[121],stage1_12[193]}
   );
   gpc606_5 gpc524 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[87],stage1_14[101],stage1_13[122],stage1_12[194]}
   );
   gpc606_5 gpc525 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[88],stage1_14[102],stage1_13[123],stage1_12[195]}
   );
   gpc606_5 gpc526 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[89],stage1_14[103],stage1_13[124],stage1_12[196]}
   );
   gpc606_5 gpc527 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[90],stage1_14[104],stage1_13[125],stage1_12[197]}
   );
   gpc606_5 gpc528 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[91],stage1_14[105],stage1_13[126],stage1_12[198]}
   );
   gpc606_5 gpc529 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[92],stage1_14[106],stage1_13[127],stage1_12[199]}
   );
   gpc606_5 gpc530 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[93],stage1_14[107],stage1_13[128],stage1_12[200]}
   );
   gpc606_5 gpc531 (
      {stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[94],stage1_14[108],stage1_13[129],stage1_12[201]}
   );
   gpc606_5 gpc532 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[95],stage1_14[109],stage1_13[130],stage1_12[202]}
   );
   gpc606_5 gpc533 (
      {stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[96],stage1_14[110],stage1_13[131],stage1_12[203]}
   );
   gpc606_5 gpc534 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[97],stage1_14[111],stage1_13[132],stage1_12[204]}
   );
   gpc606_5 gpc535 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[98],stage1_14[112],stage1_13[133],stage1_12[205]}
   );
   gpc606_5 gpc536 (
      {stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[99],stage1_14[113],stage1_13[134],stage1_12[206]}
   );
   gpc606_5 gpc537 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[100],stage1_14[114],stage1_13[135],stage1_12[207]}
   );
   gpc606_5 gpc538 (
      {stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[101],stage1_14[115],stage1_13[136],stage1_12[208]}
   );
   gpc606_5 gpc539 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[102],stage1_14[116],stage1_13[137],stage1_12[209]}
   );
   gpc606_5 gpc540 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[103],stage1_14[117],stage1_13[138],stage1_12[210]}
   );
   gpc606_5 gpc541 (
      {stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[104],stage1_14[118],stage1_13[139],stage1_12[211]}
   );
   gpc606_5 gpc542 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[105],stage1_14[119],stage1_13[140],stage1_12[212]}
   );
   gpc606_5 gpc543 (
      {stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[106],stage1_14[120],stage1_13[141],stage1_12[213]}
   );
   gpc606_5 gpc544 (
      {stage0_12[486], stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[107],stage1_14[121],stage1_13[142],stage1_12[214]}
   );
   gpc606_5 gpc545 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496], stage0_12[497]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[108],stage1_14[122],stage1_13[143],stage1_12[215]}
   );
   gpc606_5 gpc546 (
      {stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501], stage0_12[502], stage0_12[503]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[109],stage1_14[123],stage1_13[144],stage1_12[216]}
   );
   gpc606_5 gpc547 (
      {stage0_12[504], stage0_12[505], stage0_12[506], stage0_12[507], stage0_12[508], stage0_12[509]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[110],stage1_14[124],stage1_13[145],stage1_12[217]}
   );
   gpc606_5 gpc548 (
      {stage0_12[510], stage0_12[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage1_16[63],stage1_15[111],stage1_14[125],stage1_13[146],stage1_12[218]}
   );
   gpc606_5 gpc549 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[64],stage1_15[112],stage1_14[126],stage1_13[147]}
   );
   gpc606_5 gpc550 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[65],stage1_15[113],stage1_14[127],stage1_13[148]}
   );
   gpc606_5 gpc551 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[66],stage1_15[114],stage1_14[128],stage1_13[149]}
   );
   gpc606_5 gpc552 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[67],stage1_15[115],stage1_14[129],stage1_13[150]}
   );
   gpc606_5 gpc553 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[68],stage1_15[116],stage1_14[130],stage1_13[151]}
   );
   gpc606_5 gpc554 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[69],stage1_15[117],stage1_14[131],stage1_13[152]}
   );
   gpc606_5 gpc555 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[70],stage1_15[118],stage1_14[132],stage1_13[153]}
   );
   gpc606_5 gpc556 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[71],stage1_15[119],stage1_14[133],stage1_13[154]}
   );
   gpc606_5 gpc557 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[72],stage1_15[120],stage1_14[134],stage1_13[155]}
   );
   gpc606_5 gpc558 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[73],stage1_15[121],stage1_14[135],stage1_13[156]}
   );
   gpc606_5 gpc559 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[74],stage1_15[122],stage1_14[136],stage1_13[157]}
   );
   gpc606_5 gpc560 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[75],stage1_15[123],stage1_14[137],stage1_13[158]}
   );
   gpc606_5 gpc561 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[76],stage1_15[124],stage1_14[138],stage1_13[159]}
   );
   gpc606_5 gpc562 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[77],stage1_15[125],stage1_14[139],stage1_13[160]}
   );
   gpc606_5 gpc563 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[78],stage1_15[126],stage1_14[140],stage1_13[161]}
   );
   gpc606_5 gpc564 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[79],stage1_15[127],stage1_14[141],stage1_13[162]}
   );
   gpc606_5 gpc565 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[80],stage1_15[128],stage1_14[142],stage1_13[163]}
   );
   gpc606_5 gpc566 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[81],stage1_15[129],stage1_14[143],stage1_13[164]}
   );
   gpc606_5 gpc567 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[82],stage1_15[130],stage1_14[144],stage1_13[165]}
   );
   gpc606_5 gpc568 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[83],stage1_15[131],stage1_14[145],stage1_13[166]}
   );
   gpc606_5 gpc569 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[84],stage1_15[132],stage1_14[146],stage1_13[167]}
   );
   gpc606_5 gpc570 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[85],stage1_15[133],stage1_14[147],stage1_13[168]}
   );
   gpc606_5 gpc571 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[86],stage1_15[134],stage1_14[148],stage1_13[169]}
   );
   gpc606_5 gpc572 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[87],stage1_15[135],stage1_14[149],stage1_13[170]}
   );
   gpc606_5 gpc573 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[88],stage1_15[136],stage1_14[150],stage1_13[171]}
   );
   gpc606_5 gpc574 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[89],stage1_15[137],stage1_14[151],stage1_13[172]}
   );
   gpc606_5 gpc575 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[90],stage1_15[138],stage1_14[152],stage1_13[173]}
   );
   gpc606_5 gpc576 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[91],stage1_15[139],stage1_14[153],stage1_13[174]}
   );
   gpc606_5 gpc577 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[92],stage1_15[140],stage1_14[154],stage1_13[175]}
   );
   gpc606_5 gpc578 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466], stage0_13[467]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[93],stage1_15[141],stage1_14[155],stage1_13[176]}
   );
   gpc606_5 gpc579 (
      {stage0_13[468], stage0_13[469], stage0_13[470], stage0_13[471], stage0_13[472], stage0_13[473]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[94],stage1_15[142],stage1_14[156],stage1_13[177]}
   );
   gpc606_5 gpc580 (
      {stage0_13[474], stage0_13[475], stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[95],stage1_15[143],stage1_14[157],stage1_13[178]}
   );
   gpc606_5 gpc581 (
      {stage0_13[480], stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[96],stage1_15[144],stage1_14[158],stage1_13[179]}
   );
   gpc606_5 gpc582 (
      {stage0_13[486], stage0_13[487], stage0_13[488], stage0_13[489], stage0_13[490], stage0_13[491]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[97],stage1_15[145],stage1_14[159],stage1_13[180]}
   );
   gpc606_5 gpc583 (
      {stage0_13[492], stage0_13[493], stage0_13[494], stage0_13[495], stage0_13[496], stage0_13[497]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[98],stage1_15[146],stage1_14[160],stage1_13[181]}
   );
   gpc606_5 gpc584 (
      {stage0_13[498], stage0_13[499], stage0_13[500], stage0_13[501], stage0_13[502], stage0_13[503]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[99],stage1_15[147],stage1_14[161],stage1_13[182]}
   );
   gpc606_5 gpc585 (
      {stage0_13[504], stage0_13[505], stage0_13[506], stage0_13[507], stage0_13[508], stage0_13[509]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[100],stage1_15[148],stage1_14[162],stage1_13[183]}
   );
   gpc606_5 gpc586 (
      {stage0_13[510], stage0_13[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[101],stage1_15[149],stage1_14[163],stage1_13[184]}
   );
   gpc615_5 gpc587 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388]},
      {stage0_15[228]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[38],stage1_16[102],stage1_15[150],stage1_14[164]}
   );
   gpc615_5 gpc588 (
      {stage0_14[389], stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393]},
      {stage0_15[229]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[39],stage1_16[103],stage1_15[151],stage1_14[165]}
   );
   gpc615_5 gpc589 (
      {stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397], stage0_14[398]},
      {stage0_15[230]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[40],stage1_16[104],stage1_15[152],stage1_14[166]}
   );
   gpc615_5 gpc590 (
      {stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage0_15[231]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[41],stage1_16[105],stage1_15[153],stage1_14[167]}
   );
   gpc615_5 gpc591 (
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408]},
      {stage0_15[232]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[42],stage1_16[106],stage1_15[154],stage1_14[168]}
   );
   gpc615_5 gpc592 (
      {stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_15[233]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[43],stage1_16[107],stage1_15[155],stage1_14[169]}
   );
   gpc615_5 gpc593 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_15[234]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[44],stage1_16[108],stage1_15[156],stage1_14[170]}
   );
   gpc615_5 gpc594 (
      {stage0_14[419], stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423]},
      {stage0_15[235]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[45],stage1_16[109],stage1_15[157],stage1_14[171]}
   );
   gpc615_5 gpc595 (
      {stage0_14[424], stage0_14[425], stage0_14[426], stage0_14[427], stage0_14[428]},
      {stage0_15[236]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[46],stage1_16[110],stage1_15[158],stage1_14[172]}
   );
   gpc615_5 gpc596 (
      {stage0_15[237], stage0_15[238], stage0_15[239], stage0_15[240], stage0_15[241]},
      {stage0_16[54]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[9],stage1_17[47],stage1_16[111],stage1_15[159]}
   );
   gpc615_5 gpc597 (
      {stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245], stage0_15[246]},
      {stage0_16[55]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[10],stage1_17[48],stage1_16[112],stage1_15[160]}
   );
   gpc615_5 gpc598 (
      {stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage0_16[56]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[11],stage1_17[49],stage1_16[113],stage1_15[161]}
   );
   gpc615_5 gpc599 (
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256]},
      {stage0_16[57]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[12],stage1_17[50],stage1_16[114],stage1_15[162]}
   );
   gpc615_5 gpc600 (
      {stage0_15[257], stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261]},
      {stage0_16[58]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[13],stage1_17[51],stage1_16[115],stage1_15[163]}
   );
   gpc615_5 gpc601 (
      {stage0_15[262], stage0_15[263], stage0_15[264], stage0_15[265], stage0_15[266]},
      {stage0_16[59]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[14],stage1_17[52],stage1_16[116],stage1_15[164]}
   );
   gpc615_5 gpc602 (
      {stage0_15[267], stage0_15[268], stage0_15[269], stage0_15[270], stage0_15[271]},
      {stage0_16[60]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[15],stage1_17[53],stage1_16[117],stage1_15[165]}
   );
   gpc615_5 gpc603 (
      {stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275], stage0_15[276]},
      {stage0_16[61]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[16],stage1_17[54],stage1_16[118],stage1_15[166]}
   );
   gpc615_5 gpc604 (
      {stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage0_16[62]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[17],stage1_17[55],stage1_16[119],stage1_15[167]}
   );
   gpc615_5 gpc605 (
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286]},
      {stage0_16[63]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[18],stage1_17[56],stage1_16[120],stage1_15[168]}
   );
   gpc615_5 gpc606 (
      {stage0_15[287], stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291]},
      {stage0_16[64]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[19],stage1_17[57],stage1_16[121],stage1_15[169]}
   );
   gpc615_5 gpc607 (
      {stage0_15[292], stage0_15[293], stage0_15[294], stage0_15[295], stage0_15[296]},
      {stage0_16[65]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[20],stage1_17[58],stage1_16[122],stage1_15[170]}
   );
   gpc615_5 gpc608 (
      {stage0_15[297], stage0_15[298], stage0_15[299], stage0_15[300], stage0_15[301]},
      {stage0_16[66]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[21],stage1_17[59],stage1_16[123],stage1_15[171]}
   );
   gpc615_5 gpc609 (
      {stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305], stage0_15[306]},
      {stage0_16[67]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[22],stage1_17[60],stage1_16[124],stage1_15[172]}
   );
   gpc615_5 gpc610 (
      {stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage0_16[68]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[23],stage1_17[61],stage1_16[125],stage1_15[173]}
   );
   gpc615_5 gpc611 (
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316]},
      {stage0_16[69]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[24],stage1_17[62],stage1_16[126],stage1_15[174]}
   );
   gpc615_5 gpc612 (
      {stage0_15[317], stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321]},
      {stage0_16[70]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[25],stage1_17[63],stage1_16[127],stage1_15[175]}
   );
   gpc615_5 gpc613 (
      {stage0_15[322], stage0_15[323], stage0_15[324], stage0_15[325], stage0_15[326]},
      {stage0_16[71]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[26],stage1_17[64],stage1_16[128],stage1_15[176]}
   );
   gpc615_5 gpc614 (
      {stage0_15[327], stage0_15[328], stage0_15[329], stage0_15[330], stage0_15[331]},
      {stage0_16[72]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[27],stage1_17[65],stage1_16[129],stage1_15[177]}
   );
   gpc615_5 gpc615 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336]},
      {stage0_16[73]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[28],stage1_17[66],stage1_16[130],stage1_15[178]}
   );
   gpc615_5 gpc616 (
      {stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage0_16[74]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[29],stage1_17[67],stage1_16[131],stage1_15[179]}
   );
   gpc615_5 gpc617 (
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346]},
      {stage0_16[75]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[30],stage1_17[68],stage1_16[132],stage1_15[180]}
   );
   gpc615_5 gpc618 (
      {stage0_15[347], stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351]},
      {stage0_16[76]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[31],stage1_17[69],stage1_16[133],stage1_15[181]}
   );
   gpc615_5 gpc619 (
      {stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355], stage0_15[356]},
      {stage0_16[77]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[32],stage1_17[70],stage1_16[134],stage1_15[182]}
   );
   gpc615_5 gpc620 (
      {stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360], stage0_15[361]},
      {stage0_16[78]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[33],stage1_17[71],stage1_16[135],stage1_15[183]}
   );
   gpc615_5 gpc621 (
      {stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365], stage0_15[366]},
      {stage0_16[79]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[34],stage1_17[72],stage1_16[136],stage1_15[184]}
   );
   gpc615_5 gpc622 (
      {stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage0_16[80]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[35],stage1_17[73],stage1_16[137],stage1_15[185]}
   );
   gpc615_5 gpc623 (
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376]},
      {stage0_16[81]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[36],stage1_17[74],stage1_16[138],stage1_15[186]}
   );
   gpc615_5 gpc624 (
      {stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381]},
      {stage0_16[82]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[37],stage1_17[75],stage1_16[139],stage1_15[187]}
   );
   gpc615_5 gpc625 (
      {stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385], stage0_15[386]},
      {stage0_16[83]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[38],stage1_17[76],stage1_16[140],stage1_15[188]}
   );
   gpc615_5 gpc626 (
      {stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390], stage0_15[391]},
      {stage0_16[84]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[39],stage1_17[77],stage1_16[141],stage1_15[189]}
   );
   gpc615_5 gpc627 (
      {stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395], stage0_15[396]},
      {stage0_16[85]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[40],stage1_17[78],stage1_16[142],stage1_15[190]}
   );
   gpc615_5 gpc628 (
      {stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage0_16[86]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[41],stage1_17[79],stage1_16[143],stage1_15[191]}
   );
   gpc615_5 gpc629 (
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406]},
      {stage0_16[87]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[42],stage1_17[80],stage1_16[144],stage1_15[192]}
   );
   gpc615_5 gpc630 (
      {stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411]},
      {stage0_16[88]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[43],stage1_17[81],stage1_16[145],stage1_15[193]}
   );
   gpc615_5 gpc631 (
      {stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415], stage0_15[416]},
      {stage0_16[89]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[44],stage1_17[82],stage1_16[146],stage1_15[194]}
   );
   gpc615_5 gpc632 (
      {stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420], stage0_15[421]},
      {stage0_16[90]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[45],stage1_17[83],stage1_16[147],stage1_15[195]}
   );
   gpc615_5 gpc633 (
      {stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425], stage0_15[426]},
      {stage0_16[91]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[46],stage1_17[84],stage1_16[148],stage1_15[196]}
   );
   gpc615_5 gpc634 (
      {stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage0_16[92]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[47],stage1_17[85],stage1_16[149],stage1_15[197]}
   );
   gpc615_5 gpc635 (
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436]},
      {stage0_16[93]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[48],stage1_17[86],stage1_16[150],stage1_15[198]}
   );
   gpc615_5 gpc636 (
      {stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441]},
      {stage0_16[94]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[49],stage1_17[87],stage1_16[151],stage1_15[199]}
   );
   gpc615_5 gpc637 (
      {stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445], stage0_15[446]},
      {stage0_16[95]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[50],stage1_17[88],stage1_16[152],stage1_15[200]}
   );
   gpc615_5 gpc638 (
      {stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450], stage0_15[451]},
      {stage0_16[96]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[51],stage1_17[89],stage1_16[153],stage1_15[201]}
   );
   gpc615_5 gpc639 (
      {stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455], stage0_15[456]},
      {stage0_16[97]},
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage1_19[43],stage1_18[52],stage1_17[90],stage1_16[154],stage1_15[202]}
   );
   gpc606_5 gpc640 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[44],stage1_18[53],stage1_17[91],stage1_16[155]}
   );
   gpc606_5 gpc641 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[45],stage1_18[54],stage1_17[92],stage1_16[156]}
   );
   gpc606_5 gpc642 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[46],stage1_18[55],stage1_17[93],stage1_16[157]}
   );
   gpc606_5 gpc643 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[47],stage1_18[56],stage1_17[94],stage1_16[158]}
   );
   gpc606_5 gpc644 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[48],stage1_18[57],stage1_17[95],stage1_16[159]}
   );
   gpc606_5 gpc645 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[49],stage1_18[58],stage1_17[96],stage1_16[160]}
   );
   gpc606_5 gpc646 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[50],stage1_18[59],stage1_17[97],stage1_16[161]}
   );
   gpc606_5 gpc647 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[51],stage1_18[60],stage1_17[98],stage1_16[162]}
   );
   gpc606_5 gpc648 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[52],stage1_18[61],stage1_17[99],stage1_16[163]}
   );
   gpc606_5 gpc649 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[53],stage1_18[62],stage1_17[100],stage1_16[164]}
   );
   gpc606_5 gpc650 (
      {stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[54],stage1_18[63],stage1_17[101],stage1_16[165]}
   );
   gpc606_5 gpc651 (
      {stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[55],stage1_18[64],stage1_17[102],stage1_16[166]}
   );
   gpc606_5 gpc652 (
      {stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[56],stage1_18[65],stage1_17[103],stage1_16[167]}
   );
   gpc606_5 gpc653 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[57],stage1_18[66],stage1_17[104],stage1_16[168]}
   );
   gpc606_5 gpc654 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[58],stage1_18[67],stage1_17[105],stage1_16[169]}
   );
   gpc606_5 gpc655 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[59],stage1_18[68],stage1_17[106],stage1_16[170]}
   );
   gpc606_5 gpc656 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[60],stage1_18[69],stage1_17[107],stage1_16[171]}
   );
   gpc606_5 gpc657 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[61],stage1_18[70],stage1_17[108],stage1_16[172]}
   );
   gpc606_5 gpc658 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[62],stage1_18[71],stage1_17[109],stage1_16[173]}
   );
   gpc606_5 gpc659 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[63],stage1_18[72],stage1_17[110],stage1_16[174]}
   );
   gpc606_5 gpc660 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[64],stage1_18[73],stage1_17[111],stage1_16[175]}
   );
   gpc606_5 gpc661 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[65],stage1_18[74],stage1_17[112],stage1_16[176]}
   );
   gpc606_5 gpc662 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[66],stage1_18[75],stage1_17[113],stage1_16[177]}
   );
   gpc606_5 gpc663 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[67],stage1_18[76],stage1_17[114],stage1_16[178]}
   );
   gpc606_5 gpc664 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[68],stage1_18[77],stage1_17[115],stage1_16[179]}
   );
   gpc606_5 gpc665 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[69],stage1_18[78],stage1_17[116],stage1_16[180]}
   );
   gpc606_5 gpc666 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[70],stage1_18[79],stage1_17[117],stage1_16[181]}
   );
   gpc606_5 gpc667 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[71],stage1_18[80],stage1_17[118],stage1_16[182]}
   );
   gpc606_5 gpc668 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[72],stage1_18[81],stage1_17[119],stage1_16[183]}
   );
   gpc606_5 gpc669 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[73],stage1_18[82],stage1_17[120],stage1_16[184]}
   );
   gpc606_5 gpc670 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[74],stage1_18[83],stage1_17[121],stage1_16[185]}
   );
   gpc606_5 gpc671 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[75],stage1_18[84],stage1_17[122],stage1_16[186]}
   );
   gpc606_5 gpc672 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[76],stage1_18[85],stage1_17[123],stage1_16[187]}
   );
   gpc606_5 gpc673 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[77],stage1_18[86],stage1_17[124],stage1_16[188]}
   );
   gpc606_5 gpc674 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[78],stage1_18[87],stage1_17[125],stage1_16[189]}
   );
   gpc606_5 gpc675 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[79],stage1_18[88],stage1_17[126],stage1_16[190]}
   );
   gpc606_5 gpc676 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[80],stage1_18[89],stage1_17[127],stage1_16[191]}
   );
   gpc606_5 gpc677 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[81],stage1_18[90],stage1_17[128],stage1_16[192]}
   );
   gpc606_5 gpc678 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[82],stage1_18[91],stage1_17[129],stage1_16[193]}
   );
   gpc606_5 gpc679 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[83],stage1_18[92],stage1_17[130],stage1_16[194]}
   );
   gpc606_5 gpc680 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[84],stage1_18[93],stage1_17[131],stage1_16[195]}
   );
   gpc606_5 gpc681 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[85],stage1_18[94],stage1_17[132],stage1_16[196]}
   );
   gpc606_5 gpc682 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[86],stage1_18[95],stage1_17[133],stage1_16[197]}
   );
   gpc606_5 gpc683 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[87],stage1_18[96],stage1_17[134],stage1_16[198]}
   );
   gpc606_5 gpc684 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[88],stage1_18[97],stage1_17[135],stage1_16[199]}
   );
   gpc606_5 gpc685 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[89],stage1_18[98],stage1_17[136],stage1_16[200]}
   );
   gpc606_5 gpc686 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[90],stage1_18[99],stage1_17[137],stage1_16[201]}
   );
   gpc606_5 gpc687 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[91],stage1_18[100],stage1_17[138],stage1_16[202]}
   );
   gpc606_5 gpc688 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[92],stage1_18[101],stage1_17[139],stage1_16[203]}
   );
   gpc606_5 gpc689 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[93],stage1_18[102],stage1_17[140],stage1_16[204]}
   );
   gpc606_5 gpc690 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[94],stage1_18[103],stage1_17[141],stage1_16[205]}
   );
   gpc606_5 gpc691 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[95],stage1_18[104],stage1_17[142],stage1_16[206]}
   );
   gpc606_5 gpc692 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[96],stage1_18[105],stage1_17[143],stage1_16[207]}
   );
   gpc606_5 gpc693 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[97],stage1_18[106],stage1_17[144],stage1_16[208]}
   );
   gpc606_5 gpc694 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[98],stage1_18[107],stage1_17[145],stage1_16[209]}
   );
   gpc606_5 gpc695 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[99],stage1_18[108],stage1_17[146],stage1_16[210]}
   );
   gpc606_5 gpc696 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[100],stage1_18[109],stage1_17[147],stage1_16[211]}
   );
   gpc606_5 gpc697 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[101],stage1_18[110],stage1_17[148],stage1_16[212]}
   );
   gpc606_5 gpc698 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[102],stage1_18[111],stage1_17[149],stage1_16[213]}
   );
   gpc606_5 gpc699 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[103],stage1_18[112],stage1_17[150],stage1_16[214]}
   );
   gpc606_5 gpc700 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[104],stage1_18[113],stage1_17[151],stage1_16[215]}
   );
   gpc606_5 gpc701 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[105],stage1_18[114],stage1_17[152],stage1_16[216]}
   );
   gpc606_5 gpc702 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[106],stage1_18[115],stage1_17[153],stage1_16[217]}
   );
   gpc606_5 gpc703 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[107],stage1_18[116],stage1_17[154],stage1_16[218]}
   );
   gpc606_5 gpc704 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[108],stage1_18[117],stage1_17[155],stage1_16[219]}
   );
   gpc606_5 gpc705 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[109],stage1_18[118],stage1_17[156],stage1_16[220]}
   );
   gpc606_5 gpc706 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[110],stage1_18[119],stage1_17[157],stage1_16[221]}
   );
   gpc606_5 gpc707 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[111],stage1_18[120],stage1_17[158],stage1_16[222]}
   );
   gpc606_5 gpc708 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[112],stage1_18[121],stage1_17[159],stage1_16[223]}
   );
   gpc606_5 gpc709 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[69],stage1_19[113],stage1_18[122],stage1_17[160]}
   );
   gpc606_5 gpc710 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[70],stage1_19[114],stage1_18[123],stage1_17[161]}
   );
   gpc606_5 gpc711 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[71],stage1_19[115],stage1_18[124],stage1_17[162]}
   );
   gpc606_5 gpc712 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[72],stage1_19[116],stage1_18[125],stage1_17[163]}
   );
   gpc606_5 gpc713 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[73],stage1_19[117],stage1_18[126],stage1_17[164]}
   );
   gpc606_5 gpc714 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[74],stage1_19[118],stage1_18[127],stage1_17[165]}
   );
   gpc606_5 gpc715 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[75],stage1_19[119],stage1_18[128],stage1_17[166]}
   );
   gpc606_5 gpc716 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[76],stage1_19[120],stage1_18[129],stage1_17[167]}
   );
   gpc606_5 gpc717 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[77],stage1_19[121],stage1_18[130],stage1_17[168]}
   );
   gpc606_5 gpc718 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[78],stage1_19[122],stage1_18[131],stage1_17[169]}
   );
   gpc606_5 gpc719 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[79],stage1_19[123],stage1_18[132],stage1_17[170]}
   );
   gpc606_5 gpc720 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[80],stage1_19[124],stage1_18[133],stage1_17[171]}
   );
   gpc606_5 gpc721 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[81],stage1_19[125],stage1_18[134],stage1_17[172]}
   );
   gpc606_5 gpc722 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[82],stage1_19[126],stage1_18[135],stage1_17[173]}
   );
   gpc606_5 gpc723 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[83],stage1_19[127],stage1_18[136],stage1_17[174]}
   );
   gpc606_5 gpc724 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[84],stage1_19[128],stage1_18[137],stage1_17[175]}
   );
   gpc606_5 gpc725 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[85],stage1_19[129],stage1_18[138],stage1_17[176]}
   );
   gpc606_5 gpc726 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[86],stage1_19[130],stage1_18[139],stage1_17[177]}
   );
   gpc606_5 gpc727 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[87],stage1_19[131],stage1_18[140],stage1_17[178]}
   );
   gpc606_5 gpc728 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[88],stage1_19[132],stage1_18[141],stage1_17[179]}
   );
   gpc606_5 gpc729 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[89],stage1_19[133],stage1_18[142],stage1_17[180]}
   );
   gpc606_5 gpc730 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[90],stage1_19[134],stage1_18[143],stage1_17[181]}
   );
   gpc606_5 gpc731 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[91],stage1_19[135],stage1_18[144],stage1_17[182]}
   );
   gpc606_5 gpc732 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[92],stage1_19[136],stage1_18[145],stage1_17[183]}
   );
   gpc606_5 gpc733 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[93],stage1_19[137],stage1_18[146],stage1_17[184]}
   );
   gpc606_5 gpc734 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[94],stage1_19[138],stage1_18[147],stage1_17[185]}
   );
   gpc606_5 gpc735 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[95],stage1_19[139],stage1_18[148],stage1_17[186]}
   );
   gpc606_5 gpc736 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[96],stage1_19[140],stage1_18[149],stage1_17[187]}
   );
   gpc606_5 gpc737 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[97],stage1_19[141],stage1_18[150],stage1_17[188]}
   );
   gpc606_5 gpc738 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[98],stage1_19[142],stage1_18[151],stage1_17[189]}
   );
   gpc606_5 gpc739 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[99],stage1_19[143],stage1_18[152],stage1_17[190]}
   );
   gpc606_5 gpc740 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[100],stage1_19[144],stage1_18[153],stage1_17[191]}
   );
   gpc606_5 gpc741 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[101],stage1_19[145],stage1_18[154],stage1_17[192]}
   );
   gpc606_5 gpc742 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[102],stage1_19[146],stage1_18[155],stage1_17[193]}
   );
   gpc606_5 gpc743 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[103],stage1_19[147],stage1_18[156],stage1_17[194]}
   );
   gpc606_5 gpc744 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[104],stage1_19[148],stage1_18[157],stage1_17[195]}
   );
   gpc606_5 gpc745 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[105],stage1_19[149],stage1_18[158],stage1_17[196]}
   );
   gpc606_5 gpc746 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[106],stage1_19[150],stage1_18[159],stage1_17[197]}
   );
   gpc615_5 gpc747 (
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418]},
      {stage0_19[228]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[107],stage1_19[151],stage1_18[160]}
   );
   gpc615_5 gpc748 (
      {stage0_18[419], stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423]},
      {stage0_19[229]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[108],stage1_19[152],stage1_18[161]}
   );
   gpc615_5 gpc749 (
      {stage0_18[424], stage0_18[425], stage0_18[426], stage0_18[427], stage0_18[428]},
      {stage0_19[230]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[109],stage1_19[153],stage1_18[162]}
   );
   gpc615_5 gpc750 (
      {stage0_18[429], stage0_18[430], stage0_18[431], stage0_18[432], stage0_18[433]},
      {stage0_19[231]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[110],stage1_19[154],stage1_18[163]}
   );
   gpc615_5 gpc751 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[24]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[42],stage1_20[111],stage1_19[155]}
   );
   gpc615_5 gpc752 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[25]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[43],stage1_20[112],stage1_19[156]}
   );
   gpc615_5 gpc753 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[26]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[44],stage1_20[113],stage1_19[157]}
   );
   gpc615_5 gpc754 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[27]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[7],stage1_21[45],stage1_20[114],stage1_19[158]}
   );
   gpc615_5 gpc755 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[28]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[8],stage1_21[46],stage1_20[115],stage1_19[159]}
   );
   gpc615_5 gpc756 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[29]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[9],stage1_21[47],stage1_20[116],stage1_19[160]}
   );
   gpc615_5 gpc757 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[30]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[10],stage1_21[48],stage1_20[117],stage1_19[161]}
   );
   gpc615_5 gpc758 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[31]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[11],stage1_21[49],stage1_20[118],stage1_19[162]}
   );
   gpc615_5 gpc759 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[32]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[12],stage1_21[50],stage1_20[119],stage1_19[163]}
   );
   gpc615_5 gpc760 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[33]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[13],stage1_21[51],stage1_20[120],stage1_19[164]}
   );
   gpc615_5 gpc761 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[34]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[14],stage1_21[52],stage1_20[121],stage1_19[165]}
   );
   gpc615_5 gpc762 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[35]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[15],stage1_21[53],stage1_20[122],stage1_19[166]}
   );
   gpc615_5 gpc763 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[36]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[16],stage1_21[54],stage1_20[123],stage1_19[167]}
   );
   gpc615_5 gpc764 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[37]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[17],stage1_21[55],stage1_20[124],stage1_19[168]}
   );
   gpc615_5 gpc765 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[38]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[18],stage1_21[56],stage1_20[125],stage1_19[169]}
   );
   gpc615_5 gpc766 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[39]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[19],stage1_21[57],stage1_20[126],stage1_19[170]}
   );
   gpc615_5 gpc767 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[40]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[20],stage1_21[58],stage1_20[127],stage1_19[171]}
   );
   gpc615_5 gpc768 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[41]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[21],stage1_21[59],stage1_20[128],stage1_19[172]}
   );
   gpc615_5 gpc769 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[42]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[22],stage1_21[60],stage1_20[129],stage1_19[173]}
   );
   gpc615_5 gpc770 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[43]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[23],stage1_21[61],stage1_20[130],stage1_19[174]}
   );
   gpc615_5 gpc771 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[44]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[24],stage1_21[62],stage1_20[131],stage1_19[175]}
   );
   gpc615_5 gpc772 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[45]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[25],stage1_21[63],stage1_20[132],stage1_19[176]}
   );
   gpc615_5 gpc773 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[46]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[26],stage1_21[64],stage1_20[133],stage1_19[177]}
   );
   gpc615_5 gpc774 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[47]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[27],stage1_21[65],stage1_20[134],stage1_19[178]}
   );
   gpc615_5 gpc775 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[48]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[28],stage1_21[66],stage1_20[135],stage1_19[179]}
   );
   gpc615_5 gpc776 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[49]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[29],stage1_21[67],stage1_20[136],stage1_19[180]}
   );
   gpc615_5 gpc777 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[50]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[30],stage1_21[68],stage1_20[137],stage1_19[181]}
   );
   gpc615_5 gpc778 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[51]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[31],stage1_21[69],stage1_20[138],stage1_19[182]}
   );
   gpc615_5 gpc779 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[52]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[32],stage1_21[70],stage1_20[139],stage1_19[183]}
   );
   gpc615_5 gpc780 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[53]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[33],stage1_21[71],stage1_20[140],stage1_19[184]}
   );
   gpc615_5 gpc781 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[54]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[34],stage1_21[72],stage1_20[141],stage1_19[185]}
   );
   gpc615_5 gpc782 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[55]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[35],stage1_21[73],stage1_20[142],stage1_19[186]}
   );
   gpc615_5 gpc783 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[56]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[36],stage1_21[74],stage1_20[143],stage1_19[187]}
   );
   gpc615_5 gpc784 (
      {stage0_19[397], stage0_19[398], stage0_19[399], stage0_19[400], stage0_19[401]},
      {stage0_20[57]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[37],stage1_21[75],stage1_20[144],stage1_19[188]}
   );
   gpc615_5 gpc785 (
      {stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405], stage0_19[406]},
      {stage0_20[58]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[38],stage1_21[76],stage1_20[145],stage1_19[189]}
   );
   gpc615_5 gpc786 (
      {stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410], stage0_19[411]},
      {stage0_20[59]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[39],stage1_21[77],stage1_20[146],stage1_19[190]}
   );
   gpc615_5 gpc787 (
      {stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415], stage0_19[416]},
      {stage0_20[60]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[40],stage1_21[78],stage1_20[147],stage1_19[191]}
   );
   gpc615_5 gpc788 (
      {stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420], stage0_19[421]},
      {stage0_20[61]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[41],stage1_21[79],stage1_20[148],stage1_19[192]}
   );
   gpc615_5 gpc789 (
      {stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425], stage0_19[426]},
      {stage0_20[62]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[42],stage1_21[80],stage1_20[149],stage1_19[193]}
   );
   gpc615_5 gpc790 (
      {stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430], stage0_19[431]},
      {stage0_20[63]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[43],stage1_21[81],stage1_20[150],stage1_19[194]}
   );
   gpc615_5 gpc791 (
      {stage0_19[432], stage0_19[433], stage0_19[434], stage0_19[435], stage0_19[436]},
      {stage0_20[64]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[44],stage1_21[82],stage1_20[151],stage1_19[195]}
   );
   gpc615_5 gpc792 (
      {stage0_19[437], stage0_19[438], stage0_19[439], stage0_19[440], stage0_19[441]},
      {stage0_20[65]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage1_23[41],stage1_22[45],stage1_21[83],stage1_20[152],stage1_19[196]}
   );
   gpc615_5 gpc793 (
      {stage0_19[442], stage0_19[443], stage0_19[444], stage0_19[445], stage0_19[446]},
      {stage0_20[66]},
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage1_23[42],stage1_22[46],stage1_21[84],stage1_20[153],stage1_19[197]}
   );
   gpc615_5 gpc794 (
      {stage0_19[447], stage0_19[448], stage0_19[449], stage0_19[450], stage0_19[451]},
      {stage0_20[67]},
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage1_23[43],stage1_22[47],stage1_21[85],stage1_20[154],stage1_19[198]}
   );
   gpc615_5 gpc795 (
      {stage0_19[452], stage0_19[453], stage0_19[454], stage0_19[455], stage0_19[456]},
      {stage0_20[68]},
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage1_23[44],stage1_22[48],stage1_21[86],stage1_20[155],stage1_19[199]}
   );
   gpc615_5 gpc796 (
      {stage0_19[457], stage0_19[458], stage0_19[459], stage0_19[460], stage0_19[461]},
      {stage0_20[69]},
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage1_23[45],stage1_22[49],stage1_21[87],stage1_20[156],stage1_19[200]}
   );
   gpc615_5 gpc797 (
      {stage0_19[462], stage0_19[463], stage0_19[464], stage0_19[465], stage0_19[466]},
      {stage0_20[70]},
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage1_23[46],stage1_22[50],stage1_21[88],stage1_20[157],stage1_19[201]}
   );
   gpc615_5 gpc798 (
      {stage0_19[467], stage0_19[468], stage0_19[469], stage0_19[470], stage0_19[471]},
      {stage0_20[71]},
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage1_23[47],stage1_22[51],stage1_21[89],stage1_20[158],stage1_19[202]}
   );
   gpc615_5 gpc799 (
      {stage0_19[472], stage0_19[473], stage0_19[474], stage0_19[475], stage0_19[476]},
      {stage0_20[72]},
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage1_23[48],stage1_22[52],stage1_21[90],stage1_20[159],stage1_19[203]}
   );
   gpc615_5 gpc800 (
      {stage0_19[477], stage0_19[478], stage0_19[479], stage0_19[480], stage0_19[481]},
      {stage0_20[73]},
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage1_23[49],stage1_22[53],stage1_21[91],stage1_20[160],stage1_19[204]}
   );
   gpc615_5 gpc801 (
      {stage0_19[482], stage0_19[483], stage0_19[484], stage0_19[485], stage0_19[486]},
      {stage0_20[74]},
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage1_23[50],stage1_22[54],stage1_21[92],stage1_20[161],stage1_19[205]}
   );
   gpc615_5 gpc802 (
      {stage0_19[487], stage0_19[488], stage0_19[489], stage0_19[490], stage0_19[491]},
      {stage0_20[75]},
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage1_23[51],stage1_22[55],stage1_21[93],stage1_20[162],stage1_19[206]}
   );
   gpc615_5 gpc803 (
      {stage0_19[492], stage0_19[493], stage0_19[494], stage0_19[495], stage0_19[496]},
      {stage0_20[76]},
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage1_23[52],stage1_22[56],stage1_21[94],stage1_20[163],stage1_19[207]}
   );
   gpc615_5 gpc804 (
      {stage0_19[497], stage0_19[498], stage0_19[499], stage0_19[500], stage0_19[501]},
      {stage0_20[77]},
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage1_23[53],stage1_22[57],stage1_21[95],stage1_20[164],stage1_19[208]}
   );
   gpc606_5 gpc805 (
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[54],stage1_22[58],stage1_21[96],stage1_20[165]}
   );
   gpc606_5 gpc806 (
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[55],stage1_22[59],stage1_21[97],stage1_20[166]}
   );
   gpc606_5 gpc807 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[56],stage1_22[60],stage1_21[98],stage1_20[167]}
   );
   gpc606_5 gpc808 (
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[57],stage1_22[61],stage1_21[99],stage1_20[168]}
   );
   gpc606_5 gpc809 (
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[58],stage1_22[62],stage1_21[100],stage1_20[169]}
   );
   gpc606_5 gpc810 (
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[59],stage1_22[63],stage1_21[101],stage1_20[170]}
   );
   gpc606_5 gpc811 (
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[60],stage1_22[64],stage1_21[102],stage1_20[171]}
   );
   gpc606_5 gpc812 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[61],stage1_22[65],stage1_21[103],stage1_20[172]}
   );
   gpc606_5 gpc813 (
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[62],stage1_22[66],stage1_21[104],stage1_20[173]}
   );
   gpc606_5 gpc814 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[63],stage1_22[67],stage1_21[105],stage1_20[174]}
   );
   gpc606_5 gpc815 (
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[64],stage1_22[68],stage1_21[106],stage1_20[175]}
   );
   gpc606_5 gpc816 (
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[65],stage1_22[69],stage1_21[107],stage1_20[176]}
   );
   gpc606_5 gpc817 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[66],stage1_22[70],stage1_21[108],stage1_20[177]}
   );
   gpc606_5 gpc818 (
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[67],stage1_22[71],stage1_21[109],stage1_20[178]}
   );
   gpc606_5 gpc819 (
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[68],stage1_22[72],stage1_21[110],stage1_20[179]}
   );
   gpc606_5 gpc820 (
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[69],stage1_22[73],stage1_21[111],stage1_20[180]}
   );
   gpc606_5 gpc821 (
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[70],stage1_22[74],stage1_21[112],stage1_20[181]}
   );
   gpc606_5 gpc822 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[71],stage1_22[75],stage1_21[113],stage1_20[182]}
   );
   gpc606_5 gpc823 (
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[72],stage1_22[76],stage1_21[114],stage1_20[183]}
   );
   gpc606_5 gpc824 (
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[73],stage1_22[77],stage1_21[115],stage1_20[184]}
   );
   gpc606_5 gpc825 (
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[74],stage1_22[78],stage1_21[116],stage1_20[185]}
   );
   gpc606_5 gpc826 (
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[75],stage1_22[79],stage1_21[117],stage1_20[186]}
   );
   gpc606_5 gpc827 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[76],stage1_22[80],stage1_21[118],stage1_20[187]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[77],stage1_22[81],stage1_21[119],stage1_20[188]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[78],stage1_22[82],stage1_21[120],stage1_20[189]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[79],stage1_22[83],stage1_21[121],stage1_20[190]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[80],stage1_22[84],stage1_21[122],stage1_20[191]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[81],stage1_22[85],stage1_21[123],stage1_20[192]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[82],stage1_22[86],stage1_21[124],stage1_20[193]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[83],stage1_22[87],stage1_21[125],stage1_20[194]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[84],stage1_22[88],stage1_21[126],stage1_20[195]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[85],stage1_22[89],stage1_21[127],stage1_20[196]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[86],stage1_22[90],stage1_21[128],stage1_20[197]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[87],stage1_22[91],stage1_21[129],stage1_20[198]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[88],stage1_22[92],stage1_21[130],stage1_20[199]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[89],stage1_22[93],stage1_21[131],stage1_20[200]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[90],stage1_22[94],stage1_21[132],stage1_20[201]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[91],stage1_22[95],stage1_21[133],stage1_20[202]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[92],stage1_22[96],stage1_21[134],stage1_20[203]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[93],stage1_22[97],stage1_21[135],stage1_20[204]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[94],stage1_22[98],stage1_21[136],stage1_20[205]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[95],stage1_22[99],stage1_21[137],stage1_20[206]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[96],stage1_22[100],stage1_21[138],stage1_20[207]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[97],stage1_22[101],stage1_21[139],stage1_20[208]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[98],stage1_22[102],stage1_21[140],stage1_20[209]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[99],stage1_22[103],stage1_21[141],stage1_20[210]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[100],stage1_22[104],stage1_21[142],stage1_20[211]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[101],stage1_22[105],stage1_21[143],stage1_20[212]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291], stage0_22[292], stage0_22[293]},
      {stage1_24[48],stage1_23[102],stage1_22[106],stage1_21[144],stage1_20[213]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[294], stage0_22[295], stage0_22[296], stage0_22[297], stage0_22[298], stage0_22[299]},
      {stage1_24[49],stage1_23[103],stage1_22[107],stage1_21[145],stage1_20[214]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[300], stage0_22[301], stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305]},
      {stage1_24[50],stage1_23[104],stage1_22[108],stage1_21[146],stage1_20[215]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[306], stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage1_24[51],stage1_23[105],stage1_22[109],stage1_21[147],stage1_20[216]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316], stage0_22[317]},
      {stage1_24[52],stage1_23[106],stage1_22[110],stage1_21[148],stage1_20[217]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321], stage0_22[322], stage0_22[323]},
      {stage1_24[53],stage1_23[107],stage1_22[111],stage1_21[149],stage1_20[218]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[324], stage0_22[325], stage0_22[326], stage0_22[327], stage0_22[328], stage0_22[329]},
      {stage1_24[54],stage1_23[108],stage1_22[112],stage1_21[150],stage1_20[219]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[330], stage0_22[331], stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335]},
      {stage1_24[55],stage1_23[109],stage1_22[113],stage1_21[151],stage1_20[220]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[336], stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage1_24[56],stage1_23[110],stage1_22[114],stage1_21[152],stage1_20[221]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346], stage0_22[347]},
      {stage1_24[57],stage1_23[111],stage1_22[115],stage1_21[153],stage1_20[222]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351], stage0_22[352], stage0_22[353]},
      {stage1_24[58],stage1_23[112],stage1_22[116],stage1_21[154],stage1_20[223]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[354], stage0_22[355], stage0_22[356], stage0_22[357], stage0_22[358], stage0_22[359]},
      {stage1_24[59],stage1_23[113],stage1_22[117],stage1_21[155],stage1_20[224]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[360], stage0_22[361], stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365]},
      {stage1_24[60],stage1_23[114],stage1_22[118],stage1_21[156],stage1_20[225]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[366], stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage1_24[61],stage1_23[115],stage1_22[119],stage1_21[157],stage1_20[226]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376], stage0_22[377]},
      {stage1_24[62],stage1_23[116],stage1_22[120],stage1_21[158],stage1_20[227]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381], stage0_22[382], stage0_22[383]},
      {stage1_24[63],stage1_23[117],stage1_22[121],stage1_21[159],stage1_20[228]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[384], stage0_22[385], stage0_22[386], stage0_22[387], stage0_22[388], stage0_22[389]},
      {stage1_24[64],stage1_23[118],stage1_22[122],stage1_21[160],stage1_20[229]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[390], stage0_22[391], stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395]},
      {stage1_24[65],stage1_23[119],stage1_22[123],stage1_21[161],stage1_20[230]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[396], stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage1_24[66],stage1_23[120],stage1_22[124],stage1_21[162],stage1_20[231]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage1_24[67],stage1_23[121],stage1_22[125],stage1_21[163],stage1_20[232]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412], stage0_22[413]},
      {stage1_24[68],stage1_23[122],stage1_22[126],stage1_21[164],stage1_20[233]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417], stage0_22[418], stage0_22[419]},
      {stage1_24[69],stage1_23[123],stage1_22[127],stage1_21[165],stage1_20[234]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[420], stage0_22[421], stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425]},
      {stage1_24[70],stage1_23[124],stage1_22[128],stage1_21[166],stage1_20[235]}
   );
   gpc606_5 gpc876 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[71],stage1_23[125],stage1_22[129],stage1_21[167]}
   );
   gpc606_5 gpc877 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[72],stage1_23[126],stage1_22[130],stage1_21[168]}
   );
   gpc606_5 gpc878 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[73],stage1_23[127],stage1_22[131],stage1_21[169]}
   );
   gpc606_5 gpc879 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[74],stage1_23[128],stage1_22[132],stage1_21[170]}
   );
   gpc606_5 gpc880 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[75],stage1_23[129],stage1_22[133],stage1_21[171]}
   );
   gpc606_5 gpc881 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[76],stage1_23[130],stage1_22[134],stage1_21[172]}
   );
   gpc606_5 gpc882 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[77],stage1_23[131],stage1_22[135],stage1_21[173]}
   );
   gpc606_5 gpc883 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[78],stage1_23[132],stage1_22[136],stage1_21[174]}
   );
   gpc606_5 gpc884 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[79],stage1_23[133],stage1_22[137],stage1_21[175]}
   );
   gpc606_5 gpc885 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[80],stage1_23[134],stage1_22[138],stage1_21[176]}
   );
   gpc606_5 gpc886 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[81],stage1_23[135],stage1_22[139],stage1_21[177]}
   );
   gpc606_5 gpc887 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[82],stage1_23[136],stage1_22[140],stage1_21[178]}
   );
   gpc606_5 gpc888 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[83],stage1_23[137],stage1_22[141],stage1_21[179]}
   );
   gpc606_5 gpc889 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[84],stage1_23[138],stage1_22[142],stage1_21[180]}
   );
   gpc606_5 gpc890 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[85],stage1_23[139],stage1_22[143],stage1_21[181]}
   );
   gpc606_5 gpc891 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[86],stage1_23[140],stage1_22[144],stage1_21[182]}
   );
   gpc606_5 gpc892 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[87],stage1_23[141],stage1_22[145],stage1_21[183]}
   );
   gpc606_5 gpc893 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[88],stage1_23[142],stage1_22[146],stage1_21[184]}
   );
   gpc606_5 gpc894 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[89],stage1_23[143],stage1_22[147],stage1_21[185]}
   );
   gpc606_5 gpc895 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[90],stage1_23[144],stage1_22[148],stage1_21[186]}
   );
   gpc606_5 gpc896 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[91],stage1_23[145],stage1_22[149],stage1_21[187]}
   );
   gpc606_5 gpc897 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[92],stage1_23[146],stage1_22[150],stage1_21[188]}
   );
   gpc606_5 gpc898 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[93],stage1_23[147],stage1_22[151],stage1_21[189]}
   );
   gpc606_5 gpc899 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[94],stage1_23[148],stage1_22[152],stage1_21[190]}
   );
   gpc606_5 gpc900 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[95],stage1_23[149],stage1_22[153],stage1_21[191]}
   );
   gpc606_5 gpc901 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[96],stage1_23[150],stage1_22[154],stage1_21[192]}
   );
   gpc606_5 gpc902 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[97],stage1_23[151],stage1_22[155],stage1_21[193]}
   );
   gpc606_5 gpc903 (
      {stage0_21[486], stage0_21[487], stage0_21[488], stage0_21[489], stage0_21[490], stage0_21[491]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[98],stage1_23[152],stage1_22[156],stage1_21[194]}
   );
   gpc606_5 gpc904 (
      {stage0_21[492], stage0_21[493], stage0_21[494], stage0_21[495], stage0_21[496], stage0_21[497]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[99],stage1_23[153],stage1_22[157],stage1_21[195]}
   );
   gpc606_5 gpc905 (
      {stage0_21[498], stage0_21[499], stage0_21[500], stage0_21[501], stage0_21[502], stage0_21[503]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[100],stage1_23[154],stage1_22[158],stage1_21[196]}
   );
   gpc615_5 gpc906 (
      {stage0_22[426], stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430]},
      {stage0_23[180]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[30],stage1_24[101],stage1_23[155],stage1_22[159]}
   );
   gpc615_5 gpc907 (
      {stage0_22[431], stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435]},
      {stage0_23[181]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[31],stage1_24[102],stage1_23[156],stage1_22[160]}
   );
   gpc615_5 gpc908 (
      {stage0_22[436], stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440]},
      {stage0_23[182]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[32],stage1_24[103],stage1_23[157],stage1_22[161]}
   );
   gpc615_5 gpc909 (
      {stage0_22[441], stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445]},
      {stage0_23[183]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[33],stage1_24[104],stage1_23[158],stage1_22[162]}
   );
   gpc615_5 gpc910 (
      {stage0_22[446], stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450]},
      {stage0_23[184]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[34],stage1_24[105],stage1_23[159],stage1_22[163]}
   );
   gpc615_5 gpc911 (
      {stage0_22[451], stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455]},
      {stage0_23[185]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[35],stage1_24[106],stage1_23[160],stage1_22[164]}
   );
   gpc615_5 gpc912 (
      {stage0_22[456], stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460]},
      {stage0_23[186]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[36],stage1_24[107],stage1_23[161],stage1_22[165]}
   );
   gpc615_5 gpc913 (
      {stage0_22[461], stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465]},
      {stage0_23[187]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[37],stage1_24[108],stage1_23[162],stage1_22[166]}
   );
   gpc615_5 gpc914 (
      {stage0_22[466], stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470]},
      {stage0_23[188]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[38],stage1_24[109],stage1_23[163],stage1_22[167]}
   );
   gpc615_5 gpc915 (
      {stage0_22[471], stage0_22[472], stage0_22[473], stage0_22[474], stage0_22[475]},
      {stage0_23[189]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[39],stage1_24[110],stage1_23[164],stage1_22[168]}
   );
   gpc615_5 gpc916 (
      {stage0_22[476], stage0_22[477], stage0_22[478], stage0_22[479], stage0_22[480]},
      {stage0_23[190]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[40],stage1_24[111],stage1_23[165],stage1_22[169]}
   );
   gpc606_5 gpc917 (
      {stage0_23[191], stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[11],stage1_25[41],stage1_24[112],stage1_23[166]}
   );
   gpc606_5 gpc918 (
      {stage0_23[197], stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[12],stage1_25[42],stage1_24[113],stage1_23[167]}
   );
   gpc606_5 gpc919 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[13],stage1_25[43],stage1_24[114],stage1_23[168]}
   );
   gpc606_5 gpc920 (
      {stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[14],stage1_25[44],stage1_24[115],stage1_23[169]}
   );
   gpc606_5 gpc921 (
      {stage0_23[215], stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[15],stage1_25[45],stage1_24[116],stage1_23[170]}
   );
   gpc606_5 gpc922 (
      {stage0_23[221], stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[16],stage1_25[46],stage1_24[117],stage1_23[171]}
   );
   gpc606_5 gpc923 (
      {stage0_23[227], stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[17],stage1_25[47],stage1_24[118],stage1_23[172]}
   );
   gpc606_5 gpc924 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[18],stage1_25[48],stage1_24[119],stage1_23[173]}
   );
   gpc606_5 gpc925 (
      {stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[19],stage1_25[49],stage1_24[120],stage1_23[174]}
   );
   gpc606_5 gpc926 (
      {stage0_23[245], stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[20],stage1_25[50],stage1_24[121],stage1_23[175]}
   );
   gpc606_5 gpc927 (
      {stage0_23[251], stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[21],stage1_25[51],stage1_24[122],stage1_23[176]}
   );
   gpc606_5 gpc928 (
      {stage0_23[257], stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[22],stage1_25[52],stage1_24[123],stage1_23[177]}
   );
   gpc606_5 gpc929 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[23],stage1_25[53],stage1_24[124],stage1_23[178]}
   );
   gpc606_5 gpc930 (
      {stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[24],stage1_25[54],stage1_24[125],stage1_23[179]}
   );
   gpc606_5 gpc931 (
      {stage0_23[275], stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[25],stage1_25[55],stage1_24[126],stage1_23[180]}
   );
   gpc606_5 gpc932 (
      {stage0_23[281], stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[26],stage1_25[56],stage1_24[127],stage1_23[181]}
   );
   gpc606_5 gpc933 (
      {stage0_23[287], stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[27],stage1_25[57],stage1_24[128],stage1_23[182]}
   );
   gpc606_5 gpc934 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[28],stage1_25[58],stage1_24[129],stage1_23[183]}
   );
   gpc606_5 gpc935 (
      {stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[29],stage1_25[59],stage1_24[130],stage1_23[184]}
   );
   gpc606_5 gpc936 (
      {stage0_23[305], stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[30],stage1_25[60],stage1_24[131],stage1_23[185]}
   );
   gpc606_5 gpc937 (
      {stage0_23[311], stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[31],stage1_25[61],stage1_24[132],stage1_23[186]}
   );
   gpc606_5 gpc938 (
      {stage0_23[317], stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[32],stage1_25[62],stage1_24[133],stage1_23[187]}
   );
   gpc606_5 gpc939 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[33],stage1_25[63],stage1_24[134],stage1_23[188]}
   );
   gpc606_5 gpc940 (
      {stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[34],stage1_25[64],stage1_24[135],stage1_23[189]}
   );
   gpc606_5 gpc941 (
      {stage0_23[335], stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[35],stage1_25[65],stage1_24[136],stage1_23[190]}
   );
   gpc606_5 gpc942 (
      {stage0_23[341], stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[36],stage1_25[66],stage1_24[137],stage1_23[191]}
   );
   gpc606_5 gpc943 (
      {stage0_23[347], stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[37],stage1_25[67],stage1_24[138],stage1_23[192]}
   );
   gpc606_5 gpc944 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[38],stage1_25[68],stage1_24[139],stage1_23[193]}
   );
   gpc606_5 gpc945 (
      {stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[39],stage1_25[69],stage1_24[140],stage1_23[194]}
   );
   gpc606_5 gpc946 (
      {stage0_23[365], stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[40],stage1_25[70],stage1_24[141],stage1_23[195]}
   );
   gpc606_5 gpc947 (
      {stage0_23[371], stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[41],stage1_25[71],stage1_24[142],stage1_23[196]}
   );
   gpc606_5 gpc948 (
      {stage0_23[377], stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[42],stage1_25[72],stage1_24[143],stage1_23[197]}
   );
   gpc615_5 gpc949 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[66]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[43],stage1_25[73],stage1_24[144],stage1_23[198]}
   );
   gpc615_5 gpc950 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[67]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[44],stage1_25[74],stage1_24[145],stage1_23[199]}
   );
   gpc615_5 gpc951 (
      {stage0_23[393], stage0_23[394], stage0_23[395], stage0_23[396], stage0_23[397]},
      {stage0_24[68]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[45],stage1_25[75],stage1_24[146],stage1_23[200]}
   );
   gpc615_5 gpc952 (
      {stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401], stage0_23[402]},
      {stage0_24[69]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[46],stage1_25[76],stage1_24[147],stage1_23[201]}
   );
   gpc615_5 gpc953 (
      {stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage0_24[70]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[47],stage1_25[77],stage1_24[148],stage1_23[202]}
   );
   gpc615_5 gpc954 (
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412]},
      {stage0_24[71]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[48],stage1_25[78],stage1_24[149],stage1_23[203]}
   );
   gpc615_5 gpc955 (
      {stage0_23[413], stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417]},
      {stage0_24[72]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[49],stage1_25[79],stage1_24[150],stage1_23[204]}
   );
   gpc606_5 gpc956 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[39],stage1_26[50],stage1_25[80],stage1_24[151]}
   );
   gpc606_5 gpc957 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[40],stage1_26[51],stage1_25[81],stage1_24[152]}
   );
   gpc606_5 gpc958 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[41],stage1_26[52],stage1_25[82],stage1_24[153]}
   );
   gpc606_5 gpc959 (
      {stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[42],stage1_26[53],stage1_25[83],stage1_24[154]}
   );
   gpc606_5 gpc960 (
      {stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[43],stage1_26[54],stage1_25[84],stage1_24[155]}
   );
   gpc606_5 gpc961 (
      {stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[44],stage1_26[55],stage1_25[85],stage1_24[156]}
   );
   gpc606_5 gpc962 (
      {stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113], stage0_24[114]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[45],stage1_26[56],stage1_25[86],stage1_24[157]}
   );
   gpc606_5 gpc963 (
      {stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119], stage0_24[120]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[46],stage1_26[57],stage1_25[87],stage1_24[158]}
   );
   gpc606_5 gpc964 (
      {stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125], stage0_24[126]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[47],stage1_26[58],stage1_25[88],stage1_24[159]}
   );
   gpc606_5 gpc965 (
      {stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131], stage0_24[132]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[48],stage1_26[59],stage1_25[89],stage1_24[160]}
   );
   gpc606_5 gpc966 (
      {stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137], stage0_24[138]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[49],stage1_26[60],stage1_25[90],stage1_24[161]}
   );
   gpc606_5 gpc967 (
      {stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143], stage0_24[144]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[50],stage1_26[61],stage1_25[91],stage1_24[162]}
   );
   gpc606_5 gpc968 (
      {stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149], stage0_24[150]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[51],stage1_26[62],stage1_25[92],stage1_24[163]}
   );
   gpc606_5 gpc969 (
      {stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155], stage0_24[156]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[52],stage1_26[63],stage1_25[93],stage1_24[164]}
   );
   gpc606_5 gpc970 (
      {stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161], stage0_24[162]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[53],stage1_26[64],stage1_25[94],stage1_24[165]}
   );
   gpc606_5 gpc971 (
      {stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167], stage0_24[168]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[54],stage1_26[65],stage1_25[95],stage1_24[166]}
   );
   gpc606_5 gpc972 (
      {stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172], stage0_24[173], stage0_24[174]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[55],stage1_26[66],stage1_25[96],stage1_24[167]}
   );
   gpc606_5 gpc973 (
      {stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178], stage0_24[179], stage0_24[180]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[56],stage1_26[67],stage1_25[97],stage1_24[168]}
   );
   gpc606_5 gpc974 (
      {stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184], stage0_24[185], stage0_24[186]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[57],stage1_26[68],stage1_25[98],stage1_24[169]}
   );
   gpc606_5 gpc975 (
      {stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190], stage0_24[191], stage0_24[192]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[58],stage1_26[69],stage1_25[99],stage1_24[170]}
   );
   gpc606_5 gpc976 (
      {stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196], stage0_24[197], stage0_24[198]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[59],stage1_26[70],stage1_25[100],stage1_24[171]}
   );
   gpc606_5 gpc977 (
      {stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[60],stage1_26[71],stage1_25[101],stage1_24[172]}
   );
   gpc606_5 gpc978 (
      {stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[61],stage1_26[72],stage1_25[102],stage1_24[173]}
   );
   gpc606_5 gpc979 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215], stage0_24[216]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[62],stage1_26[73],stage1_25[103],stage1_24[174]}
   );
   gpc606_5 gpc980 (
      {stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220], stage0_24[221], stage0_24[222]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[63],stage1_26[74],stage1_25[104],stage1_24[175]}
   );
   gpc606_5 gpc981 (
      {stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226], stage0_24[227], stage0_24[228]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[64],stage1_26[75],stage1_25[105],stage1_24[176]}
   );
   gpc606_5 gpc982 (
      {stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[65],stage1_26[76],stage1_25[106],stage1_24[177]}
   );
   gpc606_5 gpc983 (
      {stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[66],stage1_26[77],stage1_25[107],stage1_24[178]}
   );
   gpc606_5 gpc984 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245], stage0_24[246]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[67],stage1_26[78],stage1_25[108],stage1_24[179]}
   );
   gpc606_5 gpc985 (
      {stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250], stage0_24[251], stage0_24[252]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[68],stage1_26[79],stage1_25[109],stage1_24[180]}
   );
   gpc606_5 gpc986 (
      {stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256], stage0_24[257], stage0_24[258]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[69],stage1_26[80],stage1_25[110],stage1_24[181]}
   );
   gpc606_5 gpc987 (
      {stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[70],stage1_26[81],stage1_25[111],stage1_24[182]}
   );
   gpc606_5 gpc988 (
      {stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[71],stage1_26[82],stage1_25[112],stage1_24[183]}
   );
   gpc606_5 gpc989 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275], stage0_24[276]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[72],stage1_26[83],stage1_25[113],stage1_24[184]}
   );
   gpc606_5 gpc990 (
      {stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280], stage0_24[281], stage0_24[282]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[73],stage1_26[84],stage1_25[114],stage1_24[185]}
   );
   gpc606_5 gpc991 (
      {stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286], stage0_24[287], stage0_24[288]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[74],stage1_26[85],stage1_25[115],stage1_24[186]}
   );
   gpc606_5 gpc992 (
      {stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[75],stage1_26[86],stage1_25[116],stage1_24[187]}
   );
   gpc606_5 gpc993 (
      {stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[76],stage1_26[87],stage1_25[117],stage1_24[188]}
   );
   gpc606_5 gpc994 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305], stage0_24[306]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[77],stage1_26[88],stage1_25[118],stage1_24[189]}
   );
   gpc606_5 gpc995 (
      {stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310], stage0_24[311], stage0_24[312]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[78],stage1_26[89],stage1_25[119],stage1_24[190]}
   );
   gpc606_5 gpc996 (
      {stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316], stage0_24[317], stage0_24[318]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[79],stage1_26[90],stage1_25[120],stage1_24[191]}
   );
   gpc606_5 gpc997 (
      {stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[80],stage1_26[91],stage1_25[121],stage1_24[192]}
   );
   gpc606_5 gpc998 (
      {stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[81],stage1_26[92],stage1_25[122],stage1_24[193]}
   );
   gpc606_5 gpc999 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335], stage0_24[336]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[82],stage1_26[93],stage1_25[123],stage1_24[194]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340], stage0_24[341], stage0_24[342]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[83],stage1_26[94],stage1_25[124],stage1_24[195]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346], stage0_24[347], stage0_24[348]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[84],stage1_26[95],stage1_25[125],stage1_24[196]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[85],stage1_26[96],stage1_25[126],stage1_24[197]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[86],stage1_26[97],stage1_25[127],stage1_24[198]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[87],stage1_26[98],stage1_25[128],stage1_24[199]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371], stage0_24[372]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[88],stage1_26[99],stage1_25[129],stage1_24[200]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376], stage0_24[377], stage0_24[378]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[89],stage1_26[100],stage1_25[130],stage1_24[201]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[90],stage1_26[101],stage1_25[131],stage1_24[202]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[91],stage1_26[102],stage1_25[132],stage1_24[203]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[92],stage1_26[103],stage1_25[133],stage1_24[204]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401], stage0_24[402]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[93],stage1_26[104],stage1_25[134],stage1_24[205]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406], stage0_24[407], stage0_24[408]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[94],stage1_26[105],stage1_25[135],stage1_24[206]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[95],stage1_26[106],stage1_25[136],stage1_24[207]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[96],stage1_26[107],stage1_25[137],stage1_24[208]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[97],stage1_26[108],stage1_25[138],stage1_24[209]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431], stage0_24[432]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[98],stage1_26[109],stage1_25[139],stage1_24[210]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436], stage0_24[437], stage0_24[438]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[99],stage1_26[110],stage1_25[140],stage1_24[211]}
   );
   gpc606_5 gpc1017 (
      {stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[100],stage1_26[111],stage1_25[141],stage1_24[212]}
   );
   gpc606_5 gpc1018 (
      {stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[101],stage1_26[112],stage1_25[142],stage1_24[213]}
   );
   gpc606_5 gpc1019 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[102],stage1_26[113],stage1_25[143],stage1_24[214]}
   );
   gpc606_5 gpc1020 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461], stage0_24[462]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[103],stage1_26[114],stage1_25[144],stage1_24[215]}
   );
   gpc606_5 gpc1021 (
      {stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466], stage0_24[467], stage0_24[468]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[104],stage1_26[115],stage1_25[145],stage1_24[216]}
   );
   gpc606_5 gpc1022 (
      {stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[105],stage1_26[116],stage1_25[146],stage1_24[217]}
   );
   gpc606_5 gpc1023 (
      {stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[106],stage1_26[117],stage1_25[147],stage1_24[218]}
   );
   gpc606_5 gpc1024 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[107],stage1_26[118],stage1_25[148],stage1_24[219]}
   );
   gpc606_5 gpc1025 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491], stage0_24[492]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[108],stage1_26[119],stage1_25[149],stage1_24[220]}
   );
   gpc606_5 gpc1026 (
      {stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496], stage0_24[497], stage0_24[498]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[109],stage1_26[120],stage1_25[150],stage1_24[221]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[71],stage1_27[110],stage1_26[121],stage1_25[151]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[72],stage1_27[111],stage1_26[122],stage1_25[152]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[426]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[73],stage1_27[112],stage1_26[123],stage1_25[153]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[427]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[74],stage1_27[113],stage1_26[124],stage1_25[154]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[428]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[75],stage1_27[114],stage1_26[125],stage1_25[155]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[429]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[76],stage1_27[115],stage1_26[126],stage1_25[156]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[430]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[77],stage1_27[116],stage1_26[127],stage1_25[157]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[431]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[78],stage1_27[117],stage1_26[128],stage1_25[158]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[432]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[79],stage1_27[118],stage1_26[129],stage1_25[159]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[433]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[80],stage1_27[119],stage1_26[130],stage1_25[160]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[434]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[81],stage1_27[120],stage1_26[131],stage1_25[161]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[435]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[82],stage1_27[121],stage1_26[132],stage1_25[162]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[436]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[83],stage1_27[122],stage1_26[133],stage1_25[163]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[437]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[84],stage1_27[123],stage1_26[134],stage1_25[164]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[438]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[85],stage1_27[124],stage1_26[135],stage1_25[165]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[439]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[86],stage1_27[125],stage1_26[136],stage1_25[166]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[440]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[87],stage1_27[126],stage1_26[137],stage1_25[167]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[441]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[88],stage1_27[127],stage1_26[138],stage1_25[168]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[442]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[89],stage1_27[128],stage1_26[139],stage1_25[169]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[443]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[90],stage1_27[129],stage1_26[140],stage1_25[170]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[444]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[91],stage1_27[130],stage1_26[141],stage1_25[171]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[445]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[92],stage1_27[131],stage1_26[142],stage1_25[172]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[446]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[93],stage1_27[132],stage1_26[143],stage1_25[173]}
   );
   gpc615_5 gpc1050 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[447]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[94],stage1_27[133],stage1_26[144],stage1_25[174]}
   );
   gpc615_5 gpc1051 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[448]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[95],stage1_27[134],stage1_26[145],stage1_25[175]}
   );
   gpc615_5 gpc1052 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[449]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[96],stage1_27[135],stage1_26[146],stage1_25[176]}
   );
   gpc615_5 gpc1053 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[450]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[97],stage1_27[136],stage1_26[147],stage1_25[177]}
   );
   gpc615_5 gpc1054 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[451]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[98],stage1_27[137],stage1_26[148],stage1_25[178]}
   );
   gpc615_5 gpc1055 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[452]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[99],stage1_27[138],stage1_26[149],stage1_25[179]}
   );
   gpc615_5 gpc1056 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[453]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[100],stage1_27[139],stage1_26[150],stage1_25[180]}
   );
   gpc615_5 gpc1057 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[454]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[101],stage1_27[140],stage1_26[151],stage1_25[181]}
   );
   gpc615_5 gpc1058 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[455]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[102],stage1_27[141],stage1_26[152],stage1_25[182]}
   );
   gpc615_5 gpc1059 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[456]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[103],stage1_27[142],stage1_26[153],stage1_25[183]}
   );
   gpc615_5 gpc1060 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[457]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[104],stage1_27[143],stage1_26[154],stage1_25[184]}
   );
   gpc615_5 gpc1061 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[458]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[105],stage1_27[144],stage1_26[155],stage1_25[185]}
   );
   gpc615_5 gpc1062 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[459]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[106],stage1_27[145],stage1_26[156],stage1_25[186]}
   );
   gpc615_5 gpc1063 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[460]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[107],stage1_27[146],stage1_26[157],stage1_25[187]}
   );
   gpc615_5 gpc1064 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[461]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[108],stage1_27[147],stage1_26[158],stage1_25[188]}
   );
   gpc615_5 gpc1065 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[462]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[109],stage1_27[148],stage1_26[159],stage1_25[189]}
   );
   gpc615_5 gpc1066 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[463]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[110],stage1_27[149],stage1_26[160],stage1_25[190]}
   );
   gpc615_5 gpc1067 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[464]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[111],stage1_27[150],stage1_26[161],stage1_25[191]}
   );
   gpc615_5 gpc1068 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[465]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[112],stage1_27[151],stage1_26[162],stage1_25[192]}
   );
   gpc615_5 gpc1069 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[466]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[113],stage1_27[152],stage1_26[163],stage1_25[193]}
   );
   gpc615_5 gpc1070 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[467]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[114],stage1_27[153],stage1_26[164],stage1_25[194]}
   );
   gpc615_5 gpc1071 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[468]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[115],stage1_27[154],stage1_26[165],stage1_25[195]}
   );
   gpc615_5 gpc1072 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[469]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[116],stage1_27[155],stage1_26[166],stage1_25[196]}
   );
   gpc615_5 gpc1073 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[470]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[117],stage1_27[156],stage1_26[167],stage1_25[197]}
   );
   gpc615_5 gpc1074 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[471]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[118],stage1_27[157],stage1_26[168],stage1_25[198]}
   );
   gpc615_5 gpc1075 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[472]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[119],stage1_27[158],stage1_26[169],stage1_25[199]}
   );
   gpc615_5 gpc1076 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[473]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[120],stage1_27[159],stage1_26[170],stage1_25[200]}
   );
   gpc615_5 gpc1077 (
      {stage0_25[486], stage0_25[487], stage0_25[488], stage0_25[489], stage0_25[490]},
      {stage0_26[474]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[121],stage1_27[160],stage1_26[171],stage1_25[201]}
   );
   gpc615_5 gpc1078 (
      {stage0_25[491], stage0_25[492], stage0_25[493], stage0_25[494], stage0_25[495]},
      {stage0_26[475]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[122],stage1_27[161],stage1_26[172],stage1_25[202]}
   );
   gpc615_5 gpc1079 (
      {stage0_25[496], stage0_25[497], stage0_25[498], stage0_25[499], stage0_25[500]},
      {stage0_26[476]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[123],stage1_27[162],stage1_26[173],stage1_25[203]}
   );
   gpc615_5 gpc1080 (
      {stage0_25[501], stage0_25[502], stage0_25[503], stage0_25[504], stage0_25[505]},
      {stage0_26[477]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[124],stage1_27[163],stage1_26[174],stage1_25[204]}
   );
   gpc615_5 gpc1081 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[324]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[54],stage1_28[125],stage1_27[164],stage1_26[175]}
   );
   gpc615_5 gpc1082 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[325]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[55],stage1_28[126],stage1_27[165],stage1_26[176]}
   );
   gpc615_5 gpc1083 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[326]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[56],stage1_28[127],stage1_27[166],stage1_26[177]}
   );
   gpc615_5 gpc1084 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[327]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[57],stage1_28[128],stage1_27[167],stage1_26[178]}
   );
   gpc615_5 gpc1085 (
      {stage0_26[498], stage0_26[499], stage0_26[500], stage0_26[501], stage0_26[502]},
      {stage0_27[328]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[58],stage1_28[129],stage1_27[168],stage1_26[179]}
   );
   gpc7_3 gpc1086 (
      {stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[59],stage1_28[130],stage1_27[169]}
   );
   gpc7_3 gpc1087 (
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage1_29[60],stage1_28[131],stage1_27[170]}
   );
   gpc615_5 gpc1088 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[30]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[61],stage1_28[132],stage1_27[171]}
   );
   gpc615_5 gpc1089 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[31]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[62],stage1_28[133],stage1_27[172]}
   );
   gpc615_5 gpc1090 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[32]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[63],stage1_28[134],stage1_27[173]}
   );
   gpc615_5 gpc1091 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[33]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[64],stage1_28[135],stage1_27[174]}
   );
   gpc615_5 gpc1092 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[34]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[65],stage1_28[136],stage1_27[175]}
   );
   gpc615_5 gpc1093 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[35]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[66],stage1_28[137],stage1_27[176]}
   );
   gpc615_5 gpc1094 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[36]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[67],stage1_28[138],stage1_27[177]}
   );
   gpc615_5 gpc1095 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[37]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[68],stage1_28[139],stage1_27[178]}
   );
   gpc615_5 gpc1096 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[38]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[69],stage1_28[140],stage1_27[179]}
   );
   gpc615_5 gpc1097 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[39]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[70],stage1_28[141],stage1_27[180]}
   );
   gpc615_5 gpc1098 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[40]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[15],stage1_29[71],stage1_28[142],stage1_27[181]}
   );
   gpc615_5 gpc1099 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[41]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[16],stage1_29[72],stage1_28[143],stage1_27[182]}
   );
   gpc615_5 gpc1100 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[42]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[17],stage1_29[73],stage1_28[144],stage1_27[183]}
   );
   gpc615_5 gpc1101 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[43]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[18],stage1_29[74],stage1_28[145],stage1_27[184]}
   );
   gpc615_5 gpc1102 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[44]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[19],stage1_29[75],stage1_28[146],stage1_27[185]}
   );
   gpc615_5 gpc1103 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[45]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[20],stage1_29[76],stage1_28[147],stage1_27[186]}
   );
   gpc615_5 gpc1104 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[46]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[21],stage1_29[77],stage1_28[148],stage1_27[187]}
   );
   gpc615_5 gpc1105 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[47]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[22],stage1_29[78],stage1_28[149],stage1_27[188]}
   );
   gpc615_5 gpc1106 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[48]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[23],stage1_29[79],stage1_28[150],stage1_27[189]}
   );
   gpc615_5 gpc1107 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[49]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[24],stage1_29[80],stage1_28[151],stage1_27[190]}
   );
   gpc615_5 gpc1108 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[50]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[25],stage1_29[81],stage1_28[152],stage1_27[191]}
   );
   gpc615_5 gpc1109 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[51]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[26],stage1_29[82],stage1_28[153],stage1_27[192]}
   );
   gpc615_5 gpc1110 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[52]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[27],stage1_29[83],stage1_28[154],stage1_27[193]}
   );
   gpc615_5 gpc1111 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[53]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[28],stage1_29[84],stage1_28[155],stage1_27[194]}
   );
   gpc615_5 gpc1112 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[54]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[29],stage1_29[85],stage1_28[156],stage1_27[195]}
   );
   gpc615_5 gpc1113 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[55]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[30],stage1_29[86],stage1_28[157],stage1_27[196]}
   );
   gpc615_5 gpc1114 (
      {stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477]},
      {stage0_28[56]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[31],stage1_29[87],stage1_28[158],stage1_27[197]}
   );
   gpc615_5 gpc1115 (
      {stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_28[57]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[32],stage1_29[88],stage1_28[159],stage1_27[198]}
   );
   gpc615_5 gpc1116 (
      {stage0_27[483], stage0_27[484], stage0_27[485], stage0_27[486], stage0_27[487]},
      {stage0_28[58]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[33],stage1_29[89],stage1_28[160],stage1_27[199]}
   );
   gpc615_5 gpc1117 (
      {stage0_27[488], stage0_27[489], stage0_27[490], stage0_27[491], stage0_27[492]},
      {stage0_28[59]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[34],stage1_29[90],stage1_28[161],stage1_27[200]}
   );
   gpc615_5 gpc1118 (
      {stage0_27[493], stage0_27[494], stage0_27[495], stage0_27[496], stage0_27[497]},
      {stage0_28[60]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[35],stage1_29[91],stage1_28[162],stage1_27[201]}
   );
   gpc615_5 gpc1119 (
      {stage0_27[498], stage0_27[499], stage0_27[500], stage0_27[501], stage0_27[502]},
      {stage0_28[61]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[36],stage1_29[92],stage1_28[163],stage1_27[202]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65], stage0_28[66], stage0_28[67]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[32],stage1_30[37],stage1_29[93],stage1_28[164]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71], stage0_28[72], stage0_28[73]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[33],stage1_30[38],stage1_29[94],stage1_28[165]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78], stage0_28[79]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[34],stage1_30[39],stage1_29[95],stage1_28[166]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84], stage0_28[85]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[35],stage1_30[40],stage1_29[96],stage1_28[167]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90], stage0_28[91]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[36],stage1_30[41],stage1_29[97],stage1_28[168]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[37],stage1_30[42],stage1_29[98],stage1_28[169]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[38],stage1_30[43],stage1_29[99],stage1_28[170]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[39],stage1_30[44],stage1_29[100],stage1_28[171]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[40],stage1_30[45],stage1_29[101],stage1_28[172]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[41],stage1_30[46],stage1_29[102],stage1_28[173]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[42],stage1_30[47],stage1_29[103],stage1_28[174]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[43],stage1_30[48],stage1_29[104],stage1_28[175]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[44],stage1_30[49],stage1_29[105],stage1_28[176]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144], stage0_28[145]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[45],stage1_30[50],stage1_29[106],stage1_28[177]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150], stage0_28[151]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[46],stage1_30[51],stage1_29[107],stage1_28[178]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156], stage0_28[157]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[47],stage1_30[52],stage1_29[108],stage1_28[179]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162], stage0_28[163]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[48],stage1_30[53],stage1_29[109],stage1_28[180]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168], stage0_28[169]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[49],stage1_30[54],stage1_29[110],stage1_28[181]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174], stage0_28[175]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[50],stage1_30[55],stage1_29[111],stage1_28[182]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180], stage0_28[181]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[51],stage1_30[56],stage1_29[112],stage1_28[183]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186], stage0_28[187]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[52],stage1_30[57],stage1_29[113],stage1_28[184]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192], stage0_28[193]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[53],stage1_30[58],stage1_29[114],stage1_28[185]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198], stage0_28[199]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[54],stage1_30[59],stage1_29[115],stage1_28[186]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204], stage0_28[205]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[55],stage1_30[60],stage1_29[116],stage1_28[187]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210], stage0_28[211]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[56],stage1_30[61],stage1_29[117],stage1_28[188]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216], stage0_28[217]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[57],stage1_30[62],stage1_29[118],stage1_28[189]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222], stage0_28[223]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[58],stage1_30[63],stage1_29[119],stage1_28[190]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228], stage0_28[229]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[59],stage1_30[64],stage1_29[120],stage1_28[191]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234], stage0_28[235]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[60],stage1_30[65],stage1_29[121],stage1_28[192]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240], stage0_28[241]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[61],stage1_30[66],stage1_29[122],stage1_28[193]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246], stage0_28[247]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[62],stage1_30[67],stage1_29[123],stage1_28[194]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252], stage0_28[253]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[63],stage1_30[68],stage1_29[124],stage1_28[195]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258], stage0_28[259]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[64],stage1_30[69],stage1_29[125],stage1_28[196]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264], stage0_28[265]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[65],stage1_30[70],stage1_29[126],stage1_28[197]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270], stage0_28[271]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[66],stage1_30[71],stage1_29[127],stage1_28[198]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276], stage0_28[277]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[67],stage1_30[72],stage1_29[128],stage1_28[199]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282], stage0_28[283]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[68],stage1_30[73],stage1_29[129],stage1_28[200]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288], stage0_28[289]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[69],stage1_30[74],stage1_29[130],stage1_28[201]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294], stage0_28[295]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[70],stage1_30[75],stage1_29[131],stage1_28[202]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300], stage0_28[301]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[71],stage1_30[76],stage1_29[132],stage1_28[203]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306], stage0_28[307]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[72],stage1_30[77],stage1_29[133],stage1_28[204]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312], stage0_28[313]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[73],stage1_30[78],stage1_29[134],stage1_28[205]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[74],stage1_30[79],stage1_29[135],stage1_28[206]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[75],stage1_30[80],stage1_29[136],stage1_28[207]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330], stage0_28[331]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[76],stage1_30[81],stage1_29[137],stage1_28[208]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336], stage0_28[337]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[77],stage1_30[82],stage1_29[138],stage1_28[209]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342], stage0_28[343]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[78],stage1_30[83],stage1_29[139],stage1_28[210]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[79],stage1_30[84],stage1_29[140],stage1_28[211]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[80],stage1_30[85],stage1_29[141],stage1_28[212]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360], stage0_28[361]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[81],stage1_30[86],stage1_29[142],stage1_28[213]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366], stage0_28[367]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[82],stage1_30[87],stage1_29[143],stage1_28[214]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372], stage0_28[373]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[83],stage1_30[88],stage1_29[144],stage1_28[215]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[84],stage1_30[89],stage1_29[145],stage1_28[216]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[85],stage1_30[90],stage1_29[146],stage1_28[217]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390], stage0_28[391]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[86],stage1_30[91],stage1_29[147],stage1_28[218]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396], stage0_28[397]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[87],stage1_30[92],stage1_29[148],stage1_28[219]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402], stage0_28[403]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[88],stage1_30[93],stage1_29[149],stage1_28[220]}
   );
   gpc606_5 gpc1177 (
      {stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[89],stage1_30[94],stage1_29[150],stage1_28[221]}
   );
   gpc606_5 gpc1178 (
      {stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[90],stage1_30[95],stage1_29[151],stage1_28[222]}
   );
   gpc606_5 gpc1179 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420], stage0_28[421]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[91],stage1_30[96],stage1_29[152],stage1_28[223]}
   );
   gpc606_5 gpc1180 (
      {stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426], stage0_28[427]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[92],stage1_30[97],stage1_29[153],stage1_28[224]}
   );
   gpc606_5 gpc1181 (
      {stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432], stage0_28[433]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[93],stage1_30[98],stage1_29[154],stage1_28[225]}
   );
   gpc606_5 gpc1182 (
      {stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[94],stage1_30[99],stage1_29[155],stage1_28[226]}
   );
   gpc606_5 gpc1183 (
      {stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[95],stage1_30[100],stage1_29[156],stage1_28[227]}
   );
   gpc606_5 gpc1184 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450], stage0_28[451]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[96],stage1_30[101],stage1_29[157],stage1_28[228]}
   );
   gpc606_5 gpc1185 (
      {stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456], stage0_28[457]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[97],stage1_30[102],stage1_29[158],stage1_28[229]}
   );
   gpc606_5 gpc1186 (
      {stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462], stage0_28[463]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[98],stage1_30[103],stage1_29[159],stage1_28[230]}
   );
   gpc606_5 gpc1187 (
      {stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[99],stage1_30[104],stage1_29[160],stage1_28[231]}
   );
   gpc606_5 gpc1188 (
      {stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[100],stage1_30[105],stage1_29[161],stage1_28[232]}
   );
   gpc606_5 gpc1189 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480], stage0_28[481]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[101],stage1_30[106],stage1_29[162],stage1_28[233]}
   );
   gpc606_5 gpc1190 (
      {stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485], stage0_28[486], stage0_28[487]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[102],stage1_30[107],stage1_29[163],stage1_28[234]}
   );
   gpc606_5 gpc1191 (
      {stage0_28[488], stage0_28[489], stage0_28[490], stage0_28[491], stage0_28[492], stage0_28[493]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[103],stage1_30[108],stage1_29[164],stage1_28[235]}
   );
   gpc606_5 gpc1192 (
      {stage0_28[494], stage0_28[495], stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[104],stage1_30[109],stage1_29[165],stage1_28[236]}
   );
   gpc606_5 gpc1193 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[73],stage1_31[105],stage1_30[110],stage1_29[166]}
   );
   gpc606_5 gpc1194 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[74],stage1_31[106],stage1_30[111],stage1_29[167]}
   );
   gpc606_5 gpc1195 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[75],stage1_31[107],stage1_30[112],stage1_29[168]}
   );
   gpc606_5 gpc1196 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[76],stage1_31[108],stage1_30[113],stage1_29[169]}
   );
   gpc606_5 gpc1197 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[77],stage1_31[109],stage1_30[114],stage1_29[170]}
   );
   gpc606_5 gpc1198 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[78],stage1_31[110],stage1_30[115],stage1_29[171]}
   );
   gpc606_5 gpc1199 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[79],stage1_31[111],stage1_30[116],stage1_29[172]}
   );
   gpc606_5 gpc1200 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[80],stage1_31[112],stage1_30[117],stage1_29[173]}
   );
   gpc606_5 gpc1201 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[81],stage1_31[113],stage1_30[118],stage1_29[174]}
   );
   gpc606_5 gpc1202 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[82],stage1_31[114],stage1_30[119],stage1_29[175]}
   );
   gpc606_5 gpc1203 (
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[83],stage1_31[115],stage1_30[120],stage1_29[176]}
   );
   gpc606_5 gpc1204 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[84],stage1_31[116],stage1_30[121],stage1_29[177]}
   );
   gpc606_5 gpc1205 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[85],stage1_31[117],stage1_30[122],stage1_29[178]}
   );
   gpc606_5 gpc1206 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[86],stage1_31[118],stage1_30[123],stage1_29[179]}
   );
   gpc606_5 gpc1207 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[87],stage1_31[119],stage1_30[124],stage1_29[180]}
   );
   gpc606_5 gpc1208 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[88],stage1_31[120],stage1_30[125],stage1_29[181]}
   );
   gpc606_5 gpc1209 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[89],stage1_31[121],stage1_30[126],stage1_29[182]}
   );
   gpc606_5 gpc1210 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[90],stage1_31[122],stage1_30[127],stage1_29[183]}
   );
   gpc606_5 gpc1211 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[91],stage1_31[123],stage1_30[128],stage1_29[184]}
   );
   gpc606_5 gpc1212 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[92],stage1_31[124],stage1_30[129],stage1_29[185]}
   );
   gpc606_5 gpc1213 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[93],stage1_31[125],stage1_30[130],stage1_29[186]}
   );
   gpc606_5 gpc1214 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[94],stage1_31[126],stage1_30[131],stage1_29[187]}
   );
   gpc606_5 gpc1215 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[95],stage1_31[127],stage1_30[132],stage1_29[188]}
   );
   gpc606_5 gpc1216 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[96],stage1_31[128],stage1_30[133],stage1_29[189]}
   );
   gpc606_5 gpc1217 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[97],stage1_31[129],stage1_30[134],stage1_29[190]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[98],stage1_31[130],stage1_30[135],stage1_29[191]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[99],stage1_31[131],stage1_30[136],stage1_29[192]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[100],stage1_31[132],stage1_30[137],stage1_29[193]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[101],stage1_31[133],stage1_30[138],stage1_29[194]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[102],stage1_31[134],stage1_30[139],stage1_29[195]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[103],stage1_31[135],stage1_30[140],stage1_29[196]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[104],stage1_31[136],stage1_30[141],stage1_29[197]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[105],stage1_31[137],stage1_30[142],stage1_29[198]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[106],stage1_31[138],stage1_30[143],stage1_29[199]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[107],stage1_31[139],stage1_30[144],stage1_29[200]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[108],stage1_31[140],stage1_30[145],stage1_29[201]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[109],stage1_31[141],stage1_30[146],stage1_29[202]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[110],stage1_31[142],stage1_30[147],stage1_29[203]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[111],stage1_31[143],stage1_30[148],stage1_29[204]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[112],stage1_31[144],stage1_30[149],stage1_29[205]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[113],stage1_31[145],stage1_30[150],stage1_29[206]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[114],stage1_31[146],stage1_30[151],stage1_29[207]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[115],stage1_31[147],stage1_30[152],stage1_29[208]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[116],stage1_31[148],stage1_30[153],stage1_29[209]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460], stage0_29[461]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[117],stage1_31[149],stage1_30[154],stage1_29[210]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466], stage0_29[467]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[118],stage1_31[150],stage1_30[155],stage1_29[211]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472], stage0_29[473]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[119],stage1_31[151],stage1_30[156],stage1_29[212]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[120],stage1_31[152],stage1_30[157],stage1_29[213]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[121],stage1_31[153],stage1_30[158],stage1_29[214]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490], stage0_29[491]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[122],stage1_31[154],stage1_30[159],stage1_29[215]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496], stage0_29[497]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[123],stage1_31[155],stage1_30[160],stage1_29[216]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502], stage0_29[503]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[124],stage1_31[156],stage1_30[161],stage1_29[217]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508], stage0_29[509]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[125],stage1_31[157],stage1_30[162],stage1_29[218]}
   );
   gpc1415_5 gpc1246 (
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442]},
      {stage0_31[318]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[53],stage1_32[126],stage1_31[158],stage1_30[163]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage0_32[4]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[1],stage1_33[54],stage1_32[127],stage1_31[159]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328]},
      {stage0_32[5]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[2],stage1_33[55],stage1_32[128],stage1_31[160]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[329], stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333]},
      {stage0_32[6]},
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage1_35[2],stage1_34[3],stage1_33[56],stage1_32[129],stage1_31[161]}
   );
   gpc615_5 gpc1250 (
      {stage0_31[334], stage0_31[335], stage0_31[336], stage0_31[337], stage0_31[338]},
      {stage0_32[7]},
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage1_35[3],stage1_34[4],stage1_33[57],stage1_32[130],stage1_31[162]}
   );
   gpc615_5 gpc1251 (
      {stage0_31[339], stage0_31[340], stage0_31[341], stage0_31[342], stage0_31[343]},
      {stage0_32[8]},
      {stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29], stage0_33[30]},
      {stage1_35[4],stage1_34[5],stage1_33[58],stage1_32[131],stage1_31[163]}
   );
   gpc615_5 gpc1252 (
      {stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347], stage0_31[348]},
      {stage0_32[9]},
      {stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35], stage0_33[36]},
      {stage1_35[5],stage1_34[6],stage1_33[59],stage1_32[132],stage1_31[164]}
   );
   gpc615_5 gpc1253 (
      {stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage0_32[10]},
      {stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41], stage0_33[42]},
      {stage1_35[6],stage1_34[7],stage1_33[60],stage1_32[133],stage1_31[165]}
   );
   gpc615_5 gpc1254 (
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358]},
      {stage0_32[11]},
      {stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47], stage0_33[48]},
      {stage1_35[7],stage1_34[8],stage1_33[61],stage1_32[134],stage1_31[166]}
   );
   gpc615_5 gpc1255 (
      {stage0_31[359], stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363]},
      {stage0_32[12]},
      {stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53], stage0_33[54]},
      {stage1_35[8],stage1_34[9],stage1_33[62],stage1_32[135],stage1_31[167]}
   );
   gpc615_5 gpc1256 (
      {stage0_31[364], stage0_31[365], stage0_31[366], stage0_31[367], stage0_31[368]},
      {stage0_32[13]},
      {stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59], stage0_33[60]},
      {stage1_35[9],stage1_34[10],stage1_33[63],stage1_32[136],stage1_31[168]}
   );
   gpc615_5 gpc1257 (
      {stage0_31[369], stage0_31[370], stage0_31[371], stage0_31[372], stage0_31[373]},
      {stage0_32[14]},
      {stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65], stage0_33[66]},
      {stage1_35[10],stage1_34[11],stage1_33[64],stage1_32[137],stage1_31[169]}
   );
   gpc615_5 gpc1258 (
      {stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377], stage0_31[378]},
      {stage0_32[15]},
      {stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71], stage0_33[72]},
      {stage1_35[11],stage1_34[12],stage1_33[65],stage1_32[138],stage1_31[170]}
   );
   gpc615_5 gpc1259 (
      {stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage0_32[16]},
      {stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77], stage0_33[78]},
      {stage1_35[12],stage1_34[13],stage1_33[66],stage1_32[139],stage1_31[171]}
   );
   gpc615_5 gpc1260 (
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388]},
      {stage0_32[17]},
      {stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83], stage0_33[84]},
      {stage1_35[13],stage1_34[14],stage1_33[67],stage1_32[140],stage1_31[172]}
   );
   gpc615_5 gpc1261 (
      {stage0_31[389], stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393]},
      {stage0_32[18]},
      {stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89], stage0_33[90]},
      {stage1_35[14],stage1_34[15],stage1_33[68],stage1_32[141],stage1_31[173]}
   );
   gpc615_5 gpc1262 (
      {stage0_31[394], stage0_31[395], stage0_31[396], stage0_31[397], stage0_31[398]},
      {stage0_32[19]},
      {stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95], stage0_33[96]},
      {stage1_35[15],stage1_34[16],stage1_33[69],stage1_32[142],stage1_31[174]}
   );
   gpc615_5 gpc1263 (
      {stage0_31[399], stage0_31[400], stage0_31[401], stage0_31[402], stage0_31[403]},
      {stage0_32[20]},
      {stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101], stage0_33[102]},
      {stage1_35[16],stage1_34[17],stage1_33[70],stage1_32[143],stage1_31[175]}
   );
   gpc615_5 gpc1264 (
      {stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407], stage0_31[408]},
      {stage0_32[21]},
      {stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107], stage0_33[108]},
      {stage1_35[17],stage1_34[18],stage1_33[71],stage1_32[144],stage1_31[176]}
   );
   gpc615_5 gpc1265 (
      {stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage0_32[22]},
      {stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113], stage0_33[114]},
      {stage1_35[18],stage1_34[19],stage1_33[72],stage1_32[145],stage1_31[177]}
   );
   gpc615_5 gpc1266 (
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418]},
      {stage0_32[23]},
      {stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119], stage0_33[120]},
      {stage1_35[19],stage1_34[20],stage1_33[73],stage1_32[146],stage1_31[178]}
   );
   gpc615_5 gpc1267 (
      {stage0_31[419], stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423]},
      {stage0_32[24]},
      {stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125], stage0_33[126]},
      {stage1_35[20],stage1_34[21],stage1_33[74],stage1_32[147],stage1_31[179]}
   );
   gpc615_5 gpc1268 (
      {stage0_31[424], stage0_31[425], stage0_31[426], stage0_31[427], stage0_31[428]},
      {stage0_32[25]},
      {stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131], stage0_33[132]},
      {stage1_35[21],stage1_34[22],stage1_33[75],stage1_32[148],stage1_31[180]}
   );
   gpc615_5 gpc1269 (
      {stage0_31[429], stage0_31[430], stage0_31[431], stage0_31[432], stage0_31[433]},
      {stage0_32[26]},
      {stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137], stage0_33[138]},
      {stage1_35[22],stage1_34[23],stage1_33[76],stage1_32[149],stage1_31[181]}
   );
   gpc615_5 gpc1270 (
      {stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437], stage0_31[438]},
      {stage0_32[27]},
      {stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143], stage0_33[144]},
      {stage1_35[23],stage1_34[24],stage1_33[77],stage1_32[150],stage1_31[182]}
   );
   gpc615_5 gpc1271 (
      {stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage0_32[28]},
      {stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149], stage0_33[150]},
      {stage1_35[24],stage1_34[25],stage1_33[78],stage1_32[151],stage1_31[183]}
   );
   gpc615_5 gpc1272 (
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448]},
      {stage0_32[29]},
      {stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155], stage0_33[156]},
      {stage1_35[25],stage1_34[26],stage1_33[79],stage1_32[152],stage1_31[184]}
   );
   gpc615_5 gpc1273 (
      {stage0_31[449], stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453]},
      {stage0_32[30]},
      {stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161], stage0_33[162]},
      {stage1_35[26],stage1_34[27],stage1_33[80],stage1_32[153],stage1_31[185]}
   );
   gpc615_5 gpc1274 (
      {stage0_31[454], stage0_31[455], stage0_31[456], stage0_31[457], stage0_31[458]},
      {stage0_32[31]},
      {stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167], stage0_33[168]},
      {stage1_35[27],stage1_34[28],stage1_33[81],stage1_32[154],stage1_31[186]}
   );
   gpc615_5 gpc1275 (
      {stage0_31[459], stage0_31[460], stage0_31[461], stage0_31[462], stage0_31[463]},
      {stage0_32[32]},
      {stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173], stage0_33[174]},
      {stage1_35[28],stage1_34[29],stage1_33[82],stage1_32[155],stage1_31[187]}
   );
   gpc615_5 gpc1276 (
      {stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467], stage0_31[468]},
      {stage0_32[33]},
      {stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179], stage0_33[180]},
      {stage1_35[29],stage1_34[30],stage1_33[83],stage1_32[156],stage1_31[188]}
   );
   gpc615_5 gpc1277 (
      {stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage0_32[34]},
      {stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185], stage0_33[186]},
      {stage1_35[30],stage1_34[31],stage1_33[84],stage1_32[157],stage1_31[189]}
   );
   gpc615_5 gpc1278 (
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478]},
      {stage0_32[35]},
      {stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191], stage0_33[192]},
      {stage1_35[31],stage1_34[32],stage1_33[85],stage1_32[158],stage1_31[190]}
   );
   gpc615_5 gpc1279 (
      {stage0_31[479], stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483]},
      {stage0_32[36]},
      {stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197], stage0_33[198]},
      {stage1_35[32],stage1_34[33],stage1_33[86],stage1_32[159],stage1_31[191]}
   );
   gpc615_5 gpc1280 (
      {stage0_31[484], stage0_31[485], stage0_31[486], stage0_31[487], stage0_31[488]},
      {stage0_32[37]},
      {stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203], stage0_33[204]},
      {stage1_35[33],stage1_34[34],stage1_33[87],stage1_32[160],stage1_31[192]}
   );
   gpc615_5 gpc1281 (
      {stage0_31[489], stage0_31[490], stage0_31[491], stage0_31[492], stage0_31[493]},
      {stage0_32[38]},
      {stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209], stage0_33[210]},
      {stage1_35[34],stage1_34[35],stage1_33[88],stage1_32[161],stage1_31[193]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[35],stage1_34[36],stage1_33[89],stage1_32[162]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[36],stage1_34[37],stage1_33[90],stage1_32[163]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[37],stage1_34[38],stage1_33[91],stage1_32[164]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[38],stage1_34[39],stage1_33[92],stage1_32[165]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[63], stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[39],stage1_34[40],stage1_33[93],stage1_32[166]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73], stage0_32[74]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[40],stage1_34[41],stage1_33[94],stage1_32[167]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78], stage0_32[79], stage0_32[80]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[41],stage1_34[42],stage1_33[95],stage1_32[168]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[81], stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[42],stage1_34[43],stage1_33[96],stage1_32[169]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[87], stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[43],stage1_34[44],stage1_33[97],stage1_32[170]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[93], stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[44],stage1_34[45],stage1_33[98],stage1_32[171]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103], stage0_32[104]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[45],stage1_34[46],stage1_33[99],stage1_32[172]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108], stage0_32[109], stage0_32[110]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[46],stage1_34[47],stage1_33[100],stage1_32[173]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[111], stage0_32[112], stage0_32[113], stage0_32[114], stage0_32[115], stage0_32[116]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[47],stage1_34[48],stage1_33[101],stage1_32[174]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[117], stage0_32[118], stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[48],stage1_34[49],stage1_33[102],stage1_32[175]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[123], stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[49],stage1_34[50],stage1_33[103],stage1_32[176]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[129], stage0_32[130], stage0_32[131], stage0_32[132], stage0_32[133], stage0_32[134]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[50],stage1_34[51],stage1_33[104],stage1_32[177]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[135], stage0_32[136], stage0_32[137], stage0_32[138], stage0_32[139], stage0_32[140]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[51],stage1_34[52],stage1_33[105],stage1_32[178]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[141], stage0_32[142], stage0_32[143], stage0_32[144], stage0_32[145], stage0_32[146]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[52],stage1_34[53],stage1_33[106],stage1_32[179]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[147], stage0_32[148], stage0_32[149], stage0_32[150], stage0_32[151], stage0_32[152]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[53],stage1_34[54],stage1_33[107],stage1_32[180]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[153], stage0_32[154], stage0_32[155], stage0_32[156], stage0_32[157], stage0_32[158]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[54],stage1_34[55],stage1_33[108],stage1_32[181]}
   );
   gpc606_5 gpc1302 (
      {stage0_32[159], stage0_32[160], stage0_32[161], stage0_32[162], stage0_32[163], stage0_32[164]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[55],stage1_34[56],stage1_33[109],stage1_32[182]}
   );
   gpc606_5 gpc1303 (
      {stage0_32[165], stage0_32[166], stage0_32[167], stage0_32[168], stage0_32[169], stage0_32[170]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[56],stage1_34[57],stage1_33[110],stage1_32[183]}
   );
   gpc606_5 gpc1304 (
      {stage0_32[171], stage0_32[172], stage0_32[173], stage0_32[174], stage0_32[175], stage0_32[176]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[57],stage1_34[58],stage1_33[111],stage1_32[184]}
   );
   gpc606_5 gpc1305 (
      {stage0_32[177], stage0_32[178], stage0_32[179], stage0_32[180], stage0_32[181], stage0_32[182]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[58],stage1_34[59],stage1_33[112],stage1_32[185]}
   );
   gpc606_5 gpc1306 (
      {stage0_32[183], stage0_32[184], stage0_32[185], stage0_32[186], stage0_32[187], stage0_32[188]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[59],stage1_34[60],stage1_33[113],stage1_32[186]}
   );
   gpc606_5 gpc1307 (
      {stage0_32[189], stage0_32[190], stage0_32[191], stage0_32[192], stage0_32[193], stage0_32[194]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[60],stage1_34[61],stage1_33[114],stage1_32[187]}
   );
   gpc606_5 gpc1308 (
      {stage0_32[195], stage0_32[196], stage0_32[197], stage0_32[198], stage0_32[199], stage0_32[200]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[61],stage1_34[62],stage1_33[115],stage1_32[188]}
   );
   gpc606_5 gpc1309 (
      {stage0_32[201], stage0_32[202], stage0_32[203], stage0_32[204], stage0_32[205], stage0_32[206]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[62],stage1_34[63],stage1_33[116],stage1_32[189]}
   );
   gpc606_5 gpc1310 (
      {stage0_32[207], stage0_32[208], stage0_32[209], stage0_32[210], stage0_32[211], stage0_32[212]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[63],stage1_34[64],stage1_33[117],stage1_32[190]}
   );
   gpc606_5 gpc1311 (
      {stage0_32[213], stage0_32[214], stage0_32[215], stage0_32[216], stage0_32[217], stage0_32[218]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[64],stage1_34[65],stage1_33[118],stage1_32[191]}
   );
   gpc606_5 gpc1312 (
      {stage0_32[219], stage0_32[220], stage0_32[221], stage0_32[222], stage0_32[223], stage0_32[224]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[65],stage1_34[66],stage1_33[119],stage1_32[192]}
   );
   gpc606_5 gpc1313 (
      {stage0_32[225], stage0_32[226], stage0_32[227], stage0_32[228], stage0_32[229], stage0_32[230]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[66],stage1_34[67],stage1_33[120],stage1_32[193]}
   );
   gpc606_5 gpc1314 (
      {stage0_32[231], stage0_32[232], stage0_32[233], stage0_32[234], stage0_32[235], stage0_32[236]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[67],stage1_34[68],stage1_33[121],stage1_32[194]}
   );
   gpc606_5 gpc1315 (
      {stage0_32[237], stage0_32[238], stage0_32[239], stage0_32[240], stage0_32[241], stage0_32[242]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[68],stage1_34[69],stage1_33[122],stage1_32[195]}
   );
   gpc606_5 gpc1316 (
      {stage0_32[243], stage0_32[244], stage0_32[245], stage0_32[246], stage0_32[247], stage0_32[248]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[69],stage1_34[70],stage1_33[123],stage1_32[196]}
   );
   gpc606_5 gpc1317 (
      {stage0_32[249], stage0_32[250], stage0_32[251], stage0_32[252], stage0_32[253], stage0_32[254]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[70],stage1_34[71],stage1_33[124],stage1_32[197]}
   );
   gpc606_5 gpc1318 (
      {stage0_32[255], stage0_32[256], stage0_32[257], stage0_32[258], stage0_32[259], stage0_32[260]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[71],stage1_34[72],stage1_33[125],stage1_32[198]}
   );
   gpc606_5 gpc1319 (
      {stage0_32[261], stage0_32[262], stage0_32[263], stage0_32[264], stage0_32[265], stage0_32[266]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[72],stage1_34[73],stage1_33[126],stage1_32[199]}
   );
   gpc606_5 gpc1320 (
      {stage0_32[267], stage0_32[268], stage0_32[269], stage0_32[270], stage0_32[271], stage0_32[272]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[73],stage1_34[74],stage1_33[127],stage1_32[200]}
   );
   gpc606_5 gpc1321 (
      {stage0_32[273], stage0_32[274], stage0_32[275], stage0_32[276], stage0_32[277], stage0_32[278]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[74],stage1_34[75],stage1_33[128],stage1_32[201]}
   );
   gpc606_5 gpc1322 (
      {stage0_32[279], stage0_32[280], stage0_32[281], stage0_32[282], stage0_32[283], stage0_32[284]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[75],stage1_34[76],stage1_33[129],stage1_32[202]}
   );
   gpc606_5 gpc1323 (
      {stage0_32[285], stage0_32[286], stage0_32[287], stage0_32[288], stage0_32[289], stage0_32[290]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[76],stage1_34[77],stage1_33[130],stage1_32[203]}
   );
   gpc606_5 gpc1324 (
      {stage0_32[291], stage0_32[292], stage0_32[293], stage0_32[294], stage0_32[295], stage0_32[296]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[77],stage1_34[78],stage1_33[131],stage1_32[204]}
   );
   gpc606_5 gpc1325 (
      {stage0_32[297], stage0_32[298], stage0_32[299], stage0_32[300], stage0_32[301], stage0_32[302]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[78],stage1_34[79],stage1_33[132],stage1_32[205]}
   );
   gpc615_5 gpc1326 (
      {stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage0_34[264]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[44],stage1_35[79],stage1_34[80],stage1_33[133]}
   );
   gpc615_5 gpc1327 (
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220]},
      {stage0_34[265]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[45],stage1_35[80],stage1_34[81],stage1_33[134]}
   );
   gpc615_5 gpc1328 (
      {stage0_33[221], stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225]},
      {stage0_34[266]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[46],stage1_35[81],stage1_34[82],stage1_33[135]}
   );
   gpc615_5 gpc1329 (
      {stage0_33[226], stage0_33[227], stage0_33[228], stage0_33[229], stage0_33[230]},
      {stage0_34[267]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[47],stage1_35[82],stage1_34[83],stage1_33[136]}
   );
   gpc615_5 gpc1330 (
      {stage0_33[231], stage0_33[232], stage0_33[233], stage0_33[234], stage0_33[235]},
      {stage0_34[268]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[48],stage1_35[83],stage1_34[84],stage1_33[137]}
   );
   gpc615_5 gpc1331 (
      {stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239], stage0_33[240]},
      {stage0_34[269]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[49],stage1_35[84],stage1_34[85],stage1_33[138]}
   );
   gpc615_5 gpc1332 (
      {stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage0_34[270]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[50],stage1_35[85],stage1_34[86],stage1_33[139]}
   );
   gpc615_5 gpc1333 (
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250]},
      {stage0_34[271]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[51],stage1_35[86],stage1_34[87],stage1_33[140]}
   );
   gpc615_5 gpc1334 (
      {stage0_33[251], stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255]},
      {stage0_34[272]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[52],stage1_35[87],stage1_34[88],stage1_33[141]}
   );
   gpc615_5 gpc1335 (
      {stage0_33[256], stage0_33[257], stage0_33[258], stage0_33[259], stage0_33[260]},
      {stage0_34[273]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[53],stage1_35[88],stage1_34[89],stage1_33[142]}
   );
   gpc615_5 gpc1336 (
      {stage0_33[261], stage0_33[262], stage0_33[263], stage0_33[264], stage0_33[265]},
      {stage0_34[274]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[54],stage1_35[89],stage1_34[90],stage1_33[143]}
   );
   gpc615_5 gpc1337 (
      {stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269], stage0_33[270]},
      {stage0_34[275]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[55],stage1_35[90],stage1_34[91],stage1_33[144]}
   );
   gpc615_5 gpc1338 (
      {stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage0_34[276]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[56],stage1_35[91],stage1_34[92],stage1_33[145]}
   );
   gpc615_5 gpc1339 (
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280]},
      {stage0_34[277]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[57],stage1_35[92],stage1_34[93],stage1_33[146]}
   );
   gpc615_5 gpc1340 (
      {stage0_33[281], stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285]},
      {stage0_34[278]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[58],stage1_35[93],stage1_34[94],stage1_33[147]}
   );
   gpc615_5 gpc1341 (
      {stage0_33[286], stage0_33[287], stage0_33[288], stage0_33[289], stage0_33[290]},
      {stage0_34[279]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[59],stage1_35[94],stage1_34[95],stage1_33[148]}
   );
   gpc615_5 gpc1342 (
      {stage0_33[291], stage0_33[292], stage0_33[293], stage0_33[294], stage0_33[295]},
      {stage0_34[280]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[60],stage1_35[95],stage1_34[96],stage1_33[149]}
   );
   gpc615_5 gpc1343 (
      {stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299], stage0_33[300]},
      {stage0_34[281]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[61],stage1_35[96],stage1_34[97],stage1_33[150]}
   );
   gpc615_5 gpc1344 (
      {stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage0_34[282]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage1_37[18],stage1_36[62],stage1_35[97],stage1_34[98],stage1_33[151]}
   );
   gpc615_5 gpc1345 (
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310]},
      {stage0_34[283]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage1_37[19],stage1_36[63],stage1_35[98],stage1_34[99],stage1_33[152]}
   );
   gpc615_5 gpc1346 (
      {stage0_33[311], stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315]},
      {stage0_34[284]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage1_37[20],stage1_36[64],stage1_35[99],stage1_34[100],stage1_33[153]}
   );
   gpc615_5 gpc1347 (
      {stage0_33[316], stage0_33[317], stage0_33[318], stage0_33[319], stage0_33[320]},
      {stage0_34[285]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage1_37[21],stage1_36[65],stage1_35[100],stage1_34[101],stage1_33[154]}
   );
   gpc615_5 gpc1348 (
      {stage0_33[321], stage0_33[322], stage0_33[323], stage0_33[324], stage0_33[325]},
      {stage0_34[286]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage1_37[22],stage1_36[66],stage1_35[101],stage1_34[102],stage1_33[155]}
   );
   gpc615_5 gpc1349 (
      {stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329], stage0_33[330]},
      {stage0_34[287]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage1_37[23],stage1_36[67],stage1_35[102],stage1_34[103],stage1_33[156]}
   );
   gpc615_5 gpc1350 (
      {stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_34[288]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage1_37[24],stage1_36[68],stage1_35[103],stage1_34[104],stage1_33[157]}
   );
   gpc615_5 gpc1351 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340]},
      {stage0_34[289]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage1_37[25],stage1_36[69],stage1_35[104],stage1_34[105],stage1_33[158]}
   );
   gpc615_5 gpc1352 (
      {stage0_33[341], stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345]},
      {stage0_34[290]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage1_37[26],stage1_36[70],stage1_35[105],stage1_34[106],stage1_33[159]}
   );
   gpc615_5 gpc1353 (
      {stage0_33[346], stage0_33[347], stage0_33[348], stage0_33[349], stage0_33[350]},
      {stage0_34[291]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage1_37[27],stage1_36[71],stage1_35[106],stage1_34[107],stage1_33[160]}
   );
   gpc615_5 gpc1354 (
      {stage0_33[351], stage0_33[352], stage0_33[353], stage0_33[354], stage0_33[355]},
      {stage0_34[292]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage1_37[28],stage1_36[72],stage1_35[107],stage1_34[108],stage1_33[161]}
   );
   gpc615_5 gpc1355 (
      {stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359], stage0_33[360]},
      {stage0_34[293]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage1_37[29],stage1_36[73],stage1_35[108],stage1_34[109],stage1_33[162]}
   );
   gpc615_5 gpc1356 (
      {stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_34[294]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage1_37[30],stage1_36[74],stage1_35[109],stage1_34[110],stage1_33[163]}
   );
   gpc615_5 gpc1357 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370]},
      {stage0_34[295]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage1_37[31],stage1_36[75],stage1_35[110],stage1_34[111],stage1_33[164]}
   );
   gpc615_5 gpc1358 (
      {stage0_33[371], stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375]},
      {stage0_34[296]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage1_37[32],stage1_36[76],stage1_35[111],stage1_34[112],stage1_33[165]}
   );
   gpc615_5 gpc1359 (
      {stage0_33[376], stage0_33[377], stage0_33[378], stage0_33[379], stage0_33[380]},
      {stage0_34[297]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage1_37[33],stage1_36[77],stage1_35[112],stage1_34[113],stage1_33[166]}
   );
   gpc615_5 gpc1360 (
      {stage0_33[381], stage0_33[382], stage0_33[383], stage0_33[384], stage0_33[385]},
      {stage0_34[298]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage1_37[34],stage1_36[78],stage1_35[113],stage1_34[114],stage1_33[167]}
   );
   gpc615_5 gpc1361 (
      {stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389], stage0_33[390]},
      {stage0_34[299]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage1_37[35],stage1_36[79],stage1_35[114],stage1_34[115],stage1_33[168]}
   );
   gpc615_5 gpc1362 (
      {stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_34[300]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage1_37[36],stage1_36[80],stage1_35[115],stage1_34[116],stage1_33[169]}
   );
   gpc615_5 gpc1363 (
      {stage0_33[396], stage0_33[397], stage0_33[398], stage0_33[399], stage0_33[400]},
      {stage0_34[301]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage1_37[37],stage1_36[81],stage1_35[116],stage1_34[117],stage1_33[170]}
   );
   gpc615_5 gpc1364 (
      {stage0_33[401], stage0_33[402], stage0_33[403], stage0_33[404], stage0_33[405]},
      {stage0_34[302]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage1_37[38],stage1_36[82],stage1_35[117],stage1_34[118],stage1_33[171]}
   );
   gpc615_5 gpc1365 (
      {stage0_33[406], stage0_33[407], stage0_33[408], stage0_33[409], stage0_33[410]},
      {stage0_34[303]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage1_37[39],stage1_36[83],stage1_35[118],stage1_34[119],stage1_33[172]}
   );
   gpc615_5 gpc1366 (
      {stage0_33[411], stage0_33[412], stage0_33[413], stage0_33[414], stage0_33[415]},
      {stage0_34[304]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage1_37[40],stage1_36[84],stage1_35[119],stage1_34[120],stage1_33[173]}
   );
   gpc615_5 gpc1367 (
      {stage0_33[416], stage0_33[417], stage0_33[418], stage0_33[419], stage0_33[420]},
      {stage0_34[305]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage1_37[41],stage1_36[85],stage1_35[120],stage1_34[121],stage1_33[174]}
   );
   gpc615_5 gpc1368 (
      {stage0_33[421], stage0_33[422], stage0_33[423], stage0_33[424], stage0_33[425]},
      {stage0_34[306]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage1_37[42],stage1_36[86],stage1_35[121],stage1_34[122],stage1_33[175]}
   );
   gpc615_5 gpc1369 (
      {stage0_33[426], stage0_33[427], stage0_33[428], stage0_33[429], stage0_33[430]},
      {stage0_34[307]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage1_37[43],stage1_36[87],stage1_35[122],stage1_34[123],stage1_33[176]}
   );
   gpc615_5 gpc1370 (
      {stage0_33[431], stage0_33[432], stage0_33[433], stage0_33[434], stage0_33[435]},
      {stage0_34[308]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage1_37[44],stage1_36[88],stage1_35[123],stage1_34[124],stage1_33[177]}
   );
   gpc615_5 gpc1371 (
      {stage0_33[436], stage0_33[437], stage0_33[438], stage0_33[439], stage0_33[440]},
      {stage0_34[309]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage1_37[45],stage1_36[89],stage1_35[124],stage1_34[125],stage1_33[178]}
   );
   gpc615_5 gpc1372 (
      {stage0_33[441], stage0_33[442], stage0_33[443], stage0_33[444], stage0_33[445]},
      {stage0_34[310]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage1_37[46],stage1_36[90],stage1_35[125],stage1_34[126],stage1_33[179]}
   );
   gpc615_5 gpc1373 (
      {stage0_33[446], stage0_33[447], stage0_33[448], stage0_33[449], stage0_33[450]},
      {stage0_34[311]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage1_37[47],stage1_36[91],stage1_35[126],stage1_34[127],stage1_33[180]}
   );
   gpc615_5 gpc1374 (
      {stage0_33[451], stage0_33[452], stage0_33[453], stage0_33[454], stage0_33[455]},
      {stage0_34[312]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage1_37[48],stage1_36[92],stage1_35[127],stage1_34[128],stage1_33[181]}
   );
   gpc615_5 gpc1375 (
      {stage0_33[456], stage0_33[457], stage0_33[458], stage0_33[459], stage0_33[460]},
      {stage0_34[313]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage1_37[49],stage1_36[93],stage1_35[128],stage1_34[129],stage1_33[182]}
   );
   gpc615_5 gpc1376 (
      {stage0_33[461], stage0_33[462], stage0_33[463], stage0_33[464], stage0_33[465]},
      {stage0_34[314]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage1_37[50],stage1_36[94],stage1_35[129],stage1_34[130],stage1_33[183]}
   );
   gpc615_5 gpc1377 (
      {stage0_33[466], stage0_33[467], stage0_33[468], stage0_33[469], stage0_33[470]},
      {stage0_34[315]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage1_37[51],stage1_36[95],stage1_35[130],stage1_34[131],stage1_33[184]}
   );
   gpc615_5 gpc1378 (
      {stage0_33[471], stage0_33[472], stage0_33[473], stage0_33[474], stage0_33[475]},
      {stage0_34[316]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage1_37[52],stage1_36[96],stage1_35[131],stage1_34[132],stage1_33[185]}
   );
   gpc615_5 gpc1379 (
      {stage0_33[476], stage0_33[477], stage0_33[478], stage0_33[479], stage0_33[480]},
      {stage0_34[317]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage1_37[53],stage1_36[97],stage1_35[132],stage1_34[133],stage1_33[186]}
   );
   gpc615_5 gpc1380 (
      {stage0_33[481], stage0_33[482], stage0_33[483], stage0_33[484], stage0_33[485]},
      {stage0_34[318]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage1_37[54],stage1_36[98],stage1_35[133],stage1_34[134],stage1_33[187]}
   );
   gpc615_5 gpc1381 (
      {stage0_33[486], stage0_33[487], stage0_33[488], stage0_33[489], stage0_33[490]},
      {stage0_34[319]},
      {stage0_35[330], stage0_35[331], stage0_35[332], stage0_35[333], stage0_35[334], stage0_35[335]},
      {stage1_37[55],stage1_36[99],stage1_35[134],stage1_34[135],stage1_33[188]}
   );
   gpc1163_5 gpc1382 (
      {stage0_34[320], stage0_34[321], stage0_34[322]},
      {stage0_35[336], stage0_35[337], stage0_35[338], stage0_35[339], stage0_35[340], stage0_35[341]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[56],stage1_36[100],stage1_35[135],stage1_34[136]}
   );
   gpc1163_5 gpc1383 (
      {stage0_34[323], stage0_34[324], stage0_34[325]},
      {stage0_35[342], stage0_35[343], stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[57],stage1_36[101],stage1_35[136],stage1_34[137]}
   );
   gpc615_5 gpc1384 (
      {stage0_34[326], stage0_34[327], stage0_34[328], stage0_34[329], stage0_34[330]},
      {stage0_35[348]},
      {stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5], stage0_36[6], stage0_36[7]},
      {stage1_38[2],stage1_37[58],stage1_36[102],stage1_35[137],stage1_34[138]}
   );
   gpc615_5 gpc1385 (
      {stage0_34[331], stage0_34[332], stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[349]},
      {stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13]},
      {stage1_38[3],stage1_37[59],stage1_36[103],stage1_35[138],stage1_34[139]}
   );
   gpc615_5 gpc1386 (
      {stage0_34[336], stage0_34[337], stage0_34[338], stage0_34[339], stage0_34[340]},
      {stage0_35[350]},
      {stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19]},
      {stage1_38[4],stage1_37[60],stage1_36[104],stage1_35[139],stage1_34[140]}
   );
   gpc615_5 gpc1387 (
      {stage0_34[341], stage0_34[342], stage0_34[343], stage0_34[344], stage0_34[345]},
      {stage0_35[351]},
      {stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25]},
      {stage1_38[5],stage1_37[61],stage1_36[105],stage1_35[140],stage1_34[141]}
   );
   gpc615_5 gpc1388 (
      {stage0_34[346], stage0_34[347], stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[352]},
      {stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31]},
      {stage1_38[6],stage1_37[62],stage1_36[106],stage1_35[141],stage1_34[142]}
   );
   gpc615_5 gpc1389 (
      {stage0_34[351], stage0_34[352], stage0_34[353], stage0_34[354], stage0_34[355]},
      {stage0_35[353]},
      {stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37]},
      {stage1_38[7],stage1_37[63],stage1_36[107],stage1_35[142],stage1_34[143]}
   );
   gpc615_5 gpc1390 (
      {stage0_34[356], stage0_34[357], stage0_34[358], stage0_34[359], stage0_34[360]},
      {stage0_35[354]},
      {stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43]},
      {stage1_38[8],stage1_37[64],stage1_36[108],stage1_35[143],stage1_34[144]}
   );
   gpc615_5 gpc1391 (
      {stage0_34[361], stage0_34[362], stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[355]},
      {stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48], stage0_36[49]},
      {stage1_38[9],stage1_37[65],stage1_36[109],stage1_35[144],stage1_34[145]}
   );
   gpc615_5 gpc1392 (
      {stage0_34[366], stage0_34[367], stage0_34[368], stage0_34[369], stage0_34[370]},
      {stage0_35[356]},
      {stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54], stage0_36[55]},
      {stage1_38[10],stage1_37[66],stage1_36[110],stage1_35[145],stage1_34[146]}
   );
   gpc615_5 gpc1393 (
      {stage0_34[371], stage0_34[372], stage0_34[373], stage0_34[374], stage0_34[375]},
      {stage0_35[357]},
      {stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60], stage0_36[61]},
      {stage1_38[11],stage1_37[67],stage1_36[111],stage1_35[146],stage1_34[147]}
   );
   gpc615_5 gpc1394 (
      {stage0_34[376], stage0_34[377], stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[358]},
      {stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66], stage0_36[67]},
      {stage1_38[12],stage1_37[68],stage1_36[112],stage1_35[147],stage1_34[148]}
   );
   gpc615_5 gpc1395 (
      {stage0_34[381], stage0_34[382], stage0_34[383], stage0_34[384], stage0_34[385]},
      {stage0_35[359]},
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage1_38[13],stage1_37[69],stage1_36[113],stage1_35[148],stage1_34[149]}
   );
   gpc615_5 gpc1396 (
      {stage0_34[386], stage0_34[387], stage0_34[388], stage0_34[389], stage0_34[390]},
      {stage0_35[360]},
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage1_38[14],stage1_37[70],stage1_36[114],stage1_35[149],stage1_34[150]}
   );
   gpc615_5 gpc1397 (
      {stage0_34[391], stage0_34[392], stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[361]},
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage1_38[15],stage1_37[71],stage1_36[115],stage1_35[150],stage1_34[151]}
   );
   gpc606_5 gpc1398 (
      {stage0_35[362], stage0_35[363], stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367]},
      {stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5], stage0_37[6], stage0_37[7]},
      {stage1_39[0],stage1_38[16],stage1_37[72],stage1_36[116],stage1_35[151]}
   );
   gpc606_5 gpc1399 (
      {stage0_35[368], stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12], stage0_37[13]},
      {stage1_39[1],stage1_38[17],stage1_37[73],stage1_36[117],stage1_35[152]}
   );
   gpc606_5 gpc1400 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378], stage0_35[379]},
      {stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17], stage0_37[18], stage0_37[19]},
      {stage1_39[2],stage1_38[18],stage1_37[74],stage1_36[118],stage1_35[153]}
   );
   gpc606_5 gpc1401 (
      {stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383], stage0_35[384], stage0_35[385]},
      {stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23], stage0_37[24], stage0_37[25]},
      {stage1_39[3],stage1_38[19],stage1_37[75],stage1_36[119],stage1_35[154]}
   );
   gpc606_5 gpc1402 (
      {stage0_35[386], stage0_35[387], stage0_35[388], stage0_35[389], stage0_35[390], stage0_35[391]},
      {stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29], stage0_37[30], stage0_37[31]},
      {stage1_39[4],stage1_38[20],stage1_37[76],stage1_36[120],stage1_35[155]}
   );
   gpc606_5 gpc1403 (
      {stage0_35[392], stage0_35[393], stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397]},
      {stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35], stage0_37[36], stage0_37[37]},
      {stage1_39[5],stage1_38[21],stage1_37[77],stage1_36[121],stage1_35[156]}
   );
   gpc606_5 gpc1404 (
      {stage0_35[398], stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41], stage0_37[42], stage0_37[43]},
      {stage1_39[6],stage1_38[22],stage1_37[78],stage1_36[122],stage1_35[157]}
   );
   gpc606_5 gpc1405 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408], stage0_35[409]},
      {stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48], stage0_37[49]},
      {stage1_39[7],stage1_38[23],stage1_37[79],stage1_36[123],stage1_35[158]}
   );
   gpc606_5 gpc1406 (
      {stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413], stage0_35[414], stage0_35[415]},
      {stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54], stage0_37[55]},
      {stage1_39[8],stage1_38[24],stage1_37[80],stage1_36[124],stage1_35[159]}
   );
   gpc606_5 gpc1407 (
      {stage0_35[416], stage0_35[417], stage0_35[418], stage0_35[419], stage0_35[420], stage0_35[421]},
      {stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60], stage0_37[61]},
      {stage1_39[9],stage1_38[25],stage1_37[81],stage1_36[125],stage1_35[160]}
   );
   gpc606_5 gpc1408 (
      {stage0_35[422], stage0_35[423], stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427]},
      {stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66], stage0_37[67]},
      {stage1_39[10],stage1_38[26],stage1_37[82],stage1_36[126],stage1_35[161]}
   );
   gpc606_5 gpc1409 (
      {stage0_35[428], stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72], stage0_37[73]},
      {stage1_39[11],stage1_38[27],stage1_37[83],stage1_36[127],stage1_35[162]}
   );
   gpc606_5 gpc1410 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438], stage0_35[439]},
      {stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78], stage0_37[79]},
      {stage1_39[12],stage1_38[28],stage1_37[84],stage1_36[128],stage1_35[163]}
   );
   gpc606_5 gpc1411 (
      {stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443], stage0_35[444], stage0_35[445]},
      {stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84], stage0_37[85]},
      {stage1_39[13],stage1_38[29],stage1_37[85],stage1_36[129],stage1_35[164]}
   );
   gpc606_5 gpc1412 (
      {stage0_35[446], stage0_35[447], stage0_35[448], stage0_35[449], stage0_35[450], stage0_35[451]},
      {stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90], stage0_37[91]},
      {stage1_39[14],stage1_38[30],stage1_37[86],stage1_36[130],stage1_35[165]}
   );
   gpc606_5 gpc1413 (
      {stage0_35[452], stage0_35[453], stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457]},
      {stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96], stage0_37[97]},
      {stage1_39[15],stage1_38[31],stage1_37[87],stage1_36[131],stage1_35[166]}
   );
   gpc606_5 gpc1414 (
      {stage0_35[458], stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102], stage0_37[103]},
      {stage1_39[16],stage1_38[32],stage1_37[88],stage1_36[132],stage1_35[167]}
   );
   gpc606_5 gpc1415 (
      {stage0_35[464], stage0_35[465], stage0_35[466], stage0_35[467], stage0_35[468], stage0_35[469]},
      {stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108], stage0_37[109]},
      {stage1_39[17],stage1_38[33],stage1_37[89],stage1_36[133],stage1_35[168]}
   );
   gpc615_5 gpc1416 (
      {stage0_35[470], stage0_35[471], stage0_35[472], stage0_35[473], stage0_35[474]},
      {stage0_36[86]},
      {stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114], stage0_37[115]},
      {stage1_39[18],stage1_38[34],stage1_37[90],stage1_36[134],stage1_35[169]}
   );
   gpc615_5 gpc1417 (
      {stage0_35[475], stage0_35[476], stage0_35[477], stage0_35[478], stage0_35[479]},
      {stage0_36[87]},
      {stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120], stage0_37[121]},
      {stage1_39[19],stage1_38[35],stage1_37[91],stage1_36[135],stage1_35[170]}
   );
   gpc615_5 gpc1418 (
      {stage0_35[480], stage0_35[481], stage0_35[482], stage0_35[483], stage0_35[484]},
      {stage0_36[88]},
      {stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126], stage0_37[127]},
      {stage1_39[20],stage1_38[36],stage1_37[92],stage1_36[136],stage1_35[171]}
   );
   gpc615_5 gpc1419 (
      {stage0_35[485], stage0_35[486], stage0_35[487], stage0_35[488], stage0_35[489]},
      {stage0_36[89]},
      {stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132], stage0_37[133]},
      {stage1_39[21],stage1_38[37],stage1_37[93],stage1_36[137],stage1_35[172]}
   );
   gpc615_5 gpc1420 (
      {stage0_35[490], stage0_35[491], stage0_35[492], stage0_35[493], stage0_35[494]},
      {stage0_36[90]},
      {stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138], stage0_37[139]},
      {stage1_39[22],stage1_38[38],stage1_37[94],stage1_36[138],stage1_35[173]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[23],stage1_38[39],stage1_37[95],stage1_36[139]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[97], stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[24],stage1_38[40],stage1_37[96],stage1_36[140]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[25],stage1_38[41],stage1_37[97],stage1_36[141]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[109], stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[26],stage1_38[42],stage1_37[98],stage1_36[142]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[115], stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[27],stage1_38[43],stage1_37[99],stage1_36[143]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[121], stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[28],stage1_38[44],stage1_37[100],stage1_36[144]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[127], stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[29],stage1_38[45],stage1_37[101],stage1_36[145]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[133], stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[30],stage1_38[46],stage1_37[102],stage1_36[146]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[139], stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[31],stage1_38[47],stage1_37[103],stage1_36[147]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[145], stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[32],stage1_38[48],stage1_37[104],stage1_36[148]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[151], stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[33],stage1_38[49],stage1_37[105],stage1_36[149]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[157], stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[34],stage1_38[50],stage1_37[106],stage1_36[150]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[163], stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[35],stage1_38[51],stage1_37[107],stage1_36[151]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[169], stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[36],stage1_38[52],stage1_37[108],stage1_36[152]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[175], stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[37],stage1_38[53],stage1_37[109],stage1_36[153]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[181], stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[38],stage1_38[54],stage1_37[110],stage1_36[154]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[187], stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[39],stage1_38[55],stage1_37[111],stage1_36[155]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[193], stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[40],stage1_38[56],stage1_37[112],stage1_36[156]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[199], stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[41],stage1_38[57],stage1_37[113],stage1_36[157]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[205], stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[42],stage1_38[58],stage1_37[114],stage1_36[158]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[211], stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[43],stage1_38[59],stage1_37[115],stage1_36[159]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[217], stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[44],stage1_38[60],stage1_37[116],stage1_36[160]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[223], stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[45],stage1_38[61],stage1_37[117],stage1_36[161]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[229], stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[46],stage1_38[62],stage1_37[118],stage1_36[162]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[235], stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[47],stage1_38[63],stage1_37[119],stage1_36[163]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[241], stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[48],stage1_38[64],stage1_37[120],stage1_36[164]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[247], stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[49],stage1_38[65],stage1_37[121],stage1_36[165]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[253], stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[50],stage1_38[66],stage1_37[122],stage1_36[166]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[259], stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[51],stage1_38[67],stage1_37[123],stage1_36[167]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[265], stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[52],stage1_38[68],stage1_37[124],stage1_36[168]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[271], stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[53],stage1_38[69],stage1_37[125],stage1_36[169]}
   );
   gpc606_5 gpc1452 (
      {stage0_36[277], stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[54],stage1_38[70],stage1_37[126],stage1_36[170]}
   );
   gpc606_5 gpc1453 (
      {stage0_36[283], stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[55],stage1_38[71],stage1_37[127],stage1_36[171]}
   );
   gpc606_5 gpc1454 (
      {stage0_36[289], stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[56],stage1_38[72],stage1_37[128],stage1_36[172]}
   );
   gpc606_5 gpc1455 (
      {stage0_36[295], stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[57],stage1_38[73],stage1_37[129],stage1_36[173]}
   );
   gpc606_5 gpc1456 (
      {stage0_36[301], stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[58],stage1_38[74],stage1_37[130],stage1_36[174]}
   );
   gpc606_5 gpc1457 (
      {stage0_36[307], stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[59],stage1_38[75],stage1_37[131],stage1_36[175]}
   );
   gpc606_5 gpc1458 (
      {stage0_36[313], stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[60],stage1_38[76],stage1_37[132],stage1_36[176]}
   );
   gpc606_5 gpc1459 (
      {stage0_36[319], stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[61],stage1_38[77],stage1_37[133],stage1_36[177]}
   );
   gpc606_5 gpc1460 (
      {stage0_36[325], stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[62],stage1_38[78],stage1_37[134],stage1_36[178]}
   );
   gpc606_5 gpc1461 (
      {stage0_36[331], stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[63],stage1_38[79],stage1_37[135],stage1_36[179]}
   );
   gpc615_5 gpc1462 (
      {stage0_36[337], stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341]},
      {stage0_37[140]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[64],stage1_38[80],stage1_37[136],stage1_36[180]}
   );
   gpc615_5 gpc1463 (
      {stage0_36[342], stage0_36[343], stage0_36[344], stage0_36[345], stage0_36[346]},
      {stage0_37[141]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[65],stage1_38[81],stage1_37[137],stage1_36[181]}
   );
   gpc615_5 gpc1464 (
      {stage0_36[347], stage0_36[348], stage0_36[349], stage0_36[350], stage0_36[351]},
      {stage0_37[142]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[66],stage1_38[82],stage1_37[138],stage1_36[182]}
   );
   gpc615_5 gpc1465 (
      {stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355], stage0_36[356]},
      {stage0_37[143]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[67],stage1_38[83],stage1_37[139],stage1_36[183]}
   );
   gpc615_5 gpc1466 (
      {stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_37[144]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[68],stage1_38[84],stage1_37[140],stage1_36[184]}
   );
   gpc615_5 gpc1467 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366]},
      {stage0_37[145]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[69],stage1_38[85],stage1_37[141],stage1_36[185]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150], stage0_37[151]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[47],stage1_39[70],stage1_38[86],stage1_37[142]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156], stage0_37[157]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[48],stage1_39[71],stage1_38[87],stage1_37[143]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162], stage0_37[163]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[49],stage1_39[72],stage1_38[88],stage1_37[144]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168], stage0_37[169]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[50],stage1_39[73],stage1_38[89],stage1_37[145]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174], stage0_37[175]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[51],stage1_39[74],stage1_38[90],stage1_37[146]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180], stage0_37[181]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[52],stage1_39[75],stage1_38[91],stage1_37[147]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186], stage0_37[187]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[53],stage1_39[76],stage1_38[92],stage1_37[148]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192], stage0_37[193]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[54],stage1_39[77],stage1_38[93],stage1_37[149]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198], stage0_37[199]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[55],stage1_39[78],stage1_38[94],stage1_37[150]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204], stage0_37[205]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[56],stage1_39[79],stage1_38[95],stage1_37[151]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210], stage0_37[211]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[57],stage1_39[80],stage1_38[96],stage1_37[152]}
   );
   gpc606_5 gpc1479 (
      {stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216], stage0_37[217]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[58],stage1_39[81],stage1_38[97],stage1_37[153]}
   );
   gpc606_5 gpc1480 (
      {stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222], stage0_37[223]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[59],stage1_39[82],stage1_38[98],stage1_37[154]}
   );
   gpc606_5 gpc1481 (
      {stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228], stage0_37[229]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[60],stage1_39[83],stage1_38[99],stage1_37[155]}
   );
   gpc606_5 gpc1482 (
      {stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234], stage0_37[235]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[61],stage1_39[84],stage1_38[100],stage1_37[156]}
   );
   gpc606_5 gpc1483 (
      {stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240], stage0_37[241]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[62],stage1_39[85],stage1_38[101],stage1_37[157]}
   );
   gpc606_5 gpc1484 (
      {stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246], stage0_37[247]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[63],stage1_39[86],stage1_38[102],stage1_37[158]}
   );
   gpc606_5 gpc1485 (
      {stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252], stage0_37[253]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[64],stage1_39[87],stage1_38[103],stage1_37[159]}
   );
   gpc606_5 gpc1486 (
      {stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258], stage0_37[259]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[65],stage1_39[88],stage1_38[104],stage1_37[160]}
   );
   gpc606_5 gpc1487 (
      {stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264], stage0_37[265]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[66],stage1_39[89],stage1_38[105],stage1_37[161]}
   );
   gpc606_5 gpc1488 (
      {stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270], stage0_37[271]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[67],stage1_39[90],stage1_38[106],stage1_37[162]}
   );
   gpc606_5 gpc1489 (
      {stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276], stage0_37[277]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[68],stage1_39[91],stage1_38[107],stage1_37[163]}
   );
   gpc606_5 gpc1490 (
      {stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282], stage0_37[283]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[69],stage1_39[92],stage1_38[108],stage1_37[164]}
   );
   gpc606_5 gpc1491 (
      {stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288], stage0_37[289]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[70],stage1_39[93],stage1_38[109],stage1_37[165]}
   );
   gpc606_5 gpc1492 (
      {stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294], stage0_37[295]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[71],stage1_39[94],stage1_38[110],stage1_37[166]}
   );
   gpc606_5 gpc1493 (
      {stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300], stage0_37[301]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[72],stage1_39[95],stage1_38[111],stage1_37[167]}
   );
   gpc606_5 gpc1494 (
      {stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306], stage0_37[307]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[73],stage1_39[96],stage1_38[112],stage1_37[168]}
   );
   gpc606_5 gpc1495 (
      {stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312], stage0_37[313]},
      {stage0_39[162], stage0_39[163], stage0_39[164], stage0_39[165], stage0_39[166], stage0_39[167]},
      {stage1_41[27],stage1_40[74],stage1_39[97],stage1_38[113],stage1_37[169]}
   );
   gpc606_5 gpc1496 (
      {stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318], stage0_37[319]},
      {stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171], stage0_39[172], stage0_39[173]},
      {stage1_41[28],stage1_40[75],stage1_39[98],stage1_38[114],stage1_37[170]}
   );
   gpc606_5 gpc1497 (
      {stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324], stage0_37[325]},
      {stage0_39[174], stage0_39[175], stage0_39[176], stage0_39[177], stage0_39[178], stage0_39[179]},
      {stage1_41[29],stage1_40[76],stage1_39[99],stage1_38[115],stage1_37[171]}
   );
   gpc606_5 gpc1498 (
      {stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330], stage0_37[331]},
      {stage0_39[180], stage0_39[181], stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185]},
      {stage1_41[30],stage1_40[77],stage1_39[100],stage1_38[116],stage1_37[172]}
   );
   gpc606_5 gpc1499 (
      {stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336], stage0_37[337]},
      {stage0_39[186], stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage1_41[31],stage1_40[78],stage1_39[101],stage1_38[117],stage1_37[173]}
   );
   gpc606_5 gpc1500 (
      {stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342], stage0_37[343]},
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196], stage0_39[197]},
      {stage1_41[32],stage1_40[79],stage1_39[102],stage1_38[118],stage1_37[174]}
   );
   gpc606_5 gpc1501 (
      {stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348], stage0_37[349]},
      {stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201], stage0_39[202], stage0_39[203]},
      {stage1_41[33],stage1_40[80],stage1_39[103],stage1_38[119],stage1_37[175]}
   );
   gpc606_5 gpc1502 (
      {stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354], stage0_37[355]},
      {stage0_39[204], stage0_39[205], stage0_39[206], stage0_39[207], stage0_39[208], stage0_39[209]},
      {stage1_41[34],stage1_40[81],stage1_39[104],stage1_38[120],stage1_37[176]}
   );
   gpc606_5 gpc1503 (
      {stage0_37[356], stage0_37[357], stage0_37[358], stage0_37[359], stage0_37[360], stage0_37[361]},
      {stage0_39[210], stage0_39[211], stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215]},
      {stage1_41[35],stage1_40[82],stage1_39[105],stage1_38[121],stage1_37[177]}
   );
   gpc606_5 gpc1504 (
      {stage0_37[362], stage0_37[363], stage0_37[364], stage0_37[365], stage0_37[366], stage0_37[367]},
      {stage0_39[216], stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage1_41[36],stage1_40[83],stage1_39[106],stage1_38[122],stage1_37[178]}
   );
   gpc606_5 gpc1505 (
      {stage0_37[368], stage0_37[369], stage0_37[370], stage0_37[371], stage0_37[372], stage0_37[373]},
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226], stage0_39[227]},
      {stage1_41[37],stage1_40[84],stage1_39[107],stage1_38[123],stage1_37[179]}
   );
   gpc606_5 gpc1506 (
      {stage0_37[374], stage0_37[375], stage0_37[376], stage0_37[377], stage0_37[378], stage0_37[379]},
      {stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231], stage0_39[232], stage0_39[233]},
      {stage1_41[38],stage1_40[85],stage1_39[108],stage1_38[124],stage1_37[180]}
   );
   gpc606_5 gpc1507 (
      {stage0_37[380], stage0_37[381], stage0_37[382], stage0_37[383], stage0_37[384], stage0_37[385]},
      {stage0_39[234], stage0_39[235], stage0_39[236], stage0_39[237], stage0_39[238], stage0_39[239]},
      {stage1_41[39],stage1_40[86],stage1_39[109],stage1_38[125],stage1_37[181]}
   );
   gpc606_5 gpc1508 (
      {stage0_37[386], stage0_37[387], stage0_37[388], stage0_37[389], stage0_37[390], stage0_37[391]},
      {stage0_39[240], stage0_39[241], stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245]},
      {stage1_41[40],stage1_40[87],stage1_39[110],stage1_38[126],stage1_37[182]}
   );
   gpc615_5 gpc1509 (
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286]},
      {stage0_39[246]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[41],stage1_40[88],stage1_39[111],stage1_38[127]}
   );
   gpc615_5 gpc1510 (
      {stage0_38[287], stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291]},
      {stage0_39[247]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[42],stage1_40[89],stage1_39[112],stage1_38[128]}
   );
   gpc615_5 gpc1511 (
      {stage0_38[292], stage0_38[293], stage0_38[294], stage0_38[295], stage0_38[296]},
      {stage0_39[248]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[43],stage1_40[90],stage1_39[113],stage1_38[129]}
   );
   gpc615_5 gpc1512 (
      {stage0_38[297], stage0_38[298], stage0_38[299], stage0_38[300], stage0_38[301]},
      {stage0_39[249]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[44],stage1_40[91],stage1_39[114],stage1_38[130]}
   );
   gpc615_5 gpc1513 (
      {stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305], stage0_38[306]},
      {stage0_39[250]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[45],stage1_40[92],stage1_39[115],stage1_38[131]}
   );
   gpc615_5 gpc1514 (
      {stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage0_39[251]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[46],stage1_40[93],stage1_39[116],stage1_38[132]}
   );
   gpc615_5 gpc1515 (
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316]},
      {stage0_39[252]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[47],stage1_40[94],stage1_39[117],stage1_38[133]}
   );
   gpc615_5 gpc1516 (
      {stage0_38[317], stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321]},
      {stage0_39[253]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[48],stage1_40[95],stage1_39[118],stage1_38[134]}
   );
   gpc615_5 gpc1517 (
      {stage0_38[322], stage0_38[323], stage0_38[324], stage0_38[325], stage0_38[326]},
      {stage0_39[254]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[49],stage1_40[96],stage1_39[119],stage1_38[135]}
   );
   gpc615_5 gpc1518 (
      {stage0_38[327], stage0_38[328], stage0_38[329], stage0_38[330], stage0_38[331]},
      {stage0_39[255]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[50],stage1_40[97],stage1_39[120],stage1_38[136]}
   );
   gpc615_5 gpc1519 (
      {stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335], stage0_38[336]},
      {stage0_39[256]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[51],stage1_40[98],stage1_39[121],stage1_38[137]}
   );
   gpc615_5 gpc1520 (
      {stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage0_39[257]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[52],stage1_40[99],stage1_39[122],stage1_38[138]}
   );
   gpc615_5 gpc1521 (
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346]},
      {stage0_39[258]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[53],stage1_40[100],stage1_39[123],stage1_38[139]}
   );
   gpc615_5 gpc1522 (
      {stage0_38[347], stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351]},
      {stage0_39[259]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[54],stage1_40[101],stage1_39[124],stage1_38[140]}
   );
   gpc615_5 gpc1523 (
      {stage0_38[352], stage0_38[353], stage0_38[354], stage0_38[355], stage0_38[356]},
      {stage0_39[260]},
      {stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89]},
      {stage1_42[14],stage1_41[55],stage1_40[102],stage1_39[125],stage1_38[141]}
   );
   gpc615_5 gpc1524 (
      {stage0_38[357], stage0_38[358], stage0_38[359], stage0_38[360], stage0_38[361]},
      {stage0_39[261]},
      {stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95]},
      {stage1_42[15],stage1_41[56],stage1_40[103],stage1_39[126],stage1_38[142]}
   );
   gpc615_5 gpc1525 (
      {stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365], stage0_38[366]},
      {stage0_39[262]},
      {stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101]},
      {stage1_42[16],stage1_41[57],stage1_40[104],stage1_39[127],stage1_38[143]}
   );
   gpc615_5 gpc1526 (
      {stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370], stage0_38[371]},
      {stage0_39[263]},
      {stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107]},
      {stage1_42[17],stage1_41[58],stage1_40[105],stage1_39[128],stage1_38[144]}
   );
   gpc615_5 gpc1527 (
      {stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375], stage0_38[376]},
      {stage0_39[264]},
      {stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113]},
      {stage1_42[18],stage1_41[59],stage1_40[106],stage1_39[129],stage1_38[145]}
   );
   gpc615_5 gpc1528 (
      {stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380], stage0_38[381]},
      {stage0_39[265]},
      {stage0_40[114], stage0_40[115], stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119]},
      {stage1_42[19],stage1_41[60],stage1_40[107],stage1_39[130],stage1_38[146]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[266], stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270]},
      {stage0_40[120]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[20],stage1_41[61],stage1_40[108],stage1_39[131]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[271], stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275]},
      {stage0_40[121]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[21],stage1_41[62],stage1_40[109],stage1_39[132]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[276], stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280]},
      {stage0_40[122]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[22],stage1_41[63],stage1_40[110],stage1_39[133]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[281], stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285]},
      {stage0_40[123]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[23],stage1_41[64],stage1_40[111],stage1_39[134]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[286], stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290]},
      {stage0_40[124]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[24],stage1_41[65],stage1_40[112],stage1_39[135]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[291], stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295]},
      {stage0_40[125]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[25],stage1_41[66],stage1_40[113],stage1_39[136]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[296], stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300]},
      {stage0_40[126]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[26],stage1_41[67],stage1_40[114],stage1_39[137]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[301], stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305]},
      {stage0_40[127]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[27],stage1_41[68],stage1_40[115],stage1_39[138]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[306], stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310]},
      {stage0_40[128]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[28],stage1_41[69],stage1_40[116],stage1_39[139]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[311], stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315]},
      {stage0_40[129]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[29],stage1_41[70],stage1_40[117],stage1_39[140]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[316], stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320]},
      {stage0_40[130]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[30],stage1_41[71],stage1_40[118],stage1_39[141]}
   );
   gpc615_5 gpc1540 (
      {stage0_39[321], stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325]},
      {stage0_40[131]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[31],stage1_41[72],stage1_40[119],stage1_39[142]}
   );
   gpc615_5 gpc1541 (
      {stage0_39[326], stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330]},
      {stage0_40[132]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[32],stage1_41[73],stage1_40[120],stage1_39[143]}
   );
   gpc615_5 gpc1542 (
      {stage0_39[331], stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335]},
      {stage0_40[133]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[33],stage1_41[74],stage1_40[121],stage1_39[144]}
   );
   gpc615_5 gpc1543 (
      {stage0_39[336], stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340]},
      {stage0_40[134]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[34],stage1_41[75],stage1_40[122],stage1_39[145]}
   );
   gpc615_5 gpc1544 (
      {stage0_39[341], stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345]},
      {stage0_40[135]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[35],stage1_41[76],stage1_40[123],stage1_39[146]}
   );
   gpc615_5 gpc1545 (
      {stage0_39[346], stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350]},
      {stage0_40[136]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[36],stage1_41[77],stage1_40[124],stage1_39[147]}
   );
   gpc615_5 gpc1546 (
      {stage0_39[351], stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355]},
      {stage0_40[137]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[37],stage1_41[78],stage1_40[125],stage1_39[148]}
   );
   gpc615_5 gpc1547 (
      {stage0_39[356], stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360]},
      {stage0_40[138]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[38],stage1_41[79],stage1_40[126],stage1_39[149]}
   );
   gpc615_5 gpc1548 (
      {stage0_39[361], stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365]},
      {stage0_40[139]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[39],stage1_41[80],stage1_40[127],stage1_39[150]}
   );
   gpc615_5 gpc1549 (
      {stage0_39[366], stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370]},
      {stage0_40[140]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[40],stage1_41[81],stage1_40[128],stage1_39[151]}
   );
   gpc615_5 gpc1550 (
      {stage0_39[371], stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375]},
      {stage0_40[141]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[41],stage1_41[82],stage1_40[129],stage1_39[152]}
   );
   gpc615_5 gpc1551 (
      {stage0_39[376], stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380]},
      {stage0_40[142]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[42],stage1_41[83],stage1_40[130],stage1_39[153]}
   );
   gpc615_5 gpc1552 (
      {stage0_39[381], stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385]},
      {stage0_40[143]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[43],stage1_41[84],stage1_40[131],stage1_39[154]}
   );
   gpc615_5 gpc1553 (
      {stage0_39[386], stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390]},
      {stage0_40[144]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[44],stage1_41[85],stage1_40[132],stage1_39[155]}
   );
   gpc615_5 gpc1554 (
      {stage0_39[391], stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395]},
      {stage0_40[145]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[45],stage1_41[86],stage1_40[133],stage1_39[156]}
   );
   gpc615_5 gpc1555 (
      {stage0_39[396], stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400]},
      {stage0_40[146]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[46],stage1_41[87],stage1_40[134],stage1_39[157]}
   );
   gpc615_5 gpc1556 (
      {stage0_39[401], stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405]},
      {stage0_40[147]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[47],stage1_41[88],stage1_40[135],stage1_39[158]}
   );
   gpc615_5 gpc1557 (
      {stage0_39[406], stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410]},
      {stage0_40[148]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[48],stage1_41[89],stage1_40[136],stage1_39[159]}
   );
   gpc615_5 gpc1558 (
      {stage0_39[411], stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415]},
      {stage0_40[149]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[49],stage1_41[90],stage1_40[137],stage1_39[160]}
   );
   gpc615_5 gpc1559 (
      {stage0_39[416], stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420]},
      {stage0_40[150]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[50],stage1_41[91],stage1_40[138],stage1_39[161]}
   );
   gpc615_5 gpc1560 (
      {stage0_39[421], stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425]},
      {stage0_40[151]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[51],stage1_41[92],stage1_40[139],stage1_39[162]}
   );
   gpc615_5 gpc1561 (
      {stage0_39[426], stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430]},
      {stage0_40[152]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[52],stage1_41[93],stage1_40[140],stage1_39[163]}
   );
   gpc615_5 gpc1562 (
      {stage0_39[431], stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435]},
      {stage0_40[153]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[53],stage1_41[94],stage1_40[141],stage1_39[164]}
   );
   gpc615_5 gpc1563 (
      {stage0_39[436], stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440]},
      {stage0_40[154]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[54],stage1_41[95],stage1_40[142],stage1_39[165]}
   );
   gpc615_5 gpc1564 (
      {stage0_39[441], stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445]},
      {stage0_40[155]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[55],stage1_41[96],stage1_40[143],stage1_39[166]}
   );
   gpc615_5 gpc1565 (
      {stage0_39[446], stage0_39[447], stage0_39[448], stage0_39[449], stage0_39[450]},
      {stage0_40[156]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[56],stage1_41[97],stage1_40[144],stage1_39[167]}
   );
   gpc615_5 gpc1566 (
      {stage0_39[451], stage0_39[452], stage0_39[453], stage0_39[454], stage0_39[455]},
      {stage0_40[157]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[57],stage1_41[98],stage1_40[145],stage1_39[168]}
   );
   gpc615_5 gpc1567 (
      {stage0_39[456], stage0_39[457], stage0_39[458], stage0_39[459], stage0_39[460]},
      {stage0_40[158]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[58],stage1_41[99],stage1_40[146],stage1_39[169]}
   );
   gpc615_5 gpc1568 (
      {stage0_39[461], stage0_39[462], stage0_39[463], stage0_39[464], stage0_39[465]},
      {stage0_40[159]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[59],stage1_41[100],stage1_40[147],stage1_39[170]}
   );
   gpc615_5 gpc1569 (
      {stage0_39[466], stage0_39[467], stage0_39[468], stage0_39[469], stage0_39[470]},
      {stage0_40[160]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[60],stage1_41[101],stage1_40[148],stage1_39[171]}
   );
   gpc615_5 gpc1570 (
      {stage0_39[471], stage0_39[472], stage0_39[473], stage0_39[474], stage0_39[475]},
      {stage0_40[161]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[61],stage1_41[102],stage1_40[149],stage1_39[172]}
   );
   gpc615_5 gpc1571 (
      {stage0_39[476], stage0_39[477], stage0_39[478], stage0_39[479], stage0_39[480]},
      {stage0_40[162]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[62],stage1_41[103],stage1_40[150],stage1_39[173]}
   );
   gpc615_5 gpc1572 (
      {stage0_39[481], stage0_39[482], stage0_39[483], stage0_39[484], stage0_39[485]},
      {stage0_40[163]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[63],stage1_41[104],stage1_40[151],stage1_39[174]}
   );
   gpc615_5 gpc1573 (
      {stage0_39[486], stage0_39[487], stage0_39[488], stage0_39[489], stage0_39[490]},
      {stage0_40[164]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[64],stage1_41[105],stage1_40[152],stage1_39[175]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169], stage0_40[170]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[45],stage1_42[65],stage1_41[106],stage1_40[153]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175], stage0_40[176]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[46],stage1_42[66],stage1_41[107],stage1_40[154]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181], stage0_40[182]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[47],stage1_42[67],stage1_41[108],stage1_40[155]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187], stage0_40[188]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[48],stage1_42[68],stage1_41[109],stage1_40[156]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193], stage0_40[194]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[49],stage1_42[69],stage1_41[110],stage1_40[157]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199], stage0_40[200]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[50],stage1_42[70],stage1_41[111],stage1_40[158]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205], stage0_40[206]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[51],stage1_42[71],stage1_41[112],stage1_40[159]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211], stage0_40[212]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[52],stage1_42[72],stage1_41[113],stage1_40[160]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217], stage0_40[218]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[53],stage1_42[73],stage1_41[114],stage1_40[161]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223], stage0_40[224]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[54],stage1_42[74],stage1_41[115],stage1_40[162]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229], stage0_40[230]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[55],stage1_42[75],stage1_41[116],stage1_40[163]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235], stage0_40[236]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[56],stage1_42[76],stage1_41[117],stage1_40[164]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241], stage0_40[242]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[57],stage1_42[77],stage1_41[118],stage1_40[165]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247], stage0_40[248]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[58],stage1_42[78],stage1_41[119],stage1_40[166]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253], stage0_40[254]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[59],stage1_42[79],stage1_41[120],stage1_40[167]}
   );
   gpc606_5 gpc1589 (
      {stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259], stage0_40[260]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[60],stage1_42[80],stage1_41[121],stage1_40[168]}
   );
   gpc606_5 gpc1590 (
      {stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265], stage0_40[266]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[61],stage1_42[81],stage1_41[122],stage1_40[169]}
   );
   gpc606_5 gpc1591 (
      {stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271], stage0_40[272]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[62],stage1_42[82],stage1_41[123],stage1_40[170]}
   );
   gpc606_5 gpc1592 (
      {stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277], stage0_40[278]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[63],stage1_42[83],stage1_41[124],stage1_40[171]}
   );
   gpc606_5 gpc1593 (
      {stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283], stage0_40[284]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[64],stage1_42[84],stage1_41[125],stage1_40[172]}
   );
   gpc606_5 gpc1594 (
      {stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289], stage0_40[290]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[65],stage1_42[85],stage1_41[126],stage1_40[173]}
   );
   gpc606_5 gpc1595 (
      {stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295], stage0_40[296]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[66],stage1_42[86],stage1_41[127],stage1_40[174]}
   );
   gpc606_5 gpc1596 (
      {stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301], stage0_40[302]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[67],stage1_42[87],stage1_41[128],stage1_40[175]}
   );
   gpc606_5 gpc1597 (
      {stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307], stage0_40[308]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[68],stage1_42[88],stage1_41[129],stage1_40[176]}
   );
   gpc606_5 gpc1598 (
      {stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313], stage0_40[314]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[69],stage1_42[89],stage1_41[130],stage1_40[177]}
   );
   gpc606_5 gpc1599 (
      {stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319], stage0_40[320]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[70],stage1_42[90],stage1_41[131],stage1_40[178]}
   );
   gpc606_5 gpc1600 (
      {stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325], stage0_40[326]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[71],stage1_42[91],stage1_41[132],stage1_40[179]}
   );
   gpc606_5 gpc1601 (
      {stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331], stage0_40[332]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[72],stage1_42[92],stage1_41[133],stage1_40[180]}
   );
   gpc606_5 gpc1602 (
      {stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337], stage0_40[338]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[73],stage1_42[93],stage1_41[134],stage1_40[181]}
   );
   gpc606_5 gpc1603 (
      {stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343], stage0_40[344]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[74],stage1_42[94],stage1_41[135],stage1_40[182]}
   );
   gpc606_5 gpc1604 (
      {stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349], stage0_40[350]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[75],stage1_42[95],stage1_41[136],stage1_40[183]}
   );
   gpc606_5 gpc1605 (
      {stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355], stage0_40[356]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[76],stage1_42[96],stage1_41[137],stage1_40[184]}
   );
   gpc606_5 gpc1606 (
      {stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361], stage0_40[362]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[77],stage1_42[97],stage1_41[138],stage1_40[185]}
   );
   gpc606_5 gpc1607 (
      {stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367], stage0_40[368]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[78],stage1_42[98],stage1_41[139],stage1_40[186]}
   );
   gpc606_5 gpc1608 (
      {stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373], stage0_40[374]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[79],stage1_42[99],stage1_41[140],stage1_40[187]}
   );
   gpc606_5 gpc1609 (
      {stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379], stage0_40[380]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[80],stage1_42[100],stage1_41[141],stage1_40[188]}
   );
   gpc606_5 gpc1610 (
      {stage0_40[381], stage0_40[382], stage0_40[383], stage0_40[384], stage0_40[385], stage0_40[386]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[81],stage1_42[101],stage1_41[142],stage1_40[189]}
   );
   gpc606_5 gpc1611 (
      {stage0_40[387], stage0_40[388], stage0_40[389], stage0_40[390], stage0_40[391], stage0_40[392]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[82],stage1_42[102],stage1_41[143],stage1_40[190]}
   );
   gpc606_5 gpc1612 (
      {stage0_40[393], stage0_40[394], stage0_40[395], stage0_40[396], stage0_40[397], stage0_40[398]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[83],stage1_42[103],stage1_41[144],stage1_40[191]}
   );
   gpc606_5 gpc1613 (
      {stage0_40[399], stage0_40[400], stage0_40[401], stage0_40[402], stage0_40[403], stage0_40[404]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[84],stage1_42[104],stage1_41[145],stage1_40[192]}
   );
   gpc606_5 gpc1614 (
      {stage0_40[405], stage0_40[406], stage0_40[407], stage0_40[408], stage0_40[409], stage0_40[410]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[85],stage1_42[105],stage1_41[146],stage1_40[193]}
   );
   gpc606_5 gpc1615 (
      {stage0_40[411], stage0_40[412], stage0_40[413], stage0_40[414], stage0_40[415], stage0_40[416]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[86],stage1_42[106],stage1_41[147],stage1_40[194]}
   );
   gpc606_5 gpc1616 (
      {stage0_40[417], stage0_40[418], stage0_40[419], stage0_40[420], stage0_40[421], stage0_40[422]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[87],stage1_42[107],stage1_41[148],stage1_40[195]}
   );
   gpc606_5 gpc1617 (
      {stage0_40[423], stage0_40[424], stage0_40[425], stage0_40[426], stage0_40[427], stage0_40[428]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[88],stage1_42[108],stage1_41[149],stage1_40[196]}
   );
   gpc606_5 gpc1618 (
      {stage0_40[429], stage0_40[430], stage0_40[431], stage0_40[432], stage0_40[433], stage0_40[434]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[89],stage1_42[109],stage1_41[150],stage1_40[197]}
   );
   gpc606_5 gpc1619 (
      {stage0_40[435], stage0_40[436], stage0_40[437], stage0_40[438], stage0_40[439], stage0_40[440]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[90],stage1_42[110],stage1_41[151],stage1_40[198]}
   );
   gpc606_5 gpc1620 (
      {stage0_40[441], stage0_40[442], stage0_40[443], stage0_40[444], stage0_40[445], stage0_40[446]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[91],stage1_42[111],stage1_41[152],stage1_40[199]}
   );
   gpc606_5 gpc1621 (
      {stage0_40[447], stage0_40[448], stage0_40[449], stage0_40[450], stage0_40[451], stage0_40[452]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[92],stage1_42[112],stage1_41[153],stage1_40[200]}
   );
   gpc606_5 gpc1622 (
      {stage0_40[453], stage0_40[454], stage0_40[455], stage0_40[456], stage0_40[457], stage0_40[458]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[93],stage1_42[113],stage1_41[154],stage1_40[201]}
   );
   gpc606_5 gpc1623 (
      {stage0_40[459], stage0_40[460], stage0_40[461], stage0_40[462], stage0_40[463], stage0_40[464]},
      {stage0_42[294], stage0_42[295], stage0_42[296], stage0_42[297], stage0_42[298], stage0_42[299]},
      {stage1_44[49],stage1_43[94],stage1_42[114],stage1_41[155],stage1_40[202]}
   );
   gpc606_5 gpc1624 (
      {stage0_40[465], stage0_40[466], stage0_40[467], stage0_40[468], stage0_40[469], stage0_40[470]},
      {stage0_42[300], stage0_42[301], stage0_42[302], stage0_42[303], stage0_42[304], stage0_42[305]},
      {stage1_44[50],stage1_43[95],stage1_42[115],stage1_41[156],stage1_40[203]}
   );
   gpc606_5 gpc1625 (
      {stage0_40[471], stage0_40[472], stage0_40[473], stage0_40[474], stage0_40[475], stage0_40[476]},
      {stage0_42[306], stage0_42[307], stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311]},
      {stage1_44[51],stage1_43[96],stage1_42[116],stage1_41[157],stage1_40[204]}
   );
   gpc606_5 gpc1626 (
      {stage0_40[477], stage0_40[478], stage0_40[479], stage0_40[480], stage0_40[481], stage0_40[482]},
      {stage0_42[312], stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage1_44[52],stage1_43[97],stage1_42[117],stage1_41[158],stage1_40[205]}
   );
   gpc606_5 gpc1627 (
      {stage0_40[483], stage0_40[484], stage0_40[485], stage0_40[486], stage0_40[487], stage0_40[488]},
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322], stage0_42[323]},
      {stage1_44[53],stage1_43[98],stage1_42[118],stage1_41[159],stage1_40[206]}
   );
   gpc606_5 gpc1628 (
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[54],stage1_43[99],stage1_42[119],stage1_41[160]}
   );
   gpc606_5 gpc1629 (
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[55],stage1_43[100],stage1_42[120],stage1_41[161]}
   );
   gpc606_5 gpc1630 (
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[56],stage1_43[101],stage1_42[121],stage1_41[162]}
   );
   gpc606_5 gpc1631 (
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[57],stage1_43[102],stage1_42[122],stage1_41[163]}
   );
   gpc606_5 gpc1632 (
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[58],stage1_43[103],stage1_42[123],stage1_41[164]}
   );
   gpc606_5 gpc1633 (
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[59],stage1_43[104],stage1_42[124],stage1_41[165]}
   );
   gpc606_5 gpc1634 (
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[60],stage1_43[105],stage1_42[125],stage1_41[166]}
   );
   gpc606_5 gpc1635 (
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[61],stage1_43[106],stage1_42[126],stage1_41[167]}
   );
   gpc606_5 gpc1636 (
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[62],stage1_43[107],stage1_42[127],stage1_41[168]}
   );
   gpc606_5 gpc1637 (
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[63],stage1_43[108],stage1_42[128],stage1_41[169]}
   );
   gpc606_5 gpc1638 (
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[64],stage1_43[109],stage1_42[129],stage1_41[170]}
   );
   gpc606_5 gpc1639 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[65],stage1_43[110],stage1_42[130],stage1_41[171]}
   );
   gpc606_5 gpc1640 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[66],stage1_43[111],stage1_42[131],stage1_41[172]}
   );
   gpc606_5 gpc1641 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[67],stage1_43[112],stage1_42[132],stage1_41[173]}
   );
   gpc606_5 gpc1642 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[68],stage1_43[113],stage1_42[133],stage1_41[174]}
   );
   gpc606_5 gpc1643 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[69],stage1_43[114],stage1_42[134],stage1_41[175]}
   );
   gpc606_5 gpc1644 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[70],stage1_43[115],stage1_42[135],stage1_41[176]}
   );
   gpc606_5 gpc1645 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[71],stage1_43[116],stage1_42[136],stage1_41[177]}
   );
   gpc606_5 gpc1646 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[72],stage1_43[117],stage1_42[137],stage1_41[178]}
   );
   gpc606_5 gpc1647 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[73],stage1_43[118],stage1_42[138],stage1_41[179]}
   );
   gpc606_5 gpc1648 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[74],stage1_43[119],stage1_42[139],stage1_41[180]}
   );
   gpc606_5 gpc1649 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[75],stage1_43[120],stage1_42[140],stage1_41[181]}
   );
   gpc606_5 gpc1650 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[76],stage1_43[121],stage1_42[141],stage1_41[182]}
   );
   gpc606_5 gpc1651 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[77],stage1_43[122],stage1_42[142],stage1_41[183]}
   );
   gpc606_5 gpc1652 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[78],stage1_43[123],stage1_42[143],stage1_41[184]}
   );
   gpc606_5 gpc1653 (
      {stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327], stage0_42[328], stage0_42[329]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[79],stage1_43[124],stage1_42[144]}
   );
   gpc606_5 gpc1654 (
      {stage0_42[330], stage0_42[331], stage0_42[332], stage0_42[333], stage0_42[334], stage0_42[335]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[80],stage1_43[125],stage1_42[145]}
   );
   gpc606_5 gpc1655 (
      {stage0_42[336], stage0_42[337], stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[81],stage1_43[126],stage1_42[146]}
   );
   gpc606_5 gpc1656 (
      {stage0_42[342], stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[82],stage1_43[127],stage1_42[147]}
   );
   gpc606_5 gpc1657 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352], stage0_42[353]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[83],stage1_43[128],stage1_42[148]}
   );
   gpc606_5 gpc1658 (
      {stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357], stage0_42[358], stage0_42[359]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[84],stage1_43[129],stage1_42[149]}
   );
   gpc606_5 gpc1659 (
      {stage0_42[360], stage0_42[361], stage0_42[362], stage0_42[363], stage0_42[364], stage0_42[365]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[85],stage1_43[130],stage1_42[150]}
   );
   gpc615_5 gpc1660 (
      {stage0_42[366], stage0_42[367], stage0_42[368], stage0_42[369], stage0_42[370]},
      {stage0_43[150]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[86],stage1_43[131],stage1_42[151]}
   );
   gpc615_5 gpc1661 (
      {stage0_42[371], stage0_42[372], stage0_42[373], stage0_42[374], stage0_42[375]},
      {stage0_43[151]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[87],stage1_43[132],stage1_42[152]}
   );
   gpc615_5 gpc1662 (
      {stage0_42[376], stage0_42[377], stage0_42[378], stage0_42[379], stage0_42[380]},
      {stage0_43[152]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[88],stage1_43[133],stage1_42[153]}
   );
   gpc615_5 gpc1663 (
      {stage0_42[381], stage0_42[382], stage0_42[383], stage0_42[384], stage0_42[385]},
      {stage0_43[153]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[89],stage1_43[134],stage1_42[154]}
   );
   gpc615_5 gpc1664 (
      {stage0_42[386], stage0_42[387], stage0_42[388], stage0_42[389], stage0_42[390]},
      {stage0_43[154]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[90],stage1_43[135],stage1_42[155]}
   );
   gpc615_5 gpc1665 (
      {stage0_42[391], stage0_42[392], stage0_42[393], stage0_42[394], stage0_42[395]},
      {stage0_43[155]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[91],stage1_43[136],stage1_42[156]}
   );
   gpc615_5 gpc1666 (
      {stage0_42[396], stage0_42[397], stage0_42[398], stage0_42[399], stage0_42[400]},
      {stage0_43[156]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[92],stage1_43[137],stage1_42[157]}
   );
   gpc615_5 gpc1667 (
      {stage0_42[401], stage0_42[402], stage0_42[403], stage0_42[404], stage0_42[405]},
      {stage0_43[157]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[93],stage1_43[138],stage1_42[158]}
   );
   gpc615_5 gpc1668 (
      {stage0_42[406], stage0_42[407], stage0_42[408], stage0_42[409], stage0_42[410]},
      {stage0_43[158]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[94],stage1_43[139],stage1_42[159]}
   );
   gpc615_5 gpc1669 (
      {stage0_42[411], stage0_42[412], stage0_42[413], stage0_42[414], stage0_42[415]},
      {stage0_43[159]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[95],stage1_43[140],stage1_42[160]}
   );
   gpc615_5 gpc1670 (
      {stage0_42[416], stage0_42[417], stage0_42[418], stage0_42[419], stage0_42[420]},
      {stage0_43[160]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[96],stage1_43[141],stage1_42[161]}
   );
   gpc615_5 gpc1671 (
      {stage0_42[421], stage0_42[422], stage0_42[423], stage0_42[424], stage0_42[425]},
      {stage0_43[161]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[97],stage1_43[142],stage1_42[162]}
   );
   gpc615_5 gpc1672 (
      {stage0_42[426], stage0_42[427], stage0_42[428], stage0_42[429], stage0_42[430]},
      {stage0_43[162]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[98],stage1_43[143],stage1_42[163]}
   );
   gpc615_5 gpc1673 (
      {stage0_42[431], stage0_42[432], stage0_42[433], stage0_42[434], stage0_42[435]},
      {stage0_43[163]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[99],stage1_43[144],stage1_42[164]}
   );
   gpc615_5 gpc1674 (
      {stage0_42[436], stage0_42[437], stage0_42[438], stage0_42[439], stage0_42[440]},
      {stage0_43[164]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[100],stage1_43[145],stage1_42[165]}
   );
   gpc615_5 gpc1675 (
      {stage0_42[441], stage0_42[442], stage0_42[443], stage0_42[444], stage0_42[445]},
      {stage0_43[165]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[101],stage1_43[146],stage1_42[166]}
   );
   gpc615_5 gpc1676 (
      {stage0_42[446], stage0_42[447], stage0_42[448], stage0_42[449], stage0_42[450]},
      {stage0_43[166]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[102],stage1_43[147],stage1_42[167]}
   );
   gpc606_5 gpc1677 (
      {stage0_43[167], stage0_43[168], stage0_43[169], stage0_43[170], stage0_43[171], stage0_43[172]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[24],stage1_45[49],stage1_44[103],stage1_43[148]}
   );
   gpc606_5 gpc1678 (
      {stage0_43[173], stage0_43[174], stage0_43[175], stage0_43[176], stage0_43[177], stage0_43[178]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[25],stage1_45[50],stage1_44[104],stage1_43[149]}
   );
   gpc606_5 gpc1679 (
      {stage0_43[179], stage0_43[180], stage0_43[181], stage0_43[182], stage0_43[183], stage0_43[184]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[26],stage1_45[51],stage1_44[105],stage1_43[150]}
   );
   gpc606_5 gpc1680 (
      {stage0_43[185], stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[27],stage1_45[52],stage1_44[106],stage1_43[151]}
   );
   gpc606_5 gpc1681 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195], stage0_43[196]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[28],stage1_45[53],stage1_44[107],stage1_43[152]}
   );
   gpc606_5 gpc1682 (
      {stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200], stage0_43[201], stage0_43[202]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[29],stage1_45[54],stage1_44[108],stage1_43[153]}
   );
   gpc606_5 gpc1683 (
      {stage0_43[203], stage0_43[204], stage0_43[205], stage0_43[206], stage0_43[207], stage0_43[208]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[30],stage1_45[55],stage1_44[109],stage1_43[154]}
   );
   gpc606_5 gpc1684 (
      {stage0_43[209], stage0_43[210], stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[31],stage1_45[56],stage1_44[110],stage1_43[155]}
   );
   gpc606_5 gpc1685 (
      {stage0_43[215], stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[32],stage1_45[57],stage1_44[111],stage1_43[156]}
   );
   gpc606_5 gpc1686 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225], stage0_43[226]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[33],stage1_45[58],stage1_44[112],stage1_43[157]}
   );
   gpc606_5 gpc1687 (
      {stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230], stage0_43[231], stage0_43[232]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[34],stage1_45[59],stage1_44[113],stage1_43[158]}
   );
   gpc606_5 gpc1688 (
      {stage0_43[233], stage0_43[234], stage0_43[235], stage0_43[236], stage0_43[237], stage0_43[238]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[35],stage1_45[60],stage1_44[114],stage1_43[159]}
   );
   gpc606_5 gpc1689 (
      {stage0_43[239], stage0_43[240], stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[36],stage1_45[61],stage1_44[115],stage1_43[160]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[245], stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249]},
      {stage0_44[144]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[37],stage1_45[62],stage1_44[116],stage1_43[161]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[250], stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254]},
      {stage0_44[145]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[38],stage1_45[63],stage1_44[117],stage1_43[162]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[255], stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259]},
      {stage0_44[146]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[39],stage1_45[64],stage1_44[118],stage1_43[163]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[260], stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264]},
      {stage0_44[147]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[40],stage1_45[65],stage1_44[119],stage1_43[164]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[265], stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269]},
      {stage0_44[148]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[41],stage1_45[66],stage1_44[120],stage1_43[165]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[270], stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274]},
      {stage0_44[149]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[42],stage1_45[67],stage1_44[121],stage1_43[166]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[275], stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279]},
      {stage0_44[150]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[43],stage1_45[68],stage1_44[122],stage1_43[167]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[280], stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284]},
      {stage0_44[151]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[44],stage1_45[69],stage1_44[123],stage1_43[168]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[285], stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289]},
      {stage0_44[152]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[45],stage1_45[70],stage1_44[124],stage1_43[169]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[290], stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294]},
      {stage0_44[153]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[46],stage1_45[71],stage1_44[125],stage1_43[170]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[295], stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299]},
      {stage0_44[154]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[47],stage1_45[72],stage1_44[126],stage1_43[171]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[300], stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304]},
      {stage0_44[155]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[48],stage1_45[73],stage1_44[127],stage1_43[172]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[305], stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309]},
      {stage0_44[156]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[49],stage1_45[74],stage1_44[128],stage1_43[173]}
   );
   gpc615_5 gpc1703 (
      {stage0_43[310], stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314]},
      {stage0_44[157]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[50],stage1_45[75],stage1_44[129],stage1_43[174]}
   );
   gpc615_5 gpc1704 (
      {stage0_43[315], stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319]},
      {stage0_44[158]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[51],stage1_45[76],stage1_44[130],stage1_43[175]}
   );
   gpc615_5 gpc1705 (
      {stage0_43[320], stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324]},
      {stage0_44[159]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[52],stage1_45[77],stage1_44[131],stage1_43[176]}
   );
   gpc615_5 gpc1706 (
      {stage0_43[325], stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329]},
      {stage0_44[160]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[53],stage1_45[78],stage1_44[132],stage1_43[177]}
   );
   gpc615_5 gpc1707 (
      {stage0_43[330], stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334]},
      {stage0_44[161]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[54],stage1_45[79],stage1_44[133],stage1_43[178]}
   );
   gpc615_5 gpc1708 (
      {stage0_43[335], stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339]},
      {stage0_44[162]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[55],stage1_45[80],stage1_44[134],stage1_43[179]}
   );
   gpc615_5 gpc1709 (
      {stage0_43[340], stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344]},
      {stage0_44[163]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[56],stage1_45[81],stage1_44[135],stage1_43[180]}
   );
   gpc615_5 gpc1710 (
      {stage0_43[345], stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349]},
      {stage0_44[164]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[57],stage1_45[82],stage1_44[136],stage1_43[181]}
   );
   gpc615_5 gpc1711 (
      {stage0_43[350], stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354]},
      {stage0_44[165]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[58],stage1_45[83],stage1_44[137],stage1_43[182]}
   );
   gpc615_5 gpc1712 (
      {stage0_43[355], stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359]},
      {stage0_44[166]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[59],stage1_45[84],stage1_44[138],stage1_43[183]}
   );
   gpc615_5 gpc1713 (
      {stage0_43[360], stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364]},
      {stage0_44[167]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[60],stage1_45[85],stage1_44[139],stage1_43[184]}
   );
   gpc615_5 gpc1714 (
      {stage0_43[365], stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369]},
      {stage0_44[168]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[61],stage1_45[86],stage1_44[140],stage1_43[185]}
   );
   gpc615_5 gpc1715 (
      {stage0_43[370], stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374]},
      {stage0_44[169]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[62],stage1_45[87],stage1_44[141],stage1_43[186]}
   );
   gpc615_5 gpc1716 (
      {stage0_43[375], stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379]},
      {stage0_44[170]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[63],stage1_45[88],stage1_44[142],stage1_43[187]}
   );
   gpc615_5 gpc1717 (
      {stage0_43[380], stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384]},
      {stage0_44[171]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[64],stage1_45[89],stage1_44[143],stage1_43[188]}
   );
   gpc615_5 gpc1718 (
      {stage0_43[385], stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389]},
      {stage0_44[172]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[65],stage1_45[90],stage1_44[144],stage1_43[189]}
   );
   gpc615_5 gpc1719 (
      {stage0_43[390], stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394]},
      {stage0_44[173]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[66],stage1_45[91],stage1_44[145],stage1_43[190]}
   );
   gpc615_5 gpc1720 (
      {stage0_43[395], stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399]},
      {stage0_44[174]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[67],stage1_45[92],stage1_44[146],stage1_43[191]}
   );
   gpc615_5 gpc1721 (
      {stage0_43[400], stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404]},
      {stage0_44[175]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[68],stage1_45[93],stage1_44[147],stage1_43[192]}
   );
   gpc615_5 gpc1722 (
      {stage0_43[405], stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409]},
      {stage0_44[176]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[69],stage1_45[94],stage1_44[148],stage1_43[193]}
   );
   gpc615_5 gpc1723 (
      {stage0_43[410], stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414]},
      {stage0_44[177]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[70],stage1_45[95],stage1_44[149],stage1_43[194]}
   );
   gpc615_5 gpc1724 (
      {stage0_43[415], stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419]},
      {stage0_44[178]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[71],stage1_45[96],stage1_44[150],stage1_43[195]}
   );
   gpc615_5 gpc1725 (
      {stage0_43[420], stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424]},
      {stage0_44[179]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[72],stage1_45[97],stage1_44[151],stage1_43[196]}
   );
   gpc615_5 gpc1726 (
      {stage0_43[425], stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429]},
      {stage0_44[180]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[73],stage1_45[98],stage1_44[152],stage1_43[197]}
   );
   gpc615_5 gpc1727 (
      {stage0_43[430], stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434]},
      {stage0_44[181]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[74],stage1_45[99],stage1_44[153],stage1_43[198]}
   );
   gpc615_5 gpc1728 (
      {stage0_43[435], stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439]},
      {stage0_44[182]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[75],stage1_45[100],stage1_44[154],stage1_43[199]}
   );
   gpc615_5 gpc1729 (
      {stage0_43[440], stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444]},
      {stage0_44[183]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[76],stage1_45[101],stage1_44[155],stage1_43[200]}
   );
   gpc615_5 gpc1730 (
      {stage0_43[445], stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449]},
      {stage0_44[184]},
      {stage0_45[318], stage0_45[319], stage0_45[320], stage0_45[321], stage0_45[322], stage0_45[323]},
      {stage1_47[53],stage1_46[77],stage1_45[102],stage1_44[156],stage1_43[201]}
   );
   gpc615_5 gpc1731 (
      {stage0_43[450], stage0_43[451], stage0_43[452], stage0_43[453], stage0_43[454]},
      {stage0_44[185]},
      {stage0_45[324], stage0_45[325], stage0_45[326], stage0_45[327], stage0_45[328], stage0_45[329]},
      {stage1_47[54],stage1_46[78],stage1_45[103],stage1_44[157],stage1_43[202]}
   );
   gpc615_5 gpc1732 (
      {stage0_43[455], stage0_43[456], stage0_43[457], stage0_43[458], stage0_43[459]},
      {stage0_44[186]},
      {stage0_45[330], stage0_45[331], stage0_45[332], stage0_45[333], stage0_45[334], stage0_45[335]},
      {stage1_47[55],stage1_46[79],stage1_45[104],stage1_44[158],stage1_43[203]}
   );
   gpc615_5 gpc1733 (
      {stage0_43[460], stage0_43[461], stage0_43[462], stage0_43[463], stage0_43[464]},
      {stage0_44[187]},
      {stage0_45[336], stage0_45[337], stage0_45[338], stage0_45[339], stage0_45[340], stage0_45[341]},
      {stage1_47[56],stage1_46[80],stage1_45[105],stage1_44[159],stage1_43[204]}
   );
   gpc615_5 gpc1734 (
      {stage0_43[465], stage0_43[466], stage0_43[467], stage0_43[468], stage0_43[469]},
      {stage0_44[188]},
      {stage0_45[342], stage0_45[343], stage0_45[344], stage0_45[345], stage0_45[346], stage0_45[347]},
      {stage1_47[57],stage1_46[81],stage1_45[106],stage1_44[160],stage1_43[205]}
   );
   gpc615_5 gpc1735 (
      {stage0_43[470], stage0_43[471], stage0_43[472], stage0_43[473], stage0_43[474]},
      {stage0_44[189]},
      {stage0_45[348], stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353]},
      {stage1_47[58],stage1_46[82],stage1_45[107],stage1_44[161],stage1_43[206]}
   );
   gpc606_5 gpc1736 (
      {stage0_44[190], stage0_44[191], stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[59],stage1_46[83],stage1_45[108],stage1_44[162]}
   );
   gpc606_5 gpc1737 (
      {stage0_44[196], stage0_44[197], stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[60],stage1_46[84],stage1_45[109],stage1_44[163]}
   );
   gpc606_5 gpc1738 (
      {stage0_44[202], stage0_44[203], stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[61],stage1_46[85],stage1_45[110],stage1_44[164]}
   );
   gpc606_5 gpc1739 (
      {stage0_44[208], stage0_44[209], stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[62],stage1_46[86],stage1_45[111],stage1_44[165]}
   );
   gpc606_5 gpc1740 (
      {stage0_44[214], stage0_44[215], stage0_44[216], stage0_44[217], stage0_44[218], stage0_44[219]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[63],stage1_46[87],stage1_45[112],stage1_44[166]}
   );
   gpc606_5 gpc1741 (
      {stage0_44[220], stage0_44[221], stage0_44[222], stage0_44[223], stage0_44[224], stage0_44[225]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[64],stage1_46[88],stage1_45[113],stage1_44[167]}
   );
   gpc606_5 gpc1742 (
      {stage0_44[226], stage0_44[227], stage0_44[228], stage0_44[229], stage0_44[230], stage0_44[231]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[65],stage1_46[89],stage1_45[114],stage1_44[168]}
   );
   gpc606_5 gpc1743 (
      {stage0_44[232], stage0_44[233], stage0_44[234], stage0_44[235], stage0_44[236], stage0_44[237]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[66],stage1_46[90],stage1_45[115],stage1_44[169]}
   );
   gpc606_5 gpc1744 (
      {stage0_44[238], stage0_44[239], stage0_44[240], stage0_44[241], stage0_44[242], stage0_44[243]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[67],stage1_46[91],stage1_45[116],stage1_44[170]}
   );
   gpc606_5 gpc1745 (
      {stage0_44[244], stage0_44[245], stage0_44[246], stage0_44[247], stage0_44[248], stage0_44[249]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[68],stage1_46[92],stage1_45[117],stage1_44[171]}
   );
   gpc606_5 gpc1746 (
      {stage0_44[250], stage0_44[251], stage0_44[252], stage0_44[253], stage0_44[254], stage0_44[255]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[69],stage1_46[93],stage1_45[118],stage1_44[172]}
   );
   gpc606_5 gpc1747 (
      {stage0_44[256], stage0_44[257], stage0_44[258], stage0_44[259], stage0_44[260], stage0_44[261]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[70],stage1_46[94],stage1_45[119],stage1_44[173]}
   );
   gpc606_5 gpc1748 (
      {stage0_44[262], stage0_44[263], stage0_44[264], stage0_44[265], stage0_44[266], stage0_44[267]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[71],stage1_46[95],stage1_45[120],stage1_44[174]}
   );
   gpc606_5 gpc1749 (
      {stage0_44[268], stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[72],stage1_46[96],stage1_45[121],stage1_44[175]}
   );
   gpc606_5 gpc1750 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278], stage0_44[279]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[73],stage1_46[97],stage1_45[122],stage1_44[176]}
   );
   gpc606_5 gpc1751 (
      {stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283], stage0_44[284], stage0_44[285]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[74],stage1_46[98],stage1_45[123],stage1_44[177]}
   );
   gpc606_5 gpc1752 (
      {stage0_44[286], stage0_44[287], stage0_44[288], stage0_44[289], stage0_44[290], stage0_44[291]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[75],stage1_46[99],stage1_45[124],stage1_44[178]}
   );
   gpc606_5 gpc1753 (
      {stage0_44[292], stage0_44[293], stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[76],stage1_46[100],stage1_45[125],stage1_44[179]}
   );
   gpc606_5 gpc1754 (
      {stage0_44[298], stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[77],stage1_46[101],stage1_45[126],stage1_44[180]}
   );
   gpc606_5 gpc1755 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308], stage0_44[309]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[78],stage1_46[102],stage1_45[127],stage1_44[181]}
   );
   gpc606_5 gpc1756 (
      {stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313], stage0_44[314], stage0_44[315]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[79],stage1_46[103],stage1_45[128],stage1_44[182]}
   );
   gpc606_5 gpc1757 (
      {stage0_44[316], stage0_44[317], stage0_44[318], stage0_44[319], stage0_44[320], stage0_44[321]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[80],stage1_46[104],stage1_45[129],stage1_44[183]}
   );
   gpc606_5 gpc1758 (
      {stage0_44[322], stage0_44[323], stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[81],stage1_46[105],stage1_45[130],stage1_44[184]}
   );
   gpc606_5 gpc1759 (
      {stage0_44[328], stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[82],stage1_46[106],stage1_45[131],stage1_44[185]}
   );
   gpc606_5 gpc1760 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338], stage0_44[339]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[83],stage1_46[107],stage1_45[132],stage1_44[186]}
   );
   gpc606_5 gpc1761 (
      {stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343], stage0_44[344], stage0_44[345]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[84],stage1_46[108],stage1_45[133],stage1_44[187]}
   );
   gpc606_5 gpc1762 (
      {stage0_44[346], stage0_44[347], stage0_44[348], stage0_44[349], stage0_44[350], stage0_44[351]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[85],stage1_46[109],stage1_45[134],stage1_44[188]}
   );
   gpc606_5 gpc1763 (
      {stage0_44[352], stage0_44[353], stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[86],stage1_46[110],stage1_45[135],stage1_44[189]}
   );
   gpc606_5 gpc1764 (
      {stage0_44[358], stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[87],stage1_46[111],stage1_45[136],stage1_44[190]}
   );
   gpc606_5 gpc1765 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368], stage0_44[369]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[88],stage1_46[112],stage1_45[137],stage1_44[191]}
   );
   gpc606_5 gpc1766 (
      {stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373], stage0_44[374], stage0_44[375]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[89],stage1_46[113],stage1_45[138],stage1_44[192]}
   );
   gpc606_5 gpc1767 (
      {stage0_44[376], stage0_44[377], stage0_44[378], stage0_44[379], stage0_44[380], stage0_44[381]},
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190], stage0_46[191]},
      {stage1_48[31],stage1_47[90],stage1_46[114],stage1_45[139],stage1_44[193]}
   );
   gpc606_5 gpc1768 (
      {stage0_44[382], stage0_44[383], stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387]},
      {stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195], stage0_46[196], stage0_46[197]},
      {stage1_48[32],stage1_47[91],stage1_46[115],stage1_45[140],stage1_44[194]}
   );
   gpc606_5 gpc1769 (
      {stage0_44[388], stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_46[198], stage0_46[199], stage0_46[200], stage0_46[201], stage0_46[202], stage0_46[203]},
      {stage1_48[33],stage1_47[92],stage1_46[116],stage1_45[141],stage1_44[195]}
   );
   gpc606_5 gpc1770 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398], stage0_44[399]},
      {stage0_46[204], stage0_46[205], stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209]},
      {stage1_48[34],stage1_47[93],stage1_46[117],stage1_45[142],stage1_44[196]}
   );
   gpc606_5 gpc1771 (
      {stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403], stage0_44[404], stage0_44[405]},
      {stage0_46[210], stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage1_48[35],stage1_47[94],stage1_46[118],stage1_45[143],stage1_44[197]}
   );
   gpc606_5 gpc1772 (
      {stage0_44[406], stage0_44[407], stage0_44[408], stage0_44[409], stage0_44[410], stage0_44[411]},
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220], stage0_46[221]},
      {stage1_48[36],stage1_47[95],stage1_46[119],stage1_45[144],stage1_44[198]}
   );
   gpc606_5 gpc1773 (
      {stage0_44[412], stage0_44[413], stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417]},
      {stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225], stage0_46[226], stage0_46[227]},
      {stage1_48[37],stage1_47[96],stage1_46[120],stage1_45[145],stage1_44[199]}
   );
   gpc606_5 gpc1774 (
      {stage0_44[418], stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_46[228], stage0_46[229], stage0_46[230], stage0_46[231], stage0_46[232], stage0_46[233]},
      {stage1_48[38],stage1_47[97],stage1_46[121],stage1_45[146],stage1_44[200]}
   );
   gpc606_5 gpc1775 (
      {stage0_44[424], stage0_44[425], stage0_44[426], stage0_44[427], stage0_44[428], stage0_44[429]},
      {stage0_46[234], stage0_46[235], stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239]},
      {stage1_48[39],stage1_47[98],stage1_46[122],stage1_45[147],stage1_44[201]}
   );
   gpc606_5 gpc1776 (
      {stage0_44[430], stage0_44[431], stage0_44[432], stage0_44[433], stage0_44[434], stage0_44[435]},
      {stage0_46[240], stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage1_48[40],stage1_47[99],stage1_46[123],stage1_45[148],stage1_44[202]}
   );
   gpc606_5 gpc1777 (
      {stage0_44[436], stage0_44[437], stage0_44[438], stage0_44[439], stage0_44[440], stage0_44[441]},
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250], stage0_46[251]},
      {stage1_48[41],stage1_47[100],stage1_46[124],stage1_45[149],stage1_44[203]}
   );
   gpc606_5 gpc1778 (
      {stage0_44[442], stage0_44[443], stage0_44[444], stage0_44[445], stage0_44[446], stage0_44[447]},
      {stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255], stage0_46[256], stage0_46[257]},
      {stage1_48[42],stage1_47[101],stage1_46[125],stage1_45[150],stage1_44[204]}
   );
   gpc606_5 gpc1779 (
      {stage0_45[354], stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[43],stage1_47[102],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1780 (
      {stage0_45[360], stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[44],stage1_47[103],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1781 (
      {stage0_45[366], stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[45],stage1_47[104],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1782 (
      {stage0_45[372], stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[46],stage1_47[105],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1783 (
      {stage0_45[378], stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[47],stage1_47[106],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1784 (
      {stage0_45[384], stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[48],stage1_47[107],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1785 (
      {stage0_45[390], stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[49],stage1_47[108],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1786 (
      {stage0_45[396], stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[50],stage1_47[109],stage1_46[133],stage1_45[158]}
   );
   gpc606_5 gpc1787 (
      {stage0_45[402], stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[51],stage1_47[110],stage1_46[134],stage1_45[159]}
   );
   gpc606_5 gpc1788 (
      {stage0_45[408], stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[52],stage1_47[111],stage1_46[135],stage1_45[160]}
   );
   gpc606_5 gpc1789 (
      {stage0_45[414], stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[53],stage1_47[112],stage1_46[136],stage1_45[161]}
   );
   gpc606_5 gpc1790 (
      {stage0_45[420], stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[54],stage1_47[113],stage1_46[137],stage1_45[162]}
   );
   gpc606_5 gpc1791 (
      {stage0_45[426], stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[55],stage1_47[114],stage1_46[138],stage1_45[163]}
   );
   gpc606_5 gpc1792 (
      {stage0_45[432], stage0_45[433], stage0_45[434], stage0_45[435], stage0_45[436], stage0_45[437]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[56],stage1_47[115],stage1_46[139],stage1_45[164]}
   );
   gpc606_5 gpc1793 (
      {stage0_45[438], stage0_45[439], stage0_45[440], stage0_45[441], stage0_45[442], stage0_45[443]},
      {stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage1_49[14],stage1_48[57],stage1_47[116],stage1_46[140],stage1_45[165]}
   );
   gpc606_5 gpc1794 (
      {stage0_45[444], stage0_45[445], stage0_45[446], stage0_45[447], stage0_45[448], stage0_45[449]},
      {stage0_47[90], stage0_47[91], stage0_47[92], stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage1_49[15],stage1_48[58],stage1_47[117],stage1_46[141],stage1_45[166]}
   );
   gpc606_5 gpc1795 (
      {stage0_45[450], stage0_45[451], stage0_45[452], stage0_45[453], stage0_45[454], stage0_45[455]},
      {stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage1_49[16],stage1_48[59],stage1_47[118],stage1_46[142],stage1_45[167]}
   );
   gpc606_5 gpc1796 (
      {stage0_45[456], stage0_45[457], stage0_45[458], stage0_45[459], stage0_45[460], stage0_45[461]},
      {stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage1_49[17],stage1_48[60],stage1_47[119],stage1_46[143],stage1_45[168]}
   );
   gpc606_5 gpc1797 (
      {stage0_45[462], stage0_45[463], stage0_45[464], stage0_45[465], stage0_45[466], stage0_45[467]},
      {stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage1_49[18],stage1_48[61],stage1_47[120],stage1_46[144],stage1_45[169]}
   );
   gpc606_5 gpc1798 (
      {stage0_45[468], stage0_45[469], stage0_45[470], stage0_45[471], stage0_45[472], stage0_45[473]},
      {stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117], stage0_47[118], stage0_47[119]},
      {stage1_49[19],stage1_48[62],stage1_47[121],stage1_46[145],stage1_45[170]}
   );
   gpc606_5 gpc1799 (
      {stage0_45[474], stage0_45[475], stage0_45[476], stage0_45[477], stage0_45[478], stage0_45[479]},
      {stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123], stage0_47[124], stage0_47[125]},
      {stage1_49[20],stage1_48[63],stage1_47[122],stage1_46[146],stage1_45[171]}
   );
   gpc606_5 gpc1800 (
      {stage0_45[480], stage0_45[481], stage0_45[482], stage0_45[483], stage0_45[484], stage0_45[485]},
      {stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129], stage0_47[130], stage0_47[131]},
      {stage1_49[21],stage1_48[64],stage1_47[123],stage1_46[147],stage1_45[172]}
   );
   gpc606_5 gpc1801 (
      {stage0_45[486], stage0_45[487], stage0_45[488], stage0_45[489], stage0_45[490], stage0_45[491]},
      {stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135], stage0_47[136], stage0_47[137]},
      {stage1_49[22],stage1_48[65],stage1_47[124],stage1_46[148],stage1_45[173]}
   );
   gpc606_5 gpc1802 (
      {stage0_45[492], stage0_45[493], stage0_45[494], stage0_45[495], stage0_45[496], stage0_45[497]},
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142], stage0_47[143]},
      {stage1_49[23],stage1_48[66],stage1_47[125],stage1_46[149],stage1_45[174]}
   );
   gpc615_5 gpc1803 (
      {stage0_46[258], stage0_46[259], stage0_46[260], stage0_46[261], stage0_46[262]},
      {stage0_47[144]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[24],stage1_48[67],stage1_47[126],stage1_46[150]}
   );
   gpc615_5 gpc1804 (
      {stage0_46[263], stage0_46[264], stage0_46[265], stage0_46[266], stage0_46[267]},
      {stage0_47[145]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[25],stage1_48[68],stage1_47[127],stage1_46[151]}
   );
   gpc615_5 gpc1805 (
      {stage0_46[268], stage0_46[269], stage0_46[270], stage0_46[271], stage0_46[272]},
      {stage0_47[146]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[26],stage1_48[69],stage1_47[128],stage1_46[152]}
   );
   gpc615_5 gpc1806 (
      {stage0_46[273], stage0_46[274], stage0_46[275], stage0_46[276], stage0_46[277]},
      {stage0_47[147]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[27],stage1_48[70],stage1_47[129],stage1_46[153]}
   );
   gpc615_5 gpc1807 (
      {stage0_46[278], stage0_46[279], stage0_46[280], stage0_46[281], stage0_46[282]},
      {stage0_47[148]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[28],stage1_48[71],stage1_47[130],stage1_46[154]}
   );
   gpc615_5 gpc1808 (
      {stage0_46[283], stage0_46[284], stage0_46[285], stage0_46[286], stage0_46[287]},
      {stage0_47[149]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[29],stage1_48[72],stage1_47[131],stage1_46[155]}
   );
   gpc615_5 gpc1809 (
      {stage0_46[288], stage0_46[289], stage0_46[290], stage0_46[291], stage0_46[292]},
      {stage0_47[150]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[30],stage1_48[73],stage1_47[132],stage1_46[156]}
   );
   gpc615_5 gpc1810 (
      {stage0_46[293], stage0_46[294], stage0_46[295], stage0_46[296], stage0_46[297]},
      {stage0_47[151]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[31],stage1_48[74],stage1_47[133],stage1_46[157]}
   );
   gpc615_5 gpc1811 (
      {stage0_46[298], stage0_46[299], stage0_46[300], stage0_46[301], stage0_46[302]},
      {stage0_47[152]},
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage1_50[8],stage1_49[32],stage1_48[75],stage1_47[134],stage1_46[158]}
   );
   gpc615_5 gpc1812 (
      {stage0_46[303], stage0_46[304], stage0_46[305], stage0_46[306], stage0_46[307]},
      {stage0_47[153]},
      {stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58], stage0_48[59]},
      {stage1_50[9],stage1_49[33],stage1_48[76],stage1_47[135],stage1_46[159]}
   );
   gpc615_5 gpc1813 (
      {stage0_46[308], stage0_46[309], stage0_46[310], stage0_46[311], stage0_46[312]},
      {stage0_47[154]},
      {stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64], stage0_48[65]},
      {stage1_50[10],stage1_49[34],stage1_48[77],stage1_47[136],stage1_46[160]}
   );
   gpc615_5 gpc1814 (
      {stage0_46[313], stage0_46[314], stage0_46[315], stage0_46[316], stage0_46[317]},
      {stage0_47[155]},
      {stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70], stage0_48[71]},
      {stage1_50[11],stage1_49[35],stage1_48[78],stage1_47[137],stage1_46[161]}
   );
   gpc615_5 gpc1815 (
      {stage0_46[318], stage0_46[319], stage0_46[320], stage0_46[321], stage0_46[322]},
      {stage0_47[156]},
      {stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75], stage0_48[76], stage0_48[77]},
      {stage1_50[12],stage1_49[36],stage1_48[79],stage1_47[138],stage1_46[162]}
   );
   gpc615_5 gpc1816 (
      {stage0_46[323], stage0_46[324], stage0_46[325], stage0_46[326], stage0_46[327]},
      {stage0_47[157]},
      {stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81], stage0_48[82], stage0_48[83]},
      {stage1_50[13],stage1_49[37],stage1_48[80],stage1_47[139],stage1_46[163]}
   );
   gpc615_5 gpc1817 (
      {stage0_46[328], stage0_46[329], stage0_46[330], stage0_46[331], stage0_46[332]},
      {stage0_47[158]},
      {stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89]},
      {stage1_50[14],stage1_49[38],stage1_48[81],stage1_47[140],stage1_46[164]}
   );
   gpc615_5 gpc1818 (
      {stage0_46[333], stage0_46[334], stage0_46[335], stage0_46[336], stage0_46[337]},
      {stage0_47[159]},
      {stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage1_50[15],stage1_49[39],stage1_48[82],stage1_47[141],stage1_46[165]}
   );
   gpc615_5 gpc1819 (
      {stage0_46[338], stage0_46[339], stage0_46[340], stage0_46[341], stage0_46[342]},
      {stage0_47[160]},
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100], stage0_48[101]},
      {stage1_50[16],stage1_49[40],stage1_48[83],stage1_47[142],stage1_46[166]}
   );
   gpc615_5 gpc1820 (
      {stage0_46[343], stage0_46[344], stage0_46[345], stage0_46[346], stage0_46[347]},
      {stage0_47[161]},
      {stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105], stage0_48[106], stage0_48[107]},
      {stage1_50[17],stage1_49[41],stage1_48[84],stage1_47[143],stage1_46[167]}
   );
   gpc615_5 gpc1821 (
      {stage0_46[348], stage0_46[349], stage0_46[350], stage0_46[351], stage0_46[352]},
      {stage0_47[162]},
      {stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111], stage0_48[112], stage0_48[113]},
      {stage1_50[18],stage1_49[42],stage1_48[85],stage1_47[144],stage1_46[168]}
   );
   gpc615_5 gpc1822 (
      {stage0_46[353], stage0_46[354], stage0_46[355], stage0_46[356], stage0_46[357]},
      {stage0_47[163]},
      {stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119]},
      {stage1_50[19],stage1_49[43],stage1_48[86],stage1_47[145],stage1_46[169]}
   );
   gpc615_5 gpc1823 (
      {stage0_46[358], stage0_46[359], stage0_46[360], stage0_46[361], stage0_46[362]},
      {stage0_47[164]},
      {stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage1_50[20],stage1_49[44],stage1_48[87],stage1_47[146],stage1_46[170]}
   );
   gpc615_5 gpc1824 (
      {stage0_46[363], stage0_46[364], stage0_46[365], stage0_46[366], stage0_46[367]},
      {stage0_47[165]},
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130], stage0_48[131]},
      {stage1_50[21],stage1_49[45],stage1_48[88],stage1_47[147],stage1_46[171]}
   );
   gpc615_5 gpc1825 (
      {stage0_46[368], stage0_46[369], stage0_46[370], stage0_46[371], stage0_46[372]},
      {stage0_47[166]},
      {stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135], stage0_48[136], stage0_48[137]},
      {stage1_50[22],stage1_49[46],stage1_48[89],stage1_47[148],stage1_46[172]}
   );
   gpc615_5 gpc1826 (
      {stage0_46[373], stage0_46[374], stage0_46[375], stage0_46[376], stage0_46[377]},
      {stage0_47[167]},
      {stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141], stage0_48[142], stage0_48[143]},
      {stage1_50[23],stage1_49[47],stage1_48[90],stage1_47[149],stage1_46[173]}
   );
   gpc615_5 gpc1827 (
      {stage0_46[378], stage0_46[379], stage0_46[380], stage0_46[381], stage0_46[382]},
      {stage0_47[168]},
      {stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149]},
      {stage1_50[24],stage1_49[48],stage1_48[91],stage1_47[150],stage1_46[174]}
   );
   gpc615_5 gpc1828 (
      {stage0_46[383], stage0_46[384], stage0_46[385], stage0_46[386], stage0_46[387]},
      {stage0_47[169]},
      {stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage1_50[25],stage1_49[49],stage1_48[92],stage1_47[151],stage1_46[175]}
   );
   gpc606_5 gpc1829 (
      {stage0_47[170], stage0_47[171], stage0_47[172], stage0_47[173], stage0_47[174], stage0_47[175]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[26],stage1_49[50],stage1_48[93],stage1_47[152]}
   );
   gpc606_5 gpc1830 (
      {stage0_47[176], stage0_47[177], stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[27],stage1_49[51],stage1_48[94],stage1_47[153]}
   );
   gpc606_5 gpc1831 (
      {stage0_47[182], stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[28],stage1_49[52],stage1_48[95],stage1_47[154]}
   );
   gpc606_5 gpc1832 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192], stage0_47[193]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[29],stage1_49[53],stage1_48[96],stage1_47[155]}
   );
   gpc606_5 gpc1833 (
      {stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197], stage0_47[198], stage0_47[199]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[30],stage1_49[54],stage1_48[97],stage1_47[156]}
   );
   gpc606_5 gpc1834 (
      {stage0_47[200], stage0_47[201], stage0_47[202], stage0_47[203], stage0_47[204], stage0_47[205]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[31],stage1_49[55],stage1_48[98],stage1_47[157]}
   );
   gpc606_5 gpc1835 (
      {stage0_47[206], stage0_47[207], stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[32],stage1_49[56],stage1_48[99],stage1_47[158]}
   );
   gpc606_5 gpc1836 (
      {stage0_47[212], stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[33],stage1_49[57],stage1_48[100],stage1_47[159]}
   );
   gpc606_5 gpc1837 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222], stage0_47[223]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[34],stage1_49[58],stage1_48[101],stage1_47[160]}
   );
   gpc606_5 gpc1838 (
      {stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227], stage0_47[228], stage0_47[229]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[35],stage1_49[59],stage1_48[102],stage1_47[161]}
   );
   gpc606_5 gpc1839 (
      {stage0_47[230], stage0_47[231], stage0_47[232], stage0_47[233], stage0_47[234], stage0_47[235]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[36],stage1_49[60],stage1_48[103],stage1_47[162]}
   );
   gpc606_5 gpc1840 (
      {stage0_47[236], stage0_47[237], stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[37],stage1_49[61],stage1_48[104],stage1_47[163]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[242], stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246]},
      {stage0_48[156]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[38],stage1_49[62],stage1_48[105],stage1_47[164]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[247], stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251]},
      {stage0_48[157]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[39],stage1_49[63],stage1_48[106],stage1_47[165]}
   );
   gpc615_5 gpc1843 (
      {stage0_47[252], stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256]},
      {stage0_48[158]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[40],stage1_49[64],stage1_48[107],stage1_47[166]}
   );
   gpc615_5 gpc1844 (
      {stage0_47[257], stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261]},
      {stage0_48[159]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[41],stage1_49[65],stage1_48[108],stage1_47[167]}
   );
   gpc615_5 gpc1845 (
      {stage0_47[262], stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266]},
      {stage0_48[160]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[42],stage1_49[66],stage1_48[109],stage1_47[168]}
   );
   gpc615_5 gpc1846 (
      {stage0_47[267], stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271]},
      {stage0_48[161]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[43],stage1_49[67],stage1_48[110],stage1_47[169]}
   );
   gpc615_5 gpc1847 (
      {stage0_47[272], stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276]},
      {stage0_48[162]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[44],stage1_49[68],stage1_48[111],stage1_47[170]}
   );
   gpc615_5 gpc1848 (
      {stage0_47[277], stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281]},
      {stage0_48[163]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[45],stage1_49[69],stage1_48[112],stage1_47[171]}
   );
   gpc615_5 gpc1849 (
      {stage0_47[282], stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286]},
      {stage0_48[164]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[46],stage1_49[70],stage1_48[113],stage1_47[172]}
   );
   gpc615_5 gpc1850 (
      {stage0_47[287], stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291]},
      {stage0_48[165]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[47],stage1_49[71],stage1_48[114],stage1_47[173]}
   );
   gpc615_5 gpc1851 (
      {stage0_47[292], stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296]},
      {stage0_48[166]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[48],stage1_49[72],stage1_48[115],stage1_47[174]}
   );
   gpc615_5 gpc1852 (
      {stage0_47[297], stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301]},
      {stage0_48[167]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[49],stage1_49[73],stage1_48[116],stage1_47[175]}
   );
   gpc615_5 gpc1853 (
      {stage0_47[302], stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306]},
      {stage0_48[168]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[50],stage1_49[74],stage1_48[117],stage1_47[176]}
   );
   gpc615_5 gpc1854 (
      {stage0_47[307], stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311]},
      {stage0_48[169]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[51],stage1_49[75],stage1_48[118],stage1_47[177]}
   );
   gpc615_5 gpc1855 (
      {stage0_47[312], stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316]},
      {stage0_48[170]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[52],stage1_49[76],stage1_48[119],stage1_47[178]}
   );
   gpc615_5 gpc1856 (
      {stage0_47[317], stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321]},
      {stage0_48[171]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[53],stage1_49[77],stage1_48[120],stage1_47[179]}
   );
   gpc615_5 gpc1857 (
      {stage0_47[322], stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326]},
      {stage0_48[172]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[54],stage1_49[78],stage1_48[121],stage1_47[180]}
   );
   gpc615_5 gpc1858 (
      {stage0_47[327], stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331]},
      {stage0_48[173]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[55],stage1_49[79],stage1_48[122],stage1_47[181]}
   );
   gpc615_5 gpc1859 (
      {stage0_47[332], stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336]},
      {stage0_48[174]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[56],stage1_49[80],stage1_48[123],stage1_47[182]}
   );
   gpc615_5 gpc1860 (
      {stage0_47[337], stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341]},
      {stage0_48[175]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[57],stage1_49[81],stage1_48[124],stage1_47[183]}
   );
   gpc615_5 gpc1861 (
      {stage0_47[342], stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346]},
      {stage0_48[176]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[58],stage1_49[82],stage1_48[125],stage1_47[184]}
   );
   gpc615_5 gpc1862 (
      {stage0_47[347], stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351]},
      {stage0_48[177]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[59],stage1_49[83],stage1_48[126],stage1_47[185]}
   );
   gpc615_5 gpc1863 (
      {stage0_47[352], stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356]},
      {stage0_48[178]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[60],stage1_49[84],stage1_48[127],stage1_47[186]}
   );
   gpc615_5 gpc1864 (
      {stage0_47[357], stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361]},
      {stage0_48[179]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[61],stage1_49[85],stage1_48[128],stage1_47[187]}
   );
   gpc615_5 gpc1865 (
      {stage0_47[362], stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366]},
      {stage0_48[180]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[62],stage1_49[86],stage1_48[129],stage1_47[188]}
   );
   gpc615_5 gpc1866 (
      {stage0_47[367], stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371]},
      {stage0_48[181]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[63],stage1_49[87],stage1_48[130],stage1_47[189]}
   );
   gpc615_5 gpc1867 (
      {stage0_47[372], stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376]},
      {stage0_48[182]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[64],stage1_49[88],stage1_48[131],stage1_47[190]}
   );
   gpc615_5 gpc1868 (
      {stage0_47[377], stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381]},
      {stage0_48[183]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[65],stage1_49[89],stage1_48[132],stage1_47[191]}
   );
   gpc615_5 gpc1869 (
      {stage0_47[382], stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386]},
      {stage0_48[184]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[66],stage1_49[90],stage1_48[133],stage1_47[192]}
   );
   gpc615_5 gpc1870 (
      {stage0_47[387], stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391]},
      {stage0_48[185]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[67],stage1_49[91],stage1_48[134],stage1_47[193]}
   );
   gpc615_5 gpc1871 (
      {stage0_47[392], stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396]},
      {stage0_48[186]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[68],stage1_49[92],stage1_48[135],stage1_47[194]}
   );
   gpc615_5 gpc1872 (
      {stage0_47[397], stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401]},
      {stage0_48[187]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[69],stage1_49[93],stage1_48[136],stage1_47[195]}
   );
   gpc615_5 gpc1873 (
      {stage0_47[402], stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406]},
      {stage0_48[188]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[70],stage1_49[94],stage1_48[137],stage1_47[196]}
   );
   gpc615_5 gpc1874 (
      {stage0_47[407], stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411]},
      {stage0_48[189]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[71],stage1_49[95],stage1_48[138],stage1_47[197]}
   );
   gpc615_5 gpc1875 (
      {stage0_47[412], stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416]},
      {stage0_48[190]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[72],stage1_49[96],stage1_48[139],stage1_47[198]}
   );
   gpc615_5 gpc1876 (
      {stage0_47[417], stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421]},
      {stage0_48[191]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[73],stage1_49[97],stage1_48[140],stage1_47[199]}
   );
   gpc615_5 gpc1877 (
      {stage0_47[422], stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426]},
      {stage0_48[192]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[74],stage1_49[98],stage1_48[141],stage1_47[200]}
   );
   gpc615_5 gpc1878 (
      {stage0_47[427], stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431]},
      {stage0_48[193]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[75],stage1_49[99],stage1_48[142],stage1_47[201]}
   );
   gpc615_5 gpc1879 (
      {stage0_47[432], stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436]},
      {stage0_48[194]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[76],stage1_49[100],stage1_48[143],stage1_47[202]}
   );
   gpc606_5 gpc1880 (
      {stage0_48[195], stage0_48[196], stage0_48[197], stage0_48[198], stage0_48[199], stage0_48[200]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[51],stage1_50[77],stage1_49[101],stage1_48[144]}
   );
   gpc606_5 gpc1881 (
      {stage0_48[201], stage0_48[202], stage0_48[203], stage0_48[204], stage0_48[205], stage0_48[206]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[52],stage1_50[78],stage1_49[102],stage1_48[145]}
   );
   gpc606_5 gpc1882 (
      {stage0_48[207], stage0_48[208], stage0_48[209], stage0_48[210], stage0_48[211], stage0_48[212]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[53],stage1_50[79],stage1_49[103],stage1_48[146]}
   );
   gpc606_5 gpc1883 (
      {stage0_48[213], stage0_48[214], stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[54],stage1_50[80],stage1_49[104],stage1_48[147]}
   );
   gpc606_5 gpc1884 (
      {stage0_48[219], stage0_48[220], stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[55],stage1_50[81],stage1_49[105],stage1_48[148]}
   );
   gpc606_5 gpc1885 (
      {stage0_48[225], stage0_48[226], stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[56],stage1_50[82],stage1_49[106],stage1_48[149]}
   );
   gpc606_5 gpc1886 (
      {stage0_48[231], stage0_48[232], stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[57],stage1_50[83],stage1_49[107],stage1_48[150]}
   );
   gpc606_5 gpc1887 (
      {stage0_48[237], stage0_48[238], stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[58],stage1_50[84],stage1_49[108],stage1_48[151]}
   );
   gpc606_5 gpc1888 (
      {stage0_48[243], stage0_48[244], stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[59],stage1_50[85],stage1_49[109],stage1_48[152]}
   );
   gpc606_5 gpc1889 (
      {stage0_48[249], stage0_48[250], stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[60],stage1_50[86],stage1_49[110],stage1_48[153]}
   );
   gpc606_5 gpc1890 (
      {stage0_48[255], stage0_48[256], stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[61],stage1_50[87],stage1_49[111],stage1_48[154]}
   );
   gpc606_5 gpc1891 (
      {stage0_48[261], stage0_48[262], stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[62],stage1_50[88],stage1_49[112],stage1_48[155]}
   );
   gpc606_5 gpc1892 (
      {stage0_48[267], stage0_48[268], stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[63],stage1_50[89],stage1_49[113],stage1_48[156]}
   );
   gpc606_5 gpc1893 (
      {stage0_48[273], stage0_48[274], stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[64],stage1_50[90],stage1_49[114],stage1_48[157]}
   );
   gpc606_5 gpc1894 (
      {stage0_48[279], stage0_48[280], stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[65],stage1_50[91],stage1_49[115],stage1_48[158]}
   );
   gpc606_5 gpc1895 (
      {stage0_48[285], stage0_48[286], stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[66],stage1_50[92],stage1_49[116],stage1_48[159]}
   );
   gpc606_5 gpc1896 (
      {stage0_48[291], stage0_48[292], stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[67],stage1_50[93],stage1_49[117],stage1_48[160]}
   );
   gpc606_5 gpc1897 (
      {stage0_48[297], stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[68],stage1_50[94],stage1_49[118],stage1_48[161]}
   );
   gpc606_5 gpc1898 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307], stage0_48[308]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[69],stage1_50[95],stage1_49[119],stage1_48[162]}
   );
   gpc606_5 gpc1899 (
      {stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312], stage0_48[313], stage0_48[314]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[70],stage1_50[96],stage1_49[120],stage1_48[163]}
   );
   gpc606_5 gpc1900 (
      {stage0_48[315], stage0_48[316], stage0_48[317], stage0_48[318], stage0_48[319], stage0_48[320]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[71],stage1_50[97],stage1_49[121],stage1_48[164]}
   );
   gpc606_5 gpc1901 (
      {stage0_48[321], stage0_48[322], stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[72],stage1_50[98],stage1_49[122],stage1_48[165]}
   );
   gpc606_5 gpc1902 (
      {stage0_48[327], stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[73],stage1_50[99],stage1_49[123],stage1_48[166]}
   );
   gpc606_5 gpc1903 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337], stage0_48[338]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[74],stage1_50[100],stage1_49[124],stage1_48[167]}
   );
   gpc606_5 gpc1904 (
      {stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342], stage0_48[343], stage0_48[344]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[75],stage1_50[101],stage1_49[125],stage1_48[168]}
   );
   gpc606_5 gpc1905 (
      {stage0_48[345], stage0_48[346], stage0_48[347], stage0_48[348], stage0_48[349], stage0_48[350]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[76],stage1_50[102],stage1_49[126],stage1_48[169]}
   );
   gpc606_5 gpc1906 (
      {stage0_48[351], stage0_48[352], stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[77],stage1_50[103],stage1_49[127],stage1_48[170]}
   );
   gpc606_5 gpc1907 (
      {stage0_48[357], stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[78],stage1_50[104],stage1_49[128],stage1_48[171]}
   );
   gpc606_5 gpc1908 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367], stage0_48[368]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[79],stage1_50[105],stage1_49[129],stage1_48[172]}
   );
   gpc606_5 gpc1909 (
      {stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372], stage0_48[373], stage0_48[374]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[80],stage1_50[106],stage1_49[130],stage1_48[173]}
   );
   gpc606_5 gpc1910 (
      {stage0_48[375], stage0_48[376], stage0_48[377], stage0_48[378], stage0_48[379], stage0_48[380]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[81],stage1_50[107],stage1_49[131],stage1_48[174]}
   );
   gpc606_5 gpc1911 (
      {stage0_48[381], stage0_48[382], stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[82],stage1_50[108],stage1_49[132],stage1_48[175]}
   );
   gpc606_5 gpc1912 (
      {stage0_48[387], stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[83],stage1_50[109],stage1_49[133],stage1_48[176]}
   );
   gpc606_5 gpc1913 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397], stage0_48[398]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[84],stage1_50[110],stage1_49[134],stage1_48[177]}
   );
   gpc606_5 gpc1914 (
      {stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402], stage0_48[403], stage0_48[404]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[85],stage1_50[111],stage1_49[135],stage1_48[178]}
   );
   gpc606_5 gpc1915 (
      {stage0_48[405], stage0_48[406], stage0_48[407], stage0_48[408], stage0_48[409], stage0_48[410]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[86],stage1_50[112],stage1_49[136],stage1_48[179]}
   );
   gpc606_5 gpc1916 (
      {stage0_48[411], stage0_48[412], stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[87],stage1_50[113],stage1_49[137],stage1_48[180]}
   );
   gpc606_5 gpc1917 (
      {stage0_48[417], stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[88],stage1_50[114],stage1_49[138],stage1_48[181]}
   );
   gpc606_5 gpc1918 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427], stage0_48[428]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[89],stage1_50[115],stage1_49[139],stage1_48[182]}
   );
   gpc606_5 gpc1919 (
      {stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432], stage0_48[433], stage0_48[434]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[90],stage1_50[116],stage1_49[140],stage1_48[183]}
   );
   gpc606_5 gpc1920 (
      {stage0_48[435], stage0_48[436], stage0_48[437], stage0_48[438], stage0_48[439], stage0_48[440]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[91],stage1_50[117],stage1_49[141],stage1_48[184]}
   );
   gpc606_5 gpc1921 (
      {stage0_48[441], stage0_48[442], stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[92],stage1_50[118],stage1_49[142],stage1_48[185]}
   );
   gpc606_5 gpc1922 (
      {stage0_48[447], stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[93],stage1_50[119],stage1_49[143],stage1_48[186]}
   );
   gpc606_5 gpc1923 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457], stage0_48[458]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[94],stage1_50[120],stage1_49[144],stage1_48[187]}
   );
   gpc606_5 gpc1924 (
      {stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462], stage0_48[463], stage0_48[464]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[95],stage1_50[121],stage1_49[145],stage1_48[188]}
   );
   gpc606_5 gpc1925 (
      {stage0_48[465], stage0_48[466], stage0_48[467], stage0_48[468], stage0_48[469], stage0_48[470]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[96],stage1_50[122],stage1_49[146],stage1_48[189]}
   );
   gpc606_5 gpc1926 (
      {stage0_48[471], stage0_48[472], stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[97],stage1_50[123],stage1_49[147],stage1_48[190]}
   );
   gpc606_5 gpc1927 (
      {stage0_48[477], stage0_48[478], stage0_48[479], stage0_48[480], stage0_48[481], stage0_48[482]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[98],stage1_50[124],stage1_49[148],stage1_48[191]}
   );
   gpc606_5 gpc1928 (
      {stage0_48[483], stage0_48[484], stage0_48[485], stage0_48[486], stage0_48[487], stage0_48[488]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[99],stage1_50[125],stage1_49[149],stage1_48[192]}
   );
   gpc606_5 gpc1929 (
      {stage0_48[489], stage0_48[490], stage0_48[491], stage0_48[492], stage0_48[493], stage0_48[494]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[100],stage1_50[126],stage1_49[150],stage1_48[193]}
   );
   gpc606_5 gpc1930 (
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[101],stage1_50[127],stage1_49[151]}
   );
   gpc606_5 gpc1931 (
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[102],stage1_50[128],stage1_49[152]}
   );
   gpc606_5 gpc1932 (
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[103],stage1_50[129],stage1_49[153]}
   );
   gpc606_5 gpc1933 (
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[104],stage1_50[130],stage1_49[154]}
   );
   gpc606_5 gpc1934 (
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[105],stage1_50[131],stage1_49[155]}
   );
   gpc606_5 gpc1935 (
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[106],stage1_50[132],stage1_49[156]}
   );
   gpc606_5 gpc1936 (
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[107],stage1_50[133],stage1_49[157]}
   );
   gpc606_5 gpc1937 (
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[108],stage1_50[134],stage1_49[158]}
   );
   gpc606_5 gpc1938 (
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[109],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1939 (
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[110],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1940 (
      {stage0_49[366], stage0_49[367], stage0_49[368], stage0_49[369], stage0_49[370], stage0_49[371]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[111],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1941 (
      {stage0_49[372], stage0_49[373], stage0_49[374], stage0_49[375], stage0_49[376], stage0_49[377]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[112],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1942 (
      {stage0_49[378], stage0_49[379], stage0_49[380], stage0_49[381], stage0_49[382], stage0_49[383]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[113],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1943 (
      {stage0_49[384], stage0_49[385], stage0_49[386], stage0_49[387], stage0_49[388], stage0_49[389]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[114],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1944 (
      {stage0_49[390], stage0_49[391], stage0_49[392], stage0_49[393], stage0_49[394], stage0_49[395]},
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage1_53[14],stage1_52[64],stage1_51[115],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1945 (
      {stage0_49[396], stage0_49[397], stage0_49[398], stage0_49[399], stage0_49[400], stage0_49[401]},
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage1_53[15],stage1_52[65],stage1_51[116],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1946 (
      {stage0_49[402], stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407]},
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage1_53[16],stage1_52[66],stage1_51[117],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1947 (
      {stage0_49[408], stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413]},
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage1_53[17],stage1_52[67],stage1_51[118],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1948 (
      {stage0_49[414], stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419]},
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage1_53[18],stage1_52[68],stage1_51[119],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1949 (
      {stage0_49[420], stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425]},
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage1_53[19],stage1_52[69],stage1_51[120],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1950 (
      {stage0_49[426], stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431]},
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage1_53[20],stage1_52[70],stage1_51[121],stage1_50[147],stage1_49[171]}
   );
   gpc606_5 gpc1951 (
      {stage0_49[432], stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437]},
      {stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129], stage0_51[130], stage0_51[131]},
      {stage1_53[21],stage1_52[71],stage1_51[122],stage1_50[148],stage1_49[172]}
   );
   gpc606_5 gpc1952 (
      {stage0_49[438], stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443]},
      {stage0_51[132], stage0_51[133], stage0_51[134], stage0_51[135], stage0_51[136], stage0_51[137]},
      {stage1_53[22],stage1_52[72],stage1_51[123],stage1_50[149],stage1_49[173]}
   );
   gpc606_5 gpc1953 (
      {stage0_50[300], stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[23],stage1_52[73],stage1_51[124],stage1_50[150]}
   );
   gpc606_5 gpc1954 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310], stage0_50[311]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[24],stage1_52[74],stage1_51[125],stage1_50[151]}
   );
   gpc606_5 gpc1955 (
      {stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315], stage0_50[316], stage0_50[317]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[25],stage1_52[75],stage1_51[126],stage1_50[152]}
   );
   gpc606_5 gpc1956 (
      {stage0_50[318], stage0_50[319], stage0_50[320], stage0_50[321], stage0_50[322], stage0_50[323]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[26],stage1_52[76],stage1_51[127],stage1_50[153]}
   );
   gpc606_5 gpc1957 (
      {stage0_50[324], stage0_50[325], stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[27],stage1_52[77],stage1_51[128],stage1_50[154]}
   );
   gpc606_5 gpc1958 (
      {stage0_50[330], stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[28],stage1_52[78],stage1_51[129],stage1_50[155]}
   );
   gpc606_5 gpc1959 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340], stage0_50[341]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[29],stage1_52[79],stage1_51[130],stage1_50[156]}
   );
   gpc606_5 gpc1960 (
      {stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345], stage0_50[346], stage0_50[347]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[30],stage1_52[80],stage1_51[131],stage1_50[157]}
   );
   gpc606_5 gpc1961 (
      {stage0_50[348], stage0_50[349], stage0_50[350], stage0_50[351], stage0_50[352], stage0_50[353]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[31],stage1_52[81],stage1_51[132],stage1_50[158]}
   );
   gpc606_5 gpc1962 (
      {stage0_50[354], stage0_50[355], stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[32],stage1_52[82],stage1_51[133],stage1_50[159]}
   );
   gpc606_5 gpc1963 (
      {stage0_50[360], stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[33],stage1_52[83],stage1_51[134],stage1_50[160]}
   );
   gpc606_5 gpc1964 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370], stage0_50[371]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[34],stage1_52[84],stage1_51[135],stage1_50[161]}
   );
   gpc606_5 gpc1965 (
      {stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375], stage0_50[376], stage0_50[377]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[35],stage1_52[85],stage1_51[136],stage1_50[162]}
   );
   gpc606_5 gpc1966 (
      {stage0_50[378], stage0_50[379], stage0_50[380], stage0_50[381], stage0_50[382], stage0_50[383]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[36],stage1_52[86],stage1_51[137],stage1_50[163]}
   );
   gpc606_5 gpc1967 (
      {stage0_50[384], stage0_50[385], stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[37],stage1_52[87],stage1_51[138],stage1_50[164]}
   );
   gpc606_5 gpc1968 (
      {stage0_50[390], stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[38],stage1_52[88],stage1_51[139],stage1_50[165]}
   );
   gpc606_5 gpc1969 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400], stage0_50[401]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[39],stage1_52[89],stage1_51[140],stage1_50[166]}
   );
   gpc606_5 gpc1970 (
      {stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405], stage0_50[406], stage0_50[407]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[40],stage1_52[90],stage1_51[141],stage1_50[167]}
   );
   gpc606_5 gpc1971 (
      {stage0_50[408], stage0_50[409], stage0_50[410], stage0_50[411], stage0_50[412], stage0_50[413]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[41],stage1_52[91],stage1_51[142],stage1_50[168]}
   );
   gpc606_5 gpc1972 (
      {stage0_50[414], stage0_50[415], stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[42],stage1_52[92],stage1_51[143],stage1_50[169]}
   );
   gpc606_5 gpc1973 (
      {stage0_50[420], stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[43],stage1_52[93],stage1_51[144],stage1_50[170]}
   );
   gpc606_5 gpc1974 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430], stage0_50[431]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[44],stage1_52[94],stage1_51[145],stage1_50[171]}
   );
   gpc606_5 gpc1975 (
      {stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435], stage0_50[436], stage0_50[437]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[45],stage1_52[95],stage1_51[146],stage1_50[172]}
   );
   gpc606_5 gpc1976 (
      {stage0_50[438], stage0_50[439], stage0_50[440], stage0_50[441], stage0_50[442], stage0_50[443]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[46],stage1_52[96],stage1_51[147],stage1_50[173]}
   );
   gpc606_5 gpc1977 (
      {stage0_50[444], stage0_50[445], stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[47],stage1_52[97],stage1_51[148],stage1_50[174]}
   );
   gpc606_5 gpc1978 (
      {stage0_50[450], stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[48],stage1_52[98],stage1_51[149],stage1_50[175]}
   );
   gpc606_5 gpc1979 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460], stage0_50[461]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[49],stage1_52[99],stage1_51[150],stage1_50[176]}
   );
   gpc606_5 gpc1980 (
      {stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465], stage0_50[466], stage0_50[467]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[50],stage1_52[100],stage1_51[151],stage1_50[177]}
   );
   gpc606_5 gpc1981 (
      {stage0_50[468], stage0_50[469], stage0_50[470], stage0_50[471], stage0_50[472], stage0_50[473]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[51],stage1_52[101],stage1_51[152],stage1_50[178]}
   );
   gpc606_5 gpc1982 (
      {stage0_51[138], stage0_51[139], stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[29],stage1_53[52],stage1_52[102],stage1_51[153]}
   );
   gpc606_5 gpc1983 (
      {stage0_51[144], stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[30],stage1_53[53],stage1_52[103],stage1_51[154]}
   );
   gpc606_5 gpc1984 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154], stage0_51[155]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[31],stage1_53[54],stage1_52[104],stage1_51[155]}
   );
   gpc606_5 gpc1985 (
      {stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159], stage0_51[160], stage0_51[161]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[32],stage1_53[55],stage1_52[105],stage1_51[156]}
   );
   gpc606_5 gpc1986 (
      {stage0_51[162], stage0_51[163], stage0_51[164], stage0_51[165], stage0_51[166], stage0_51[167]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[33],stage1_53[56],stage1_52[106],stage1_51[157]}
   );
   gpc606_5 gpc1987 (
      {stage0_51[168], stage0_51[169], stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[34],stage1_53[57],stage1_52[107],stage1_51[158]}
   );
   gpc606_5 gpc1988 (
      {stage0_51[174], stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[35],stage1_53[58],stage1_52[108],stage1_51[159]}
   );
   gpc606_5 gpc1989 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184], stage0_51[185]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[36],stage1_53[59],stage1_52[109],stage1_51[160]}
   );
   gpc606_5 gpc1990 (
      {stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189], stage0_51[190], stage0_51[191]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[37],stage1_53[60],stage1_52[110],stage1_51[161]}
   );
   gpc606_5 gpc1991 (
      {stage0_51[192], stage0_51[193], stage0_51[194], stage0_51[195], stage0_51[196], stage0_51[197]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[38],stage1_53[61],stage1_52[111],stage1_51[162]}
   );
   gpc606_5 gpc1992 (
      {stage0_51[198], stage0_51[199], stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[39],stage1_53[62],stage1_52[112],stage1_51[163]}
   );
   gpc606_5 gpc1993 (
      {stage0_51[204], stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[40],stage1_53[63],stage1_52[113],stage1_51[164]}
   );
   gpc606_5 gpc1994 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214], stage0_51[215]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[41],stage1_53[64],stage1_52[114],stage1_51[165]}
   );
   gpc606_5 gpc1995 (
      {stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219], stage0_51[220], stage0_51[221]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[42],stage1_53[65],stage1_52[115],stage1_51[166]}
   );
   gpc606_5 gpc1996 (
      {stage0_51[222], stage0_51[223], stage0_51[224], stage0_51[225], stage0_51[226], stage0_51[227]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[43],stage1_53[66],stage1_52[116],stage1_51[167]}
   );
   gpc606_5 gpc1997 (
      {stage0_51[228], stage0_51[229], stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[44],stage1_53[67],stage1_52[117],stage1_51[168]}
   );
   gpc606_5 gpc1998 (
      {stage0_51[234], stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[45],stage1_53[68],stage1_52[118],stage1_51[169]}
   );
   gpc606_5 gpc1999 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244], stage0_51[245]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[46],stage1_53[69],stage1_52[119],stage1_51[170]}
   );
   gpc606_5 gpc2000 (
      {stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249], stage0_51[250], stage0_51[251]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[47],stage1_53[70],stage1_52[120],stage1_51[171]}
   );
   gpc606_5 gpc2001 (
      {stage0_51[252], stage0_51[253], stage0_51[254], stage0_51[255], stage0_51[256], stage0_51[257]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[48],stage1_53[71],stage1_52[121],stage1_51[172]}
   );
   gpc606_5 gpc2002 (
      {stage0_51[258], stage0_51[259], stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[49],stage1_53[72],stage1_52[122],stage1_51[173]}
   );
   gpc606_5 gpc2003 (
      {stage0_51[264], stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[50],stage1_53[73],stage1_52[123],stage1_51[174]}
   );
   gpc606_5 gpc2004 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274], stage0_51[275]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[51],stage1_53[74],stage1_52[124],stage1_51[175]}
   );
   gpc606_5 gpc2005 (
      {stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279], stage0_51[280], stage0_51[281]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[52],stage1_53[75],stage1_52[125],stage1_51[176]}
   );
   gpc606_5 gpc2006 (
      {stage0_51[282], stage0_51[283], stage0_51[284], stage0_51[285], stage0_51[286], stage0_51[287]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[53],stage1_53[76],stage1_52[126],stage1_51[177]}
   );
   gpc606_5 gpc2007 (
      {stage0_51[288], stage0_51[289], stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[54],stage1_53[77],stage1_52[127],stage1_51[178]}
   );
   gpc606_5 gpc2008 (
      {stage0_51[294], stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[55],stage1_53[78],stage1_52[128],stage1_51[179]}
   );
   gpc606_5 gpc2009 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304], stage0_51[305]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[56],stage1_53[79],stage1_52[129],stage1_51[180]}
   );
   gpc606_5 gpc2010 (
      {stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309], stage0_51[310], stage0_51[311]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[57],stage1_53[80],stage1_52[130],stage1_51[181]}
   );
   gpc606_5 gpc2011 (
      {stage0_51[312], stage0_51[313], stage0_51[314], stage0_51[315], stage0_51[316], stage0_51[317]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[58],stage1_53[81],stage1_52[131],stage1_51[182]}
   );
   gpc606_5 gpc2012 (
      {stage0_51[318], stage0_51[319], stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[59],stage1_53[82],stage1_52[132],stage1_51[183]}
   );
   gpc606_5 gpc2013 (
      {stage0_51[324], stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[60],stage1_53[83],stage1_52[133],stage1_51[184]}
   );
   gpc606_5 gpc2014 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334], stage0_51[335]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[61],stage1_53[84],stage1_52[134],stage1_51[185]}
   );
   gpc606_5 gpc2015 (
      {stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339], stage0_51[340], stage0_51[341]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[62],stage1_53[85],stage1_52[135],stage1_51[186]}
   );
   gpc606_5 gpc2016 (
      {stage0_51[342], stage0_51[343], stage0_51[344], stage0_51[345], stage0_51[346], stage0_51[347]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[63],stage1_53[86],stage1_52[136],stage1_51[187]}
   );
   gpc606_5 gpc2017 (
      {stage0_51[348], stage0_51[349], stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[64],stage1_53[87],stage1_52[137],stage1_51[188]}
   );
   gpc606_5 gpc2018 (
      {stage0_51[354], stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[65],stage1_53[88],stage1_52[138],stage1_51[189]}
   );
   gpc606_5 gpc2019 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364], stage0_51[365]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[66],stage1_53[89],stage1_52[139],stage1_51[190]}
   );
   gpc606_5 gpc2020 (
      {stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369], stage0_51[370], stage0_51[371]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[67],stage1_53[90],stage1_52[140],stage1_51[191]}
   );
   gpc606_5 gpc2021 (
      {stage0_51[372], stage0_51[373], stage0_51[374], stage0_51[375], stage0_51[376], stage0_51[377]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[68],stage1_53[91],stage1_52[141],stage1_51[192]}
   );
   gpc606_5 gpc2022 (
      {stage0_51[378], stage0_51[379], stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[69],stage1_53[92],stage1_52[142],stage1_51[193]}
   );
   gpc606_5 gpc2023 (
      {stage0_51[384], stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[70],stage1_53[93],stage1_52[143],stage1_51[194]}
   );
   gpc606_5 gpc2024 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394], stage0_51[395]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[71],stage1_53[94],stage1_52[144],stage1_51[195]}
   );
   gpc606_5 gpc2025 (
      {stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399], stage0_51[400], stage0_51[401]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[72],stage1_53[95],stage1_52[145],stage1_51[196]}
   );
   gpc606_5 gpc2026 (
      {stage0_51[402], stage0_51[403], stage0_51[404], stage0_51[405], stage0_51[406], stage0_51[407]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[73],stage1_53[96],stage1_52[146],stage1_51[197]}
   );
   gpc606_5 gpc2027 (
      {stage0_51[408], stage0_51[409], stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[74],stage1_53[97],stage1_52[147],stage1_51[198]}
   );
   gpc606_5 gpc2028 (
      {stage0_51[414], stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[75],stage1_53[98],stage1_52[148],stage1_51[199]}
   );
   gpc606_5 gpc2029 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424], stage0_51[425]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[76],stage1_53[99],stage1_52[149],stage1_51[200]}
   );
   gpc606_5 gpc2030 (
      {stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429], stage0_51[430], stage0_51[431]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[77],stage1_53[100],stage1_52[150],stage1_51[201]}
   );
   gpc606_5 gpc2031 (
      {stage0_51[432], stage0_51[433], stage0_51[434], stage0_51[435], stage0_51[436], stage0_51[437]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[78],stage1_53[101],stage1_52[151],stage1_51[202]}
   );
   gpc615_5 gpc2032 (
      {stage0_51[438], stage0_51[439], stage0_51[440], stage0_51[441], stage0_51[442]},
      {stage0_52[174]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[79],stage1_53[102],stage1_52[152],stage1_51[203]}
   );
   gpc615_5 gpc2033 (
      {stage0_51[443], stage0_51[444], stage0_51[445], stage0_51[446], stage0_51[447]},
      {stage0_52[175]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[80],stage1_53[103],stage1_52[153],stage1_51[204]}
   );
   gpc615_5 gpc2034 (
      {stage0_51[448], stage0_51[449], stage0_51[450], stage0_51[451], stage0_51[452]},
      {stage0_52[176]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[81],stage1_53[104],stage1_52[154],stage1_51[205]}
   );
   gpc615_5 gpc2035 (
      {stage0_51[453], stage0_51[454], stage0_51[455], stage0_51[456], stage0_51[457]},
      {stage0_52[177]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[82],stage1_53[105],stage1_52[155],stage1_51[206]}
   );
   gpc615_5 gpc2036 (
      {stage0_51[458], stage0_51[459], stage0_51[460], stage0_51[461], stage0_51[462]},
      {stage0_52[178]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[83],stage1_53[106],stage1_52[156],stage1_51[207]}
   );
   gpc615_5 gpc2037 (
      {stage0_51[463], stage0_51[464], stage0_51[465], stage0_51[466], stage0_51[467]},
      {stage0_52[179]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[84],stage1_53[107],stage1_52[157],stage1_51[208]}
   );
   gpc615_5 gpc2038 (
      {stage0_51[468], stage0_51[469], stage0_51[470], stage0_51[471], stage0_51[472]},
      {stage0_52[180]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[85],stage1_53[108],stage1_52[158],stage1_51[209]}
   );
   gpc615_5 gpc2039 (
      {stage0_51[473], stage0_51[474], stage0_51[475], stage0_51[476], stage0_51[477]},
      {stage0_52[181]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[86],stage1_53[109],stage1_52[159],stage1_51[210]}
   );
   gpc615_5 gpc2040 (
      {stage0_51[478], stage0_51[479], stage0_51[480], stage0_51[481], stage0_51[482]},
      {stage0_52[182]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[87],stage1_53[110],stage1_52[160],stage1_51[211]}
   );
   gpc615_5 gpc2041 (
      {stage0_51[483], stage0_51[484], stage0_51[485], stage0_51[486], stage0_51[487]},
      {stage0_52[183]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[88],stage1_53[111],stage1_52[161],stage1_51[212]}
   );
   gpc615_5 gpc2042 (
      {stage0_51[488], stage0_51[489], stage0_51[490], stage0_51[491], stage0_51[492]},
      {stage0_52[184]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[89],stage1_53[112],stage1_52[162],stage1_51[213]}
   );
   gpc615_5 gpc2043 (
      {stage0_51[493], stage0_51[494], stage0_51[495], stage0_51[496], stage0_51[497]},
      {stage0_52[185]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[90],stage1_53[113],stage1_52[163],stage1_51[214]}
   );
   gpc623_5 gpc2044 (
      {stage0_51[498], stage0_51[499], stage0_51[500]},
      {stage0_52[186], stage0_52[187]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[91],stage1_53[114],stage1_52[164],stage1_51[215]}
   );
   gpc606_5 gpc2045 (
      {stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191], stage0_52[192], stage0_52[193]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[92],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2046 (
      {stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197], stage0_52[198], stage0_52[199]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[93],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2047 (
      {stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203], stage0_52[204], stage0_52[205]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[94],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2048 (
      {stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209], stage0_52[210], stage0_52[211]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[95],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2049 (
      {stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215], stage0_52[216], stage0_52[217]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[96],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2050 (
      {stage0_52[218], stage0_52[219], stage0_52[220], stage0_52[221], stage0_52[222], stage0_52[223]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[97],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2051 (
      {stage0_52[224], stage0_52[225], stage0_52[226], stage0_52[227], stage0_52[228], stage0_52[229]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[98],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2052 (
      {stage0_52[230], stage0_52[231], stage0_52[232], stage0_52[233], stage0_52[234], stage0_52[235]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[99],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2053 (
      {stage0_52[236], stage0_52[237], stage0_52[238], stage0_52[239], stage0_52[240], stage0_52[241]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[100],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2054 (
      {stage0_52[242], stage0_52[243], stage0_52[244], stage0_52[245], stage0_52[246], stage0_52[247]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[101],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2055 (
      {stage0_52[248], stage0_52[249], stage0_52[250], stage0_52[251], stage0_52[252], stage0_52[253]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[102],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2056 (
      {stage0_52[254], stage0_52[255], stage0_52[256], stage0_52[257], stage0_52[258], stage0_52[259]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[103],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2057 (
      {stage0_52[260], stage0_52[261], stage0_52[262], stage0_52[263], stage0_52[264], stage0_52[265]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[104],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2058 (
      {stage0_52[266], stage0_52[267], stage0_52[268], stage0_52[269], stage0_52[270], stage0_52[271]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[105],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2059 (
      {stage0_52[272], stage0_52[273], stage0_52[274], stage0_52[275], stage0_52[276], stage0_52[277]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[106],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2060 (
      {stage0_52[278], stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[107],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2061 (
      {stage0_52[284], stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[108],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2062 (
      {stage0_52[290], stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[109],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2063 (
      {stage0_52[296], stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[110],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2064 (
      {stage0_52[302], stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[111],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2065 (
      {stage0_52[308], stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[112],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2066 (
      {stage0_52[314], stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[113],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2067 (
      {stage0_52[320], stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[114],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2068 (
      {stage0_52[326], stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[115],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2069 (
      {stage0_52[332], stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[116],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2070 (
      {stage0_52[338], stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[117],stage1_53[140],stage1_52[190]}
   );
   gpc606_5 gpc2071 (
      {stage0_52[344], stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[118],stage1_53[141],stage1_52[191]}
   );
   gpc606_5 gpc2072 (
      {stage0_52[350], stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[119],stage1_53[142],stage1_52[192]}
   );
   gpc606_5 gpc2073 (
      {stage0_52[356], stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[120],stage1_53[143],stage1_52[193]}
   );
   gpc606_5 gpc2074 (
      {stage0_52[362], stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[121],stage1_53[144],stage1_52[194]}
   );
   gpc606_5 gpc2075 (
      {stage0_52[368], stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[122],stage1_53[145],stage1_52[195]}
   );
   gpc606_5 gpc2076 (
      {stage0_52[374], stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[123],stage1_53[146],stage1_52[196]}
   );
   gpc606_5 gpc2077 (
      {stage0_52[380], stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[124],stage1_53[147],stage1_52[197]}
   );
   gpc606_5 gpc2078 (
      {stage0_52[386], stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[125],stage1_53[148],stage1_52[198]}
   );
   gpc606_5 gpc2079 (
      {stage0_52[392], stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[126],stage1_53[149],stage1_52[199]}
   );
   gpc606_5 gpc2080 (
      {stage0_52[398], stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[127],stage1_53[150],stage1_52[200]}
   );
   gpc606_5 gpc2081 (
      {stage0_52[404], stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409]},
      {stage0_54[216], stage0_54[217], stage0_54[218], stage0_54[219], stage0_54[220], stage0_54[221]},
      {stage1_56[36],stage1_55[99],stage1_54[128],stage1_53[151],stage1_52[201]}
   );
   gpc606_5 gpc2082 (
      {stage0_53[378], stage0_53[379], stage0_53[380], stage0_53[381], stage0_53[382], stage0_53[383]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[37],stage1_55[100],stage1_54[129],stage1_53[152]}
   );
   gpc606_5 gpc2083 (
      {stage0_53[384], stage0_53[385], stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[38],stage1_55[101],stage1_54[130],stage1_53[153]}
   );
   gpc606_5 gpc2084 (
      {stage0_53[390], stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[39],stage1_55[102],stage1_54[131],stage1_53[154]}
   );
   gpc606_5 gpc2085 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400], stage0_53[401]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[40],stage1_55[103],stage1_54[132],stage1_53[155]}
   );
   gpc606_5 gpc2086 (
      {stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405], stage0_53[406], stage0_53[407]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[41],stage1_55[104],stage1_54[133],stage1_53[156]}
   );
   gpc606_5 gpc2087 (
      {stage0_53[408], stage0_53[409], stage0_53[410], stage0_53[411], stage0_53[412], stage0_53[413]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[42],stage1_55[105],stage1_54[134],stage1_53[157]}
   );
   gpc606_5 gpc2088 (
      {stage0_53[414], stage0_53[415], stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[43],stage1_55[106],stage1_54[135],stage1_53[158]}
   );
   gpc606_5 gpc2089 (
      {stage0_53[420], stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[44],stage1_55[107],stage1_54[136],stage1_53[159]}
   );
   gpc606_5 gpc2090 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430], stage0_53[431]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[45],stage1_55[108],stage1_54[137],stage1_53[160]}
   );
   gpc606_5 gpc2091 (
      {stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435], stage0_53[436], stage0_53[437]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[46],stage1_55[109],stage1_54[138],stage1_53[161]}
   );
   gpc606_5 gpc2092 (
      {stage0_53[438], stage0_53[439], stage0_53[440], stage0_53[441], stage0_53[442], stage0_53[443]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[47],stage1_55[110],stage1_54[139],stage1_53[162]}
   );
   gpc606_5 gpc2093 (
      {stage0_53[444], stage0_53[445], stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[48],stage1_55[111],stage1_54[140],stage1_53[163]}
   );
   gpc606_5 gpc2094 (
      {stage0_53[450], stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[49],stage1_55[112],stage1_54[141],stage1_53[164]}
   );
   gpc606_5 gpc2095 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460], stage0_53[461]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[50],stage1_55[113],stage1_54[142],stage1_53[165]}
   );
   gpc606_5 gpc2096 (
      {stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465], stage0_53[466], stage0_53[467]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[51],stage1_55[114],stage1_54[143],stage1_53[166]}
   );
   gpc606_5 gpc2097 (
      {stage0_53[468], stage0_53[469], stage0_53[470], stage0_53[471], stage0_53[472], stage0_53[473]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[52],stage1_55[115],stage1_54[144],stage1_53[167]}
   );
   gpc606_5 gpc2098 (
      {stage0_53[474], stage0_53[475], stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[53],stage1_55[116],stage1_54[145],stage1_53[168]}
   );
   gpc606_5 gpc2099 (
      {stage0_53[480], stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[54],stage1_55[117],stage1_54[146],stage1_53[169]}
   );
   gpc606_5 gpc2100 (
      {stage0_53[486], stage0_53[487], stage0_53[488], stage0_53[489], stage0_53[490], stage0_53[491]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[55],stage1_55[118],stage1_54[147],stage1_53[170]}
   );
   gpc615_5 gpc2101 (
      {stage0_53[492], stage0_53[493], stage0_53[494], stage0_53[495], stage0_53[496]},
      {stage0_54[222]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[56],stage1_55[119],stage1_54[148],stage1_53[171]}
   );
   gpc606_5 gpc2102 (
      {stage0_54[223], stage0_54[224], stage0_54[225], stage0_54[226], stage0_54[227], stage0_54[228]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[20],stage1_56[57],stage1_55[120],stage1_54[149]}
   );
   gpc606_5 gpc2103 (
      {stage0_54[229], stage0_54[230], stage0_54[231], stage0_54[232], stage0_54[233], stage0_54[234]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[21],stage1_56[58],stage1_55[121],stage1_54[150]}
   );
   gpc606_5 gpc2104 (
      {stage0_54[235], stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[22],stage1_56[59],stage1_55[122],stage1_54[151]}
   );
   gpc615_5 gpc2105 (
      {stage0_54[241], stage0_54[242], stage0_54[243], stage0_54[244], stage0_54[245]},
      {stage0_55[120]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[23],stage1_56[60],stage1_55[123],stage1_54[152]}
   );
   gpc615_5 gpc2106 (
      {stage0_54[246], stage0_54[247], stage0_54[248], stage0_54[249], stage0_54[250]},
      {stage0_55[121]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[24],stage1_56[61],stage1_55[124],stage1_54[153]}
   );
   gpc615_5 gpc2107 (
      {stage0_54[251], stage0_54[252], stage0_54[253], stage0_54[254], stage0_54[255]},
      {stage0_55[122]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[25],stage1_56[62],stage1_55[125],stage1_54[154]}
   );
   gpc615_5 gpc2108 (
      {stage0_54[256], stage0_54[257], stage0_54[258], stage0_54[259], stage0_54[260]},
      {stage0_55[123]},
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage1_58[6],stage1_57[26],stage1_56[63],stage1_55[126],stage1_54[155]}
   );
   gpc615_5 gpc2109 (
      {stage0_54[261], stage0_54[262], stage0_54[263], stage0_54[264], stage0_54[265]},
      {stage0_55[124]},
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage1_58[7],stage1_57[27],stage1_56[64],stage1_55[127],stage1_54[156]}
   );
   gpc615_5 gpc2110 (
      {stage0_54[266], stage0_54[267], stage0_54[268], stage0_54[269], stage0_54[270]},
      {stage0_55[125]},
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage1_58[8],stage1_57[28],stage1_56[65],stage1_55[128],stage1_54[157]}
   );
   gpc615_5 gpc2111 (
      {stage0_54[271], stage0_54[272], stage0_54[273], stage0_54[274], stage0_54[275]},
      {stage0_55[126]},
      {stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59]},
      {stage1_58[9],stage1_57[29],stage1_56[66],stage1_55[129],stage1_54[158]}
   );
   gpc615_5 gpc2112 (
      {stage0_54[276], stage0_54[277], stage0_54[278], stage0_54[279], stage0_54[280]},
      {stage0_55[127]},
      {stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65]},
      {stage1_58[10],stage1_57[30],stage1_56[67],stage1_55[130],stage1_54[159]}
   );
   gpc615_5 gpc2113 (
      {stage0_54[281], stage0_54[282], stage0_54[283], stage0_54[284], stage0_54[285]},
      {stage0_55[128]},
      {stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71]},
      {stage1_58[11],stage1_57[31],stage1_56[68],stage1_55[131],stage1_54[160]}
   );
   gpc615_5 gpc2114 (
      {stage0_54[286], stage0_54[287], stage0_54[288], stage0_54[289], stage0_54[290]},
      {stage0_55[129]},
      {stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77]},
      {stage1_58[12],stage1_57[32],stage1_56[69],stage1_55[132],stage1_54[161]}
   );
   gpc615_5 gpc2115 (
      {stage0_54[291], stage0_54[292], stage0_54[293], stage0_54[294], stage0_54[295]},
      {stage0_55[130]},
      {stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83]},
      {stage1_58[13],stage1_57[33],stage1_56[70],stage1_55[133],stage1_54[162]}
   );
   gpc615_5 gpc2116 (
      {stage0_54[296], stage0_54[297], stage0_54[298], stage0_54[299], stage0_54[300]},
      {stage0_55[131]},
      {stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89]},
      {stage1_58[14],stage1_57[34],stage1_56[71],stage1_55[134],stage1_54[163]}
   );
   gpc615_5 gpc2117 (
      {stage0_54[301], stage0_54[302], stage0_54[303], stage0_54[304], stage0_54[305]},
      {stage0_55[132]},
      {stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95]},
      {stage1_58[15],stage1_57[35],stage1_56[72],stage1_55[135],stage1_54[164]}
   );
   gpc615_5 gpc2118 (
      {stage0_54[306], stage0_54[307], stage0_54[308], stage0_54[309], stage0_54[310]},
      {stage0_55[133]},
      {stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101]},
      {stage1_58[16],stage1_57[36],stage1_56[73],stage1_55[136],stage1_54[165]}
   );
   gpc615_5 gpc2119 (
      {stage0_54[311], stage0_54[312], stage0_54[313], stage0_54[314], stage0_54[315]},
      {stage0_55[134]},
      {stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107]},
      {stage1_58[17],stage1_57[37],stage1_56[74],stage1_55[137],stage1_54[166]}
   );
   gpc615_5 gpc2120 (
      {stage0_54[316], stage0_54[317], stage0_54[318], stage0_54[319], stage0_54[320]},
      {stage0_55[135]},
      {stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113]},
      {stage1_58[18],stage1_57[38],stage1_56[75],stage1_55[138],stage1_54[167]}
   );
   gpc615_5 gpc2121 (
      {stage0_54[321], stage0_54[322], stage0_54[323], stage0_54[324], stage0_54[325]},
      {stage0_55[136]},
      {stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119]},
      {stage1_58[19],stage1_57[39],stage1_56[76],stage1_55[139],stage1_54[168]}
   );
   gpc615_5 gpc2122 (
      {stage0_54[326], stage0_54[327], stage0_54[328], stage0_54[329], stage0_54[330]},
      {stage0_55[137]},
      {stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125]},
      {stage1_58[20],stage1_57[40],stage1_56[77],stage1_55[140],stage1_54[169]}
   );
   gpc615_5 gpc2123 (
      {stage0_54[331], stage0_54[332], stage0_54[333], stage0_54[334], stage0_54[335]},
      {stage0_55[138]},
      {stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131]},
      {stage1_58[21],stage1_57[41],stage1_56[78],stage1_55[141],stage1_54[170]}
   );
   gpc615_5 gpc2124 (
      {stage0_54[336], stage0_54[337], stage0_54[338], stage0_54[339], stage0_54[340]},
      {stage0_55[139]},
      {stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137]},
      {stage1_58[22],stage1_57[42],stage1_56[79],stage1_55[142],stage1_54[171]}
   );
   gpc615_5 gpc2125 (
      {stage0_54[341], stage0_54[342], stage0_54[343], stage0_54[344], stage0_54[345]},
      {stage0_55[140]},
      {stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143]},
      {stage1_58[23],stage1_57[43],stage1_56[80],stage1_55[143],stage1_54[172]}
   );
   gpc615_5 gpc2126 (
      {stage0_54[346], stage0_54[347], stage0_54[348], stage0_54[349], stage0_54[350]},
      {stage0_55[141]},
      {stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149]},
      {stage1_58[24],stage1_57[44],stage1_56[81],stage1_55[144],stage1_54[173]}
   );
   gpc615_5 gpc2127 (
      {stage0_54[351], stage0_54[352], stage0_54[353], stage0_54[354], stage0_54[355]},
      {stage0_55[142]},
      {stage0_56[150], stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155]},
      {stage1_58[25],stage1_57[45],stage1_56[82],stage1_55[145],stage1_54[174]}
   );
   gpc615_5 gpc2128 (
      {stage0_54[356], stage0_54[357], stage0_54[358], stage0_54[359], stage0_54[360]},
      {stage0_55[143]},
      {stage0_56[156], stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161]},
      {stage1_58[26],stage1_57[46],stage1_56[83],stage1_55[146],stage1_54[175]}
   );
   gpc615_5 gpc2129 (
      {stage0_54[361], stage0_54[362], stage0_54[363], stage0_54[364], stage0_54[365]},
      {stage0_55[144]},
      {stage0_56[162], stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167]},
      {stage1_58[27],stage1_57[47],stage1_56[84],stage1_55[147],stage1_54[176]}
   );
   gpc615_5 gpc2130 (
      {stage0_54[366], stage0_54[367], stage0_54[368], stage0_54[369], stage0_54[370]},
      {stage0_55[145]},
      {stage0_56[168], stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173]},
      {stage1_58[28],stage1_57[48],stage1_56[85],stage1_55[148],stage1_54[177]}
   );
   gpc615_5 gpc2131 (
      {stage0_54[371], stage0_54[372], stage0_54[373], stage0_54[374], stage0_54[375]},
      {stage0_55[146]},
      {stage0_56[174], stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179]},
      {stage1_58[29],stage1_57[49],stage1_56[86],stage1_55[149],stage1_54[178]}
   );
   gpc615_5 gpc2132 (
      {stage0_54[376], stage0_54[377], stage0_54[378], stage0_54[379], stage0_54[380]},
      {stage0_55[147]},
      {stage0_56[180], stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185]},
      {stage1_58[30],stage1_57[50],stage1_56[87],stage1_55[150],stage1_54[179]}
   );
   gpc615_5 gpc2133 (
      {stage0_54[381], stage0_54[382], stage0_54[383], stage0_54[384], stage0_54[385]},
      {stage0_55[148]},
      {stage0_56[186], stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191]},
      {stage1_58[31],stage1_57[51],stage1_56[88],stage1_55[151],stage1_54[180]}
   );
   gpc615_5 gpc2134 (
      {stage0_54[386], stage0_54[387], stage0_54[388], stage0_54[389], stage0_54[390]},
      {stage0_55[149]},
      {stage0_56[192], stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197]},
      {stage1_58[32],stage1_57[52],stage1_56[89],stage1_55[152],stage1_54[181]}
   );
   gpc615_5 gpc2135 (
      {stage0_54[391], stage0_54[392], stage0_54[393], stage0_54[394], stage0_54[395]},
      {stage0_55[150]},
      {stage0_56[198], stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203]},
      {stage1_58[33],stage1_57[53],stage1_56[90],stage1_55[153],stage1_54[182]}
   );
   gpc615_5 gpc2136 (
      {stage0_54[396], stage0_54[397], stage0_54[398], stage0_54[399], stage0_54[400]},
      {stage0_55[151]},
      {stage0_56[204], stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209]},
      {stage1_58[34],stage1_57[54],stage1_56[91],stage1_55[154],stage1_54[183]}
   );
   gpc615_5 gpc2137 (
      {stage0_54[401], stage0_54[402], stage0_54[403], stage0_54[404], stage0_54[405]},
      {stage0_55[152]},
      {stage0_56[210], stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215]},
      {stage1_58[35],stage1_57[55],stage1_56[92],stage1_55[155],stage1_54[184]}
   );
   gpc615_5 gpc2138 (
      {stage0_54[406], stage0_54[407], stage0_54[408], stage0_54[409], stage0_54[410]},
      {stage0_55[153]},
      {stage0_56[216], stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221]},
      {stage1_58[36],stage1_57[56],stage1_56[93],stage1_55[156],stage1_54[185]}
   );
   gpc615_5 gpc2139 (
      {stage0_54[411], stage0_54[412], stage0_54[413], stage0_54[414], stage0_54[415]},
      {stage0_55[154]},
      {stage0_56[222], stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227]},
      {stage1_58[37],stage1_57[57],stage1_56[94],stage1_55[157],stage1_54[186]}
   );
   gpc615_5 gpc2140 (
      {stage0_54[416], stage0_54[417], stage0_54[418], stage0_54[419], stage0_54[420]},
      {stage0_55[155]},
      {stage0_56[228], stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233]},
      {stage1_58[38],stage1_57[58],stage1_56[95],stage1_55[158],stage1_54[187]}
   );
   gpc615_5 gpc2141 (
      {stage0_54[421], stage0_54[422], stage0_54[423], stage0_54[424], stage0_54[425]},
      {stage0_55[156]},
      {stage0_56[234], stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239]},
      {stage1_58[39],stage1_57[59],stage1_56[96],stage1_55[159],stage1_54[188]}
   );
   gpc615_5 gpc2142 (
      {stage0_54[426], stage0_54[427], stage0_54[428], stage0_54[429], stage0_54[430]},
      {stage0_55[157]},
      {stage0_56[240], stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245]},
      {stage1_58[40],stage1_57[60],stage1_56[97],stage1_55[160],stage1_54[189]}
   );
   gpc615_5 gpc2143 (
      {stage0_54[431], stage0_54[432], stage0_54[433], stage0_54[434], stage0_54[435]},
      {stage0_55[158]},
      {stage0_56[246], stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251]},
      {stage1_58[41],stage1_57[61],stage1_56[98],stage1_55[161],stage1_54[190]}
   );
   gpc615_5 gpc2144 (
      {stage0_54[436], stage0_54[437], stage0_54[438], stage0_54[439], stage0_54[440]},
      {stage0_55[159]},
      {stage0_56[252], stage0_56[253], stage0_56[254], stage0_56[255], stage0_56[256], stage0_56[257]},
      {stage1_58[42],stage1_57[62],stage1_56[99],stage1_55[162],stage1_54[191]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[160], stage0_55[161], stage0_55[162], stage0_55[163], stage0_55[164], stage0_55[165]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[43],stage1_57[63],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[166], stage0_55[167], stage0_55[168], stage0_55[169], stage0_55[170], stage0_55[171]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[44],stage1_57[64],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2147 (
      {stage0_55[172], stage0_55[173], stage0_55[174], stage0_55[175], stage0_55[176], stage0_55[177]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[45],stage1_57[65],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2148 (
      {stage0_55[178], stage0_55[179], stage0_55[180], stage0_55[181], stage0_55[182], stage0_55[183]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[46],stage1_57[66],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2149 (
      {stage0_55[184], stage0_55[185], stage0_55[186], stage0_55[187], stage0_55[188], stage0_55[189]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[47],stage1_57[67],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2150 (
      {stage0_55[190], stage0_55[191], stage0_55[192], stage0_55[193], stage0_55[194], stage0_55[195]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[48],stage1_57[68],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2151 (
      {stage0_55[196], stage0_55[197], stage0_55[198], stage0_55[199], stage0_55[200], stage0_55[201]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[49],stage1_57[69],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2152 (
      {stage0_55[202], stage0_55[203], stage0_55[204], stage0_55[205], stage0_55[206], stage0_55[207]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[50],stage1_57[70],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2153 (
      {stage0_55[208], stage0_55[209], stage0_55[210], stage0_55[211], stage0_55[212], stage0_55[213]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[51],stage1_57[71],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2154 (
      {stage0_55[214], stage0_55[215], stage0_55[216], stage0_55[217], stage0_55[218], stage0_55[219]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[52],stage1_57[72],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2155 (
      {stage0_55[220], stage0_55[221], stage0_55[222], stage0_55[223], stage0_55[224], stage0_55[225]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[53],stage1_57[73],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2156 (
      {stage0_55[226], stage0_55[227], stage0_55[228], stage0_55[229], stage0_55[230], stage0_55[231]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[54],stage1_57[74],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2157 (
      {stage0_55[232], stage0_55[233], stage0_55[234], stage0_55[235], stage0_55[236], stage0_55[237]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[55],stage1_57[75],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2158 (
      {stage0_55[238], stage0_55[239], stage0_55[240], stage0_55[241], stage0_55[242], stage0_55[243]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[56],stage1_57[76],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2159 (
      {stage0_55[244], stage0_55[245], stage0_55[246], stage0_55[247], stage0_55[248], stage0_55[249]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[57],stage1_57[77],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2160 (
      {stage0_55[250], stage0_55[251], stage0_55[252], stage0_55[253], stage0_55[254], stage0_55[255]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[58],stage1_57[78],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2161 (
      {stage0_55[256], stage0_55[257], stage0_55[258], stage0_55[259], stage0_55[260], stage0_55[261]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[59],stage1_57[79],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2162 (
      {stage0_55[262], stage0_55[263], stage0_55[264], stage0_55[265], stage0_55[266], stage0_55[267]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[60],stage1_57[80],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2163 (
      {stage0_55[268], stage0_55[269], stage0_55[270], stage0_55[271], stage0_55[272], stage0_55[273]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[61],stage1_57[81],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2164 (
      {stage0_55[274], stage0_55[275], stage0_55[276], stage0_55[277], stage0_55[278], stage0_55[279]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[62],stage1_57[82],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2165 (
      {stage0_55[280], stage0_55[281], stage0_55[282], stage0_55[283], stage0_55[284], stage0_55[285]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[63],stage1_57[83],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2166 (
      {stage0_55[286], stage0_55[287], stage0_55[288], stage0_55[289], stage0_55[290], stage0_55[291]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[64],stage1_57[84],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2167 (
      {stage0_55[292], stage0_55[293], stage0_55[294], stage0_55[295], stage0_55[296], stage0_55[297]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[65],stage1_57[85],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2168 (
      {stage0_55[298], stage0_55[299], stage0_55[300], stage0_55[301], stage0_55[302], stage0_55[303]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[66],stage1_57[86],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2169 (
      {stage0_55[304], stage0_55[305], stage0_55[306], stage0_55[307], stage0_55[308], stage0_55[309]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[67],stage1_57[87],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2170 (
      {stage0_55[310], stage0_55[311], stage0_55[312], stage0_55[313], stage0_55[314], stage0_55[315]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[68],stage1_57[88],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2171 (
      {stage0_55[316], stage0_55[317], stage0_55[318], stage0_55[319], stage0_55[320], stage0_55[321]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[69],stage1_57[89],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2172 (
      {stage0_55[322], stage0_55[323], stage0_55[324], stage0_55[325], stage0_55[326], stage0_55[327]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[70],stage1_57[90],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2173 (
      {stage0_55[328], stage0_55[329], stage0_55[330], stage0_55[331], stage0_55[332], stage0_55[333]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[71],stage1_57[91],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2174 (
      {stage0_55[334], stage0_55[335], stage0_55[336], stage0_55[337], stage0_55[338], stage0_55[339]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[72],stage1_57[92],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2175 (
      {stage0_55[340], stage0_55[341], stage0_55[342], stage0_55[343], stage0_55[344], stage0_55[345]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[73],stage1_57[93],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2176 (
      {stage0_55[346], stage0_55[347], stage0_55[348], stage0_55[349], stage0_55[350], stage0_55[351]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[74],stage1_57[94],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2177 (
      {stage0_55[352], stage0_55[353], stage0_55[354], stage0_55[355], stage0_55[356], stage0_55[357]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[75],stage1_57[95],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2178 (
      {stage0_55[358], stage0_55[359], stage0_55[360], stage0_55[361], stage0_55[362], stage0_55[363]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[76],stage1_57[96],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2179 (
      {stage0_55[364], stage0_55[365], stage0_55[366], stage0_55[367], stage0_55[368], stage0_55[369]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[77],stage1_57[97],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2180 (
      {stage0_55[370], stage0_55[371], stage0_55[372], stage0_55[373], stage0_55[374], stage0_55[375]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[78],stage1_57[98],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2181 (
      {stage0_55[376], stage0_55[377], stage0_55[378], stage0_55[379], stage0_55[380], stage0_55[381]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[79],stage1_57[99],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2182 (
      {stage0_55[382], stage0_55[383], stage0_55[384], stage0_55[385], stage0_55[386], stage0_55[387]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[80],stage1_57[100],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2183 (
      {stage0_55[388], stage0_55[389], stage0_55[390], stage0_55[391], stage0_55[392], stage0_55[393]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[81],stage1_57[101],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2184 (
      {stage0_55[394], stage0_55[395], stage0_55[396], stage0_55[397], stage0_55[398], stage0_55[399]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[82],stage1_57[102],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2185 (
      {stage0_55[400], stage0_55[401], stage0_55[402], stage0_55[403], stage0_55[404], stage0_55[405]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[83],stage1_57[103],stage1_56[140],stage1_55[203]}
   );
   gpc606_5 gpc2186 (
      {stage0_55[406], stage0_55[407], stage0_55[408], stage0_55[409], stage0_55[410], stage0_55[411]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[84],stage1_57[104],stage1_56[141],stage1_55[204]}
   );
   gpc606_5 gpc2187 (
      {stage0_55[412], stage0_55[413], stage0_55[414], stage0_55[415], stage0_55[416], stage0_55[417]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[85],stage1_57[105],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2188 (
      {stage0_55[418], stage0_55[419], stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[86],stage1_57[106],stage1_56[143],stage1_55[206]}
   );
   gpc606_5 gpc2189 (
      {stage0_55[424], stage0_55[425], stage0_55[426], stage0_55[427], stage0_55[428], stage0_55[429]},
      {stage0_57[264], stage0_57[265], stage0_57[266], stage0_57[267], stage0_57[268], stage0_57[269]},
      {stage1_59[44],stage1_58[87],stage1_57[107],stage1_56[144],stage1_55[207]}
   );
   gpc606_5 gpc2190 (
      {stage0_55[430], stage0_55[431], stage0_55[432], stage0_55[433], stage0_55[434], stage0_55[435]},
      {stage0_57[270], stage0_57[271], stage0_57[272], stage0_57[273], stage0_57[274], stage0_57[275]},
      {stage1_59[45],stage1_58[88],stage1_57[108],stage1_56[145],stage1_55[208]}
   );
   gpc606_5 gpc2191 (
      {stage0_55[436], stage0_55[437], stage0_55[438], stage0_55[439], stage0_55[440], stage0_55[441]},
      {stage0_57[276], stage0_57[277], stage0_57[278], stage0_57[279], stage0_57[280], stage0_57[281]},
      {stage1_59[46],stage1_58[89],stage1_57[109],stage1_56[146],stage1_55[209]}
   );
   gpc606_5 gpc2192 (
      {stage0_55[442], stage0_55[443], stage0_55[444], stage0_55[445], stage0_55[446], stage0_55[447]},
      {stage0_57[282], stage0_57[283], stage0_57[284], stage0_57[285], stage0_57[286], stage0_57[287]},
      {stage1_59[47],stage1_58[90],stage1_57[110],stage1_56[147],stage1_55[210]}
   );
   gpc606_5 gpc2193 (
      {stage0_55[448], stage0_55[449], stage0_55[450], stage0_55[451], stage0_55[452], stage0_55[453]},
      {stage0_57[288], stage0_57[289], stage0_57[290], stage0_57[291], stage0_57[292], stage0_57[293]},
      {stage1_59[48],stage1_58[91],stage1_57[111],stage1_56[148],stage1_55[211]}
   );
   gpc606_5 gpc2194 (
      {stage0_55[454], stage0_55[455], stage0_55[456], stage0_55[457], stage0_55[458], stage0_55[459]},
      {stage0_57[294], stage0_57[295], stage0_57[296], stage0_57[297], stage0_57[298], stage0_57[299]},
      {stage1_59[49],stage1_58[92],stage1_57[112],stage1_56[149],stage1_55[212]}
   );
   gpc606_5 gpc2195 (
      {stage0_55[460], stage0_55[461], stage0_55[462], stage0_55[463], stage0_55[464], stage0_55[465]},
      {stage0_57[300], stage0_57[301], stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305]},
      {stage1_59[50],stage1_58[93],stage1_57[113],stage1_56[150],stage1_55[213]}
   );
   gpc606_5 gpc2196 (
      {stage0_55[466], stage0_55[467], stage0_55[468], stage0_55[469], stage0_55[470], stage0_55[471]},
      {stage0_57[306], stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage1_59[51],stage1_58[94],stage1_57[114],stage1_56[151],stage1_55[214]}
   );
   gpc606_5 gpc2197 (
      {stage0_55[472], stage0_55[473], stage0_55[474], stage0_55[475], stage0_55[476], stage0_55[477]},
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316], stage0_57[317]},
      {stage1_59[52],stage1_58[95],stage1_57[115],stage1_56[152],stage1_55[215]}
   );
   gpc615_5 gpc2198 (
      {stage0_55[478], stage0_55[479], stage0_55[480], stage0_55[481], stage0_55[482]},
      {stage0_56[258]},
      {stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321], stage0_57[322], stage0_57[323]},
      {stage1_59[53],stage1_58[96],stage1_57[116],stage1_56[153],stage1_55[216]}
   );
   gpc615_5 gpc2199 (
      {stage0_55[483], stage0_55[484], stage0_55[485], stage0_55[486], stage0_55[487]},
      {stage0_56[259]},
      {stage0_57[324], stage0_57[325], stage0_57[326], stage0_57[327], stage0_57[328], stage0_57[329]},
      {stage1_59[54],stage1_58[97],stage1_57[117],stage1_56[154],stage1_55[217]}
   );
   gpc615_5 gpc2200 (
      {stage0_55[488], stage0_55[489], stage0_55[490], stage0_55[491], stage0_55[492]},
      {stage0_56[260]},
      {stage0_57[330], stage0_57[331], stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335]},
      {stage1_59[55],stage1_58[98],stage1_57[118],stage1_56[155],stage1_55[218]}
   );
   gpc615_5 gpc2201 (
      {stage0_55[493], stage0_55[494], stage0_55[495], stage0_55[496], stage0_55[497]},
      {stage0_56[261]},
      {stage0_57[336], stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage1_59[56],stage1_58[99],stage1_57[119],stage1_56[156],stage1_55[219]}
   );
   gpc615_5 gpc2202 (
      {stage0_55[498], stage0_55[499], stage0_55[500], stage0_55[501], stage0_55[502]},
      {stage0_56[262]},
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346], stage0_57[347]},
      {stage1_59[57],stage1_58[100],stage1_57[120],stage1_56[157],stage1_55[220]}
   );
   gpc615_5 gpc2203 (
      {stage0_55[503], stage0_55[504], stage0_55[505], stage0_55[506], stage0_55[507]},
      {stage0_56[263]},
      {stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351], stage0_57[352], stage0_57[353]},
      {stage1_59[58],stage1_58[101],stage1_57[121],stage1_56[158],stage1_55[221]}
   );
   gpc606_5 gpc2204 (
      {stage0_56[264], stage0_56[265], stage0_56[266], stage0_56[267], stage0_56[268], stage0_56[269]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[59],stage1_58[102],stage1_57[122],stage1_56[159]}
   );
   gpc606_5 gpc2205 (
      {stage0_56[270], stage0_56[271], stage0_56[272], stage0_56[273], stage0_56[274], stage0_56[275]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[60],stage1_58[103],stage1_57[123],stage1_56[160]}
   );
   gpc606_5 gpc2206 (
      {stage0_56[276], stage0_56[277], stage0_56[278], stage0_56[279], stage0_56[280], stage0_56[281]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[61],stage1_58[104],stage1_57[124],stage1_56[161]}
   );
   gpc606_5 gpc2207 (
      {stage0_56[282], stage0_56[283], stage0_56[284], stage0_56[285], stage0_56[286], stage0_56[287]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[62],stage1_58[105],stage1_57[125],stage1_56[162]}
   );
   gpc606_5 gpc2208 (
      {stage0_56[288], stage0_56[289], stage0_56[290], stage0_56[291], stage0_56[292], stage0_56[293]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[63],stage1_58[106],stage1_57[126],stage1_56[163]}
   );
   gpc606_5 gpc2209 (
      {stage0_56[294], stage0_56[295], stage0_56[296], stage0_56[297], stage0_56[298], stage0_56[299]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[64],stage1_58[107],stage1_57[127],stage1_56[164]}
   );
   gpc606_5 gpc2210 (
      {stage0_56[300], stage0_56[301], stage0_56[302], stage0_56[303], stage0_56[304], stage0_56[305]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[65],stage1_58[108],stage1_57[128],stage1_56[165]}
   );
   gpc606_5 gpc2211 (
      {stage0_56[306], stage0_56[307], stage0_56[308], stage0_56[309], stage0_56[310], stage0_56[311]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[66],stage1_58[109],stage1_57[129],stage1_56[166]}
   );
   gpc606_5 gpc2212 (
      {stage0_56[312], stage0_56[313], stage0_56[314], stage0_56[315], stage0_56[316], stage0_56[317]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[67],stage1_58[110],stage1_57[130],stage1_56[167]}
   );
   gpc606_5 gpc2213 (
      {stage0_56[318], stage0_56[319], stage0_56[320], stage0_56[321], stage0_56[322], stage0_56[323]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[68],stage1_58[111],stage1_57[131],stage1_56[168]}
   );
   gpc606_5 gpc2214 (
      {stage0_56[324], stage0_56[325], stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[69],stage1_58[112],stage1_57[132],stage1_56[169]}
   );
   gpc606_5 gpc2215 (
      {stage0_56[330], stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[70],stage1_58[113],stage1_57[133],stage1_56[170]}
   );
   gpc606_5 gpc2216 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340], stage0_56[341]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[71],stage1_58[114],stage1_57[134],stage1_56[171]}
   );
   gpc606_5 gpc2217 (
      {stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345], stage0_56[346], stage0_56[347]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[72],stage1_58[115],stage1_57[135],stage1_56[172]}
   );
   gpc606_5 gpc2218 (
      {stage0_56[348], stage0_56[349], stage0_56[350], stage0_56[351], stage0_56[352], stage0_56[353]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[73],stage1_58[116],stage1_57[136],stage1_56[173]}
   );
   gpc606_5 gpc2219 (
      {stage0_56[354], stage0_56[355], stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[74],stage1_58[117],stage1_57[137],stage1_56[174]}
   );
   gpc606_5 gpc2220 (
      {stage0_56[360], stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[75],stage1_58[118],stage1_57[138],stage1_56[175]}
   );
   gpc606_5 gpc2221 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370], stage0_56[371]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[76],stage1_58[119],stage1_57[139],stage1_56[176]}
   );
   gpc606_5 gpc2222 (
      {stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375], stage0_56[376], stage0_56[377]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[77],stage1_58[120],stage1_57[140],stage1_56[177]}
   );
   gpc606_5 gpc2223 (
      {stage0_56[378], stage0_56[379], stage0_56[380], stage0_56[381], stage0_56[382], stage0_56[383]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[78],stage1_58[121],stage1_57[141],stage1_56[178]}
   );
   gpc606_5 gpc2224 (
      {stage0_56[384], stage0_56[385], stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[79],stage1_58[122],stage1_57[142],stage1_56[179]}
   );
   gpc606_5 gpc2225 (
      {stage0_56[390], stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[80],stage1_58[123],stage1_57[143],stage1_56[180]}
   );
   gpc606_5 gpc2226 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400], stage0_56[401]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[81],stage1_58[124],stage1_57[144],stage1_56[181]}
   );
   gpc606_5 gpc2227 (
      {stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405], stage0_56[406], stage0_56[407]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[82],stage1_58[125],stage1_57[145],stage1_56[182]}
   );
   gpc606_5 gpc2228 (
      {stage0_56[408], stage0_56[409], stage0_56[410], stage0_56[411], stage0_56[412], stage0_56[413]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[83],stage1_58[126],stage1_57[146],stage1_56[183]}
   );
   gpc606_5 gpc2229 (
      {stage0_56[414], stage0_56[415], stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[84],stage1_58[127],stage1_57[147],stage1_56[184]}
   );
   gpc606_5 gpc2230 (
      {stage0_56[420], stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[85],stage1_58[128],stage1_57[148],stage1_56[185]}
   );
   gpc606_5 gpc2231 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430], stage0_56[431]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[86],stage1_58[129],stage1_57[149],stage1_56[186]}
   );
   gpc606_5 gpc2232 (
      {stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435], stage0_56[436], stage0_56[437]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[87],stage1_58[130],stage1_57[150],stage1_56[187]}
   );
   gpc606_5 gpc2233 (
      {stage0_56[438], stage0_56[439], stage0_56[440], stage0_56[441], stage0_56[442], stage0_56[443]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[88],stage1_58[131],stage1_57[151],stage1_56[188]}
   );
   gpc606_5 gpc2234 (
      {stage0_57[354], stage0_57[355], stage0_57[356], stage0_57[357], stage0_57[358], stage0_57[359]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[30],stage1_59[89],stage1_58[132],stage1_57[152]}
   );
   gpc606_5 gpc2235 (
      {stage0_57[360], stage0_57[361], stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[31],stage1_59[90],stage1_58[133],stage1_57[153]}
   );
   gpc606_5 gpc2236 (
      {stage0_57[366], stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[32],stage1_59[91],stage1_58[134],stage1_57[154]}
   );
   gpc606_5 gpc2237 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376], stage0_57[377]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[33],stage1_59[92],stage1_58[135],stage1_57[155]}
   );
   gpc606_5 gpc2238 (
      {stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381], stage0_57[382], stage0_57[383]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[34],stage1_59[93],stage1_58[136],stage1_57[156]}
   );
   gpc606_5 gpc2239 (
      {stage0_57[384], stage0_57[385], stage0_57[386], stage0_57[387], stage0_57[388], stage0_57[389]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[35],stage1_59[94],stage1_58[137],stage1_57[157]}
   );
   gpc606_5 gpc2240 (
      {stage0_57[390], stage0_57[391], stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[36],stage1_59[95],stage1_58[138],stage1_57[158]}
   );
   gpc606_5 gpc2241 (
      {stage0_57[396], stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[37],stage1_59[96],stage1_58[139],stage1_57[159]}
   );
   gpc606_5 gpc2242 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406], stage0_57[407]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[38],stage1_59[97],stage1_58[140],stage1_57[160]}
   );
   gpc606_5 gpc2243 (
      {stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411], stage0_57[412], stage0_57[413]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[39],stage1_59[98],stage1_58[141],stage1_57[161]}
   );
   gpc606_5 gpc2244 (
      {stage0_57[414], stage0_57[415], stage0_57[416], stage0_57[417], stage0_57[418], stage0_57[419]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[40],stage1_59[99],stage1_58[142],stage1_57[162]}
   );
   gpc606_5 gpc2245 (
      {stage0_57[420], stage0_57[421], stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[41],stage1_59[100],stage1_58[143],stage1_57[163]}
   );
   gpc606_5 gpc2246 (
      {stage0_57[426], stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[42],stage1_59[101],stage1_58[144],stage1_57[164]}
   );
   gpc606_5 gpc2247 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436], stage0_57[437]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[43],stage1_59[102],stage1_58[145],stage1_57[165]}
   );
   gpc606_5 gpc2248 (
      {stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441], stage0_57[442], stage0_57[443]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[44],stage1_59[103],stage1_58[146],stage1_57[166]}
   );
   gpc606_5 gpc2249 (
      {stage0_57[444], stage0_57[445], stage0_57[446], stage0_57[447], stage0_57[448], stage0_57[449]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[45],stage1_59[104],stage1_58[147],stage1_57[167]}
   );
   gpc606_5 gpc2250 (
      {stage0_57[450], stage0_57[451], stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[46],stage1_59[105],stage1_58[148],stage1_57[168]}
   );
   gpc606_5 gpc2251 (
      {stage0_57[456], stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[47],stage1_59[106],stage1_58[149],stage1_57[169]}
   );
   gpc606_5 gpc2252 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466], stage0_57[467]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[48],stage1_59[107],stage1_58[150],stage1_57[170]}
   );
   gpc606_5 gpc2253 (
      {stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471], stage0_57[472], stage0_57[473]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[49],stage1_59[108],stage1_58[151],stage1_57[171]}
   );
   gpc606_5 gpc2254 (
      {stage0_57[474], stage0_57[475], stage0_57[476], stage0_57[477], stage0_57[478], stage0_57[479]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[50],stage1_59[109],stage1_58[152],stage1_57[172]}
   );
   gpc606_5 gpc2255 (
      {stage0_57[480], stage0_57[481], stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[51],stage1_59[110],stage1_58[153],stage1_57[173]}
   );
   gpc606_5 gpc2256 (
      {stage0_57[486], stage0_57[487], stage0_57[488], stage0_57[489], stage0_57[490], stage0_57[491]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[52],stage1_59[111],stage1_58[154],stage1_57[174]}
   );
   gpc606_5 gpc2257 (
      {stage0_57[492], stage0_57[493], stage0_57[494], stage0_57[495], stage0_57[496], stage0_57[497]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[53],stage1_59[112],stage1_58[155],stage1_57[175]}
   );
   gpc606_5 gpc2258 (
      {stage0_57[498], stage0_57[499], stage0_57[500], stage0_57[501], stage0_57[502], stage0_57[503]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[54],stage1_59[113],stage1_58[156],stage1_57[176]}
   );
   gpc606_5 gpc2259 (
      {stage0_57[504], stage0_57[505], stage0_57[506], stage0_57[507], stage0_57[508], stage0_57[509]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[55],stage1_59[114],stage1_58[157],stage1_57[177]}
   );
   gpc2135_5 gpc2260 (
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184]},
      {stage0_59[156], stage0_59[157], stage0_59[158]},
      {stage0_60[0]},
      {stage0_61[0], stage0_61[1]},
      {stage1_62[0],stage1_61[26],stage1_60[56],stage1_59[115],stage1_58[158]}
   );
   gpc2135_5 gpc2261 (
      {stage0_58[185], stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189]},
      {stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage0_60[1]},
      {stage0_61[2], stage0_61[3]},
      {stage1_62[1],stage1_61[27],stage1_60[57],stage1_59[116],stage1_58[159]}
   );
   gpc2135_5 gpc2262 (
      {stage0_58[190], stage0_58[191], stage0_58[192], stage0_58[193], stage0_58[194]},
      {stage0_59[162], stage0_59[163], stage0_59[164]},
      {stage0_60[2]},
      {stage0_61[4], stage0_61[5]},
      {stage1_62[2],stage1_61[28],stage1_60[58],stage1_59[117],stage1_58[160]}
   );
   gpc2135_5 gpc2263 (
      {stage0_58[195], stage0_58[196], stage0_58[197], stage0_58[198], stage0_58[199]},
      {stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage0_60[3]},
      {stage0_61[6], stage0_61[7]},
      {stage1_62[3],stage1_61[29],stage1_60[59],stage1_59[118],stage1_58[161]}
   );
   gpc2135_5 gpc2264 (
      {stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203], stage0_58[204]},
      {stage0_59[168], stage0_59[169], stage0_59[170]},
      {stage0_60[4]},
      {stage0_61[8], stage0_61[9]},
      {stage1_62[4],stage1_61[30],stage1_60[60],stage1_59[119],stage1_58[162]}
   );
   gpc2135_5 gpc2265 (
      {stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage0_60[5]},
      {stage0_61[10], stage0_61[11]},
      {stage1_62[5],stage1_61[31],stage1_60[61],stage1_59[120],stage1_58[163]}
   );
   gpc2135_5 gpc2266 (
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214]},
      {stage0_59[174], stage0_59[175], stage0_59[176]},
      {stage0_60[6]},
      {stage0_61[12], stage0_61[13]},
      {stage1_62[6],stage1_61[32],stage1_60[62],stage1_59[121],stage1_58[164]}
   );
   gpc2135_5 gpc2267 (
      {stage0_58[215], stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219]},
      {stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage0_60[7]},
      {stage0_61[14], stage0_61[15]},
      {stage1_62[7],stage1_61[33],stage1_60[63],stage1_59[122],stage1_58[165]}
   );
   gpc2135_5 gpc2268 (
      {stage0_58[220], stage0_58[221], stage0_58[222], stage0_58[223], stage0_58[224]},
      {stage0_59[180], stage0_59[181], stage0_59[182]},
      {stage0_60[8]},
      {stage0_61[16], stage0_61[17]},
      {stage1_62[8],stage1_61[34],stage1_60[64],stage1_59[123],stage1_58[166]}
   );
   gpc2135_5 gpc2269 (
      {stage0_58[225], stage0_58[226], stage0_58[227], stage0_58[228], stage0_58[229]},
      {stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage0_60[9]},
      {stage0_61[18], stage0_61[19]},
      {stage1_62[9],stage1_61[35],stage1_60[65],stage1_59[124],stage1_58[167]}
   );
   gpc2135_5 gpc2270 (
      {stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233], stage0_58[234]},
      {stage0_59[186], stage0_59[187], stage0_59[188]},
      {stage0_60[10]},
      {stage0_61[20], stage0_61[21]},
      {stage1_62[10],stage1_61[36],stage1_60[66],stage1_59[125],stage1_58[168]}
   );
   gpc2135_5 gpc2271 (
      {stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage0_60[11]},
      {stage0_61[22], stage0_61[23]},
      {stage1_62[11],stage1_61[37],stage1_60[67],stage1_59[126],stage1_58[169]}
   );
   gpc2135_5 gpc2272 (
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244]},
      {stage0_59[192], stage0_59[193], stage0_59[194]},
      {stage0_60[12]},
      {stage0_61[24], stage0_61[25]},
      {stage1_62[12],stage1_61[38],stage1_60[68],stage1_59[127],stage1_58[170]}
   );
   gpc2135_5 gpc2273 (
      {stage0_58[245], stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249]},
      {stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage0_60[13]},
      {stage0_61[26], stage0_61[27]},
      {stage1_62[13],stage1_61[39],stage1_60[69],stage1_59[128],stage1_58[171]}
   );
   gpc2135_5 gpc2274 (
      {stage0_58[250], stage0_58[251], stage0_58[252], stage0_58[253], stage0_58[254]},
      {stage0_59[198], stage0_59[199], stage0_59[200]},
      {stage0_60[14]},
      {stage0_61[28], stage0_61[29]},
      {stage1_62[14],stage1_61[40],stage1_60[70],stage1_59[129],stage1_58[172]}
   );
   gpc2135_5 gpc2275 (
      {stage0_58[255], stage0_58[256], stage0_58[257], stage0_58[258], stage0_58[259]},
      {stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage0_60[15]},
      {stage0_61[30], stage0_61[31]},
      {stage1_62[15],stage1_61[41],stage1_60[71],stage1_59[130],stage1_58[173]}
   );
   gpc1163_5 gpc2276 (
      {stage0_58[260], stage0_58[261], stage0_58[262]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage0_60[16]},
      {stage0_61[32]},
      {stage1_62[16],stage1_61[42],stage1_60[72],stage1_59[131],stage1_58[174]}
   );
   gpc1163_5 gpc2277 (
      {stage0_58[263], stage0_58[264], stage0_58[265]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage0_60[17]},
      {stage0_61[33]},
      {stage1_62[17],stage1_61[43],stage1_60[73],stage1_59[132],stage1_58[175]}
   );
   gpc1163_5 gpc2278 (
      {stage0_58[266], stage0_58[267], stage0_58[268]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage0_60[18]},
      {stage0_61[34]},
      {stage1_62[18],stage1_61[44],stage1_60[74],stage1_59[133],stage1_58[176]}
   );
   gpc1163_5 gpc2279 (
      {stage0_58[269], stage0_58[270], stage0_58[271]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage0_60[19]},
      {stage0_61[35]},
      {stage1_62[19],stage1_61[45],stage1_60[75],stage1_59[134],stage1_58[177]}
   );
   gpc1163_5 gpc2280 (
      {stage0_58[272], stage0_58[273], stage0_58[274]},
      {stage0_59[228], stage0_59[229], stage0_59[230], stage0_59[231], stage0_59[232], stage0_59[233]},
      {stage0_60[20]},
      {stage0_61[36]},
      {stage1_62[20],stage1_61[46],stage1_60[76],stage1_59[135],stage1_58[178]}
   );
   gpc1163_5 gpc2281 (
      {stage0_58[275], stage0_58[276], stage0_58[277]},
      {stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238], stage0_59[239]},
      {stage0_60[21]},
      {stage0_61[37]},
      {stage1_62[21],stage1_61[47],stage1_60[77],stage1_59[136],stage1_58[179]}
   );
   gpc1163_5 gpc2282 (
      {stage0_58[278], stage0_58[279], stage0_58[280]},
      {stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[22]},
      {stage0_61[38]},
      {stage1_62[22],stage1_61[48],stage1_60[78],stage1_59[137],stage1_58[180]}
   );
   gpc1163_5 gpc2283 (
      {stage0_58[281], stage0_58[282], stage0_58[283]},
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251]},
      {stage0_60[23]},
      {stage0_61[39]},
      {stage1_62[23],stage1_61[49],stage1_60[79],stage1_59[138],stage1_58[181]}
   );
   gpc1163_5 gpc2284 (
      {stage0_58[284], stage0_58[285], stage0_58[286]},
      {stage0_59[252], stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257]},
      {stage0_60[24]},
      {stage0_61[40]},
      {stage1_62[24],stage1_61[50],stage1_60[80],stage1_59[139],stage1_58[182]}
   );
   gpc1163_5 gpc2285 (
      {stage0_58[287], stage0_58[288], stage0_58[289]},
      {stage0_59[258], stage0_59[259], stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263]},
      {stage0_60[25]},
      {stage0_61[41]},
      {stage1_62[25],stage1_61[51],stage1_60[81],stage1_59[140],stage1_58[183]}
   );
   gpc1163_5 gpc2286 (
      {stage0_58[290], stage0_58[291], stage0_58[292]},
      {stage0_59[264], stage0_59[265], stage0_59[266], stage0_59[267], stage0_59[268], stage0_59[269]},
      {stage0_60[26]},
      {stage0_61[42]},
      {stage1_62[26],stage1_61[52],stage1_60[82],stage1_59[141],stage1_58[184]}
   );
   gpc1163_5 gpc2287 (
      {stage0_58[293], stage0_58[294], stage0_58[295]},
      {stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273], stage0_59[274], stage0_59[275]},
      {stage0_60[27]},
      {stage0_61[43]},
      {stage1_62[27],stage1_61[53],stage1_60[83],stage1_59[142],stage1_58[185]}
   );
   gpc1163_5 gpc2288 (
      {stage0_58[296], stage0_58[297], stage0_58[298]},
      {stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280], stage0_59[281]},
      {stage0_60[28]},
      {stage0_61[44]},
      {stage1_62[28],stage1_61[54],stage1_60[84],stage1_59[143],stage1_58[186]}
   );
   gpc1163_5 gpc2289 (
      {stage0_58[299], stage0_58[300], stage0_58[301]},
      {stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[29]},
      {stage0_61[45]},
      {stage1_62[29],stage1_61[55],stage1_60[85],stage1_59[144],stage1_58[187]}
   );
   gpc1163_5 gpc2290 (
      {stage0_58[302], stage0_58[303], stage0_58[304]},
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293]},
      {stage0_60[30]},
      {stage0_61[46]},
      {stage1_62[30],stage1_61[56],stage1_60[86],stage1_59[145],stage1_58[188]}
   );
   gpc1163_5 gpc2291 (
      {stage0_58[305], stage0_58[306], stage0_58[307]},
      {stage0_59[294], stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299]},
      {stage0_60[31]},
      {stage0_61[47]},
      {stage1_62[31],stage1_61[57],stage1_60[87],stage1_59[146],stage1_58[189]}
   );
   gpc1163_5 gpc2292 (
      {stage0_58[308], stage0_58[309], stage0_58[310]},
      {stage0_59[300], stage0_59[301], stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305]},
      {stage0_60[32]},
      {stage0_61[48]},
      {stage1_62[32],stage1_61[58],stage1_60[88],stage1_59[147],stage1_58[190]}
   );
   gpc1163_5 gpc2293 (
      {stage0_58[311], stage0_58[312], stage0_58[313]},
      {stage0_59[306], stage0_59[307], stage0_59[308], stage0_59[309], stage0_59[310], stage0_59[311]},
      {stage0_60[33]},
      {stage0_61[49]},
      {stage1_62[33],stage1_61[59],stage1_60[89],stage1_59[148],stage1_58[191]}
   );
   gpc1163_5 gpc2294 (
      {stage0_58[314], stage0_58[315], stage0_58[316]},
      {stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315], stage0_59[316], stage0_59[317]},
      {stage0_60[34]},
      {stage0_61[50]},
      {stage1_62[34],stage1_61[60],stage1_60[90],stage1_59[149],stage1_58[192]}
   );
   gpc1163_5 gpc2295 (
      {stage0_58[317], stage0_58[318], stage0_58[319]},
      {stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322], stage0_59[323]},
      {stage0_60[35]},
      {stage0_61[51]},
      {stage1_62[35],stage1_61[61],stage1_60[91],stage1_59[150],stage1_58[193]}
   );
   gpc1163_5 gpc2296 (
      {stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[36]},
      {stage0_61[52]},
      {stage1_62[36],stage1_61[62],stage1_60[92],stage1_59[151],stage1_58[194]}
   );
   gpc606_5 gpc2297 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328]},
      {stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41], stage0_60[42]},
      {stage1_62[37],stage1_61[63],stage1_60[93],stage1_59[152],stage1_58[195]}
   );
   gpc606_5 gpc2298 (
      {stage0_58[329], stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334]},
      {stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47], stage0_60[48]},
      {stage1_62[38],stage1_61[64],stage1_60[94],stage1_59[153],stage1_58[196]}
   );
   gpc606_5 gpc2299 (
      {stage0_58[335], stage0_58[336], stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340]},
      {stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53], stage0_60[54]},
      {stage1_62[39],stage1_61[65],stage1_60[95],stage1_59[154],stage1_58[197]}
   );
   gpc606_5 gpc2300 (
      {stage0_58[341], stage0_58[342], stage0_58[343], stage0_58[344], stage0_58[345], stage0_58[346]},
      {stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59], stage0_60[60]},
      {stage1_62[40],stage1_61[66],stage1_60[96],stage1_59[155],stage1_58[198]}
   );
   gpc606_5 gpc2301 (
      {stage0_58[347], stage0_58[348], stage0_58[349], stage0_58[350], stage0_58[351], stage0_58[352]},
      {stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65], stage0_60[66]},
      {stage1_62[41],stage1_61[67],stage1_60[97],stage1_59[156],stage1_58[199]}
   );
   gpc606_5 gpc2302 (
      {stage0_58[353], stage0_58[354], stage0_58[355], stage0_58[356], stage0_58[357], stage0_58[358]},
      {stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71], stage0_60[72]},
      {stage1_62[42],stage1_61[68],stage1_60[98],stage1_59[157],stage1_58[200]}
   );
   gpc606_5 gpc2303 (
      {stage0_58[359], stage0_58[360], stage0_58[361], stage0_58[362], stage0_58[363], stage0_58[364]},
      {stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77], stage0_60[78]},
      {stage1_62[43],stage1_61[69],stage1_60[99],stage1_59[158],stage1_58[201]}
   );
   gpc606_5 gpc2304 (
      {stage0_58[365], stage0_58[366], stage0_58[367], stage0_58[368], stage0_58[369], stage0_58[370]},
      {stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83], stage0_60[84]},
      {stage1_62[44],stage1_61[70],stage1_60[100],stage1_59[159],stage1_58[202]}
   );
   gpc606_5 gpc2305 (
      {stage0_58[371], stage0_58[372], stage0_58[373], stage0_58[374], stage0_58[375], stage0_58[376]},
      {stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89], stage0_60[90]},
      {stage1_62[45],stage1_61[71],stage1_60[101],stage1_59[160],stage1_58[203]}
   );
   gpc606_5 gpc2306 (
      {stage0_58[377], stage0_58[378], stage0_58[379], stage0_58[380], stage0_58[381], stage0_58[382]},
      {stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95], stage0_60[96]},
      {stage1_62[46],stage1_61[72],stage1_60[102],stage1_59[161],stage1_58[204]}
   );
   gpc606_5 gpc2307 (
      {stage0_58[383], stage0_58[384], stage0_58[385], stage0_58[386], stage0_58[387], stage0_58[388]},
      {stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101], stage0_60[102]},
      {stage1_62[47],stage1_61[73],stage1_60[103],stage1_59[162],stage1_58[205]}
   );
   gpc606_5 gpc2308 (
      {stage0_58[389], stage0_58[390], stage0_58[391], stage0_58[392], stage0_58[393], stage0_58[394]},
      {stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107], stage0_60[108]},
      {stage1_62[48],stage1_61[74],stage1_60[104],stage1_59[163],stage1_58[206]}
   );
   gpc606_5 gpc2309 (
      {stage0_58[395], stage0_58[396], stage0_58[397], stage0_58[398], stage0_58[399], stage0_58[400]},
      {stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113], stage0_60[114]},
      {stage1_62[49],stage1_61[75],stage1_60[105],stage1_59[164],stage1_58[207]}
   );
   gpc606_5 gpc2310 (
      {stage0_58[401], stage0_58[402], stage0_58[403], stage0_58[404], stage0_58[405], stage0_58[406]},
      {stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119], stage0_60[120]},
      {stage1_62[50],stage1_61[76],stage1_60[106],stage1_59[165],stage1_58[208]}
   );
   gpc606_5 gpc2311 (
      {stage0_58[407], stage0_58[408], stage0_58[409], stage0_58[410], stage0_58[411], stage0_58[412]},
      {stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125], stage0_60[126]},
      {stage1_62[51],stage1_61[77],stage1_60[107],stage1_59[166],stage1_58[209]}
   );
   gpc606_5 gpc2312 (
      {stage0_58[413], stage0_58[414], stage0_58[415], stage0_58[416], stage0_58[417], stage0_58[418]},
      {stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131], stage0_60[132]},
      {stage1_62[52],stage1_61[78],stage1_60[108],stage1_59[167],stage1_58[210]}
   );
   gpc606_5 gpc2313 (
      {stage0_58[419], stage0_58[420], stage0_58[421], stage0_58[422], stage0_58[423], stage0_58[424]},
      {stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138]},
      {stage1_62[53],stage1_61[79],stage1_60[109],stage1_59[168],stage1_58[211]}
   );
   gpc606_5 gpc2314 (
      {stage0_58[425], stage0_58[426], stage0_58[427], stage0_58[428], stage0_58[429], stage0_58[430]},
      {stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144]},
      {stage1_62[54],stage1_61[80],stage1_60[110],stage1_59[169],stage1_58[212]}
   );
   gpc606_5 gpc2315 (
      {stage0_58[431], stage0_58[432], stage0_58[433], stage0_58[434], stage0_58[435], stage0_58[436]},
      {stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage1_62[55],stage1_61[81],stage1_60[111],stage1_59[170],stage1_58[213]}
   );
   gpc606_5 gpc2316 (
      {stage0_58[437], stage0_58[438], stage0_58[439], stage0_58[440], stage0_58[441], stage0_58[442]},
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155], stage0_60[156]},
      {stage1_62[56],stage1_61[82],stage1_60[112],stage1_59[171],stage1_58[214]}
   );
   gpc606_5 gpc2317 (
      {stage0_58[443], stage0_58[444], stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448]},
      {stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161], stage0_60[162]},
      {stage1_62[57],stage1_61[83],stage1_60[113],stage1_59[172],stage1_58[215]}
   );
   gpc606_5 gpc2318 (
      {stage0_58[449], stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_60[163], stage0_60[164], stage0_60[165], stage0_60[166], stage0_60[167], stage0_60[168]},
      {stage1_62[58],stage1_61[84],stage1_60[114],stage1_59[173],stage1_58[216]}
   );
   gpc606_5 gpc2319 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459], stage0_58[460]},
      {stage0_60[169], stage0_60[170], stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174]},
      {stage1_62[59],stage1_61[85],stage1_60[115],stage1_59[174],stage1_58[217]}
   );
   gpc606_5 gpc2320 (
      {stage0_58[461], stage0_58[462], stage0_58[463], stage0_58[464], stage0_58[465], stage0_58[466]},
      {stage0_60[175], stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage1_62[60],stage1_61[86],stage1_60[116],stage1_59[175],stage1_58[218]}
   );
   gpc606_5 gpc2321 (
      {stage0_58[467], stage0_58[468], stage0_58[469], stage0_58[470], stage0_58[471], stage0_58[472]},
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185], stage0_60[186]},
      {stage1_62[61],stage1_61[87],stage1_60[117],stage1_59[176],stage1_58[219]}
   );
   gpc615_5 gpc2322 (
      {stage0_58[473], stage0_58[474], stage0_58[475], stage0_58[476], stage0_58[477]},
      {stage0_59[330]},
      {stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190], stage0_60[191], stage0_60[192]},
      {stage1_62[62],stage1_61[88],stage1_60[118],stage1_59[177],stage1_58[220]}
   );
   gpc615_5 gpc2323 (
      {stage0_58[478], stage0_58[479], stage0_58[480], stage0_58[481], stage0_58[482]},
      {stage0_59[331]},
      {stage0_60[193], stage0_60[194], stage0_60[195], stage0_60[196], stage0_60[197], stage0_60[198]},
      {stage1_62[63],stage1_61[89],stage1_60[119],stage1_59[178],stage1_58[221]}
   );
   gpc615_5 gpc2324 (
      {stage0_58[483], stage0_58[484], stage0_58[485], stage0_58[486], stage0_58[487]},
      {stage0_59[332]},
      {stage0_60[199], stage0_60[200], stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204]},
      {stage1_62[64],stage1_61[90],stage1_60[120],stage1_59[179],stage1_58[222]}
   );
   gpc615_5 gpc2325 (
      {stage0_58[488], stage0_58[489], stage0_58[490], stage0_58[491], stage0_58[492]},
      {stage0_59[333]},
      {stage0_60[205], stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage1_62[65],stage1_61[91],stage1_60[121],stage1_59[180],stage1_58[223]}
   );
   gpc606_5 gpc2326 (
      {stage0_59[334], stage0_59[335], stage0_59[336], stage0_59[337], stage0_59[338], stage0_59[339]},
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58]},
      {stage1_63[0],stage1_62[66],stage1_61[92],stage1_60[122],stage1_59[181]}
   );
   gpc606_5 gpc2327 (
      {stage0_59[340], stage0_59[341], stage0_59[342], stage0_59[343], stage0_59[344], stage0_59[345]},
      {stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64]},
      {stage1_63[1],stage1_62[67],stage1_61[93],stage1_60[123],stage1_59[182]}
   );
   gpc606_5 gpc2328 (
      {stage0_59[346], stage0_59[347], stage0_59[348], stage0_59[349], stage0_59[350], stage0_59[351]},
      {stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70]},
      {stage1_63[2],stage1_62[68],stage1_61[94],stage1_60[124],stage1_59[183]}
   );
   gpc606_5 gpc2329 (
      {stage0_59[352], stage0_59[353], stage0_59[354], stage0_59[355], stage0_59[356], stage0_59[357]},
      {stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76]},
      {stage1_63[3],stage1_62[69],stage1_61[95],stage1_60[125],stage1_59[184]}
   );
   gpc606_5 gpc2330 (
      {stage0_59[358], stage0_59[359], stage0_59[360], stage0_59[361], stage0_59[362], stage0_59[363]},
      {stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82]},
      {stage1_63[4],stage1_62[70],stage1_61[96],stage1_60[126],stage1_59[185]}
   );
   gpc606_5 gpc2331 (
      {stage0_59[364], stage0_59[365], stage0_59[366], stage0_59[367], stage0_59[368], stage0_59[369]},
      {stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88]},
      {stage1_63[5],stage1_62[71],stage1_61[97],stage1_60[127],stage1_59[186]}
   );
   gpc606_5 gpc2332 (
      {stage0_59[370], stage0_59[371], stage0_59[372], stage0_59[373], stage0_59[374], stage0_59[375]},
      {stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94]},
      {stage1_63[6],stage1_62[72],stage1_61[98],stage1_60[128],stage1_59[187]}
   );
   gpc606_5 gpc2333 (
      {stage0_59[376], stage0_59[377], stage0_59[378], stage0_59[379], stage0_59[380], stage0_59[381]},
      {stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100]},
      {stage1_63[7],stage1_62[73],stage1_61[99],stage1_60[129],stage1_59[188]}
   );
   gpc606_5 gpc2334 (
      {stage0_59[382], stage0_59[383], stage0_59[384], stage0_59[385], stage0_59[386], stage0_59[387]},
      {stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106]},
      {stage1_63[8],stage1_62[74],stage1_61[100],stage1_60[130],stage1_59[189]}
   );
   gpc606_5 gpc2335 (
      {stage0_59[388], stage0_59[389], stage0_59[390], stage0_59[391], stage0_59[392], stage0_59[393]},
      {stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112]},
      {stage1_63[9],stage1_62[75],stage1_61[101],stage1_60[131],stage1_59[190]}
   );
   gpc606_5 gpc2336 (
      {stage0_59[394], stage0_59[395], stage0_59[396], stage0_59[397], stage0_59[398], stage0_59[399]},
      {stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118]},
      {stage1_63[10],stage1_62[76],stage1_61[102],stage1_60[132],stage1_59[191]}
   );
   gpc606_5 gpc2337 (
      {stage0_59[400], stage0_59[401], stage0_59[402], stage0_59[403], stage0_59[404], stage0_59[405]},
      {stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124]},
      {stage1_63[11],stage1_62[77],stage1_61[103],stage1_60[133],stage1_59[192]}
   );
   gpc606_5 gpc2338 (
      {stage0_59[406], stage0_59[407], stage0_59[408], stage0_59[409], stage0_59[410], stage0_59[411]},
      {stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130]},
      {stage1_63[12],stage1_62[78],stage1_61[104],stage1_60[134],stage1_59[193]}
   );
   gpc606_5 gpc2339 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215], stage0_60[216]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[13],stage1_62[79],stage1_61[105],stage1_60[135]}
   );
   gpc606_5 gpc2340 (
      {stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220], stage0_60[221], stage0_60[222]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[14],stage1_62[80],stage1_61[106],stage1_60[136]}
   );
   gpc606_5 gpc2341 (
      {stage0_60[223], stage0_60[224], stage0_60[225], stage0_60[226], stage0_60[227], stage0_60[228]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[15],stage1_62[81],stage1_61[107],stage1_60[137]}
   );
   gpc606_5 gpc2342 (
      {stage0_60[229], stage0_60[230], stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[16],stage1_62[82],stage1_61[108],stage1_60[138]}
   );
   gpc606_5 gpc2343 (
      {stage0_60[235], stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[17],stage1_62[83],stage1_61[109],stage1_60[139]}
   );
   gpc606_5 gpc2344 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245], stage0_60[246]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[18],stage1_62[84],stage1_61[110],stage1_60[140]}
   );
   gpc606_5 gpc2345 (
      {stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250], stage0_60[251], stage0_60[252]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[19],stage1_62[85],stage1_61[111],stage1_60[141]}
   );
   gpc606_5 gpc2346 (
      {stage0_60[253], stage0_60[254], stage0_60[255], stage0_60[256], stage0_60[257], stage0_60[258]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[20],stage1_62[86],stage1_61[112],stage1_60[142]}
   );
   gpc606_5 gpc2347 (
      {stage0_60[259], stage0_60[260], stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[21],stage1_62[87],stage1_61[113],stage1_60[143]}
   );
   gpc606_5 gpc2348 (
      {stage0_60[265], stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[22],stage1_62[88],stage1_61[114],stage1_60[144]}
   );
   gpc606_5 gpc2349 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275], stage0_60[276]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[23],stage1_62[89],stage1_61[115],stage1_60[145]}
   );
   gpc606_5 gpc2350 (
      {stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280], stage0_60[281], stage0_60[282]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[24],stage1_62[90],stage1_61[116],stage1_60[146]}
   );
   gpc606_5 gpc2351 (
      {stage0_60[283], stage0_60[284], stage0_60[285], stage0_60[286], stage0_60[287], stage0_60[288]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[25],stage1_62[91],stage1_61[117],stage1_60[147]}
   );
   gpc606_5 gpc2352 (
      {stage0_60[289], stage0_60[290], stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[26],stage1_62[92],stage1_61[118],stage1_60[148]}
   );
   gpc606_5 gpc2353 (
      {stage0_60[295], stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[27],stage1_62[93],stage1_61[119],stage1_60[149]}
   );
   gpc606_5 gpc2354 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305], stage0_60[306]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[28],stage1_62[94],stage1_61[120],stage1_60[150]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310], stage0_60[311]},
      {stage0_61[131]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[29],stage1_62[95],stage1_61[121],stage1_60[151]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315], stage0_60[316]},
      {stage0_61[132]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[30],stage1_62[96],stage1_61[122],stage1_60[152]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320], stage0_60[321]},
      {stage0_61[133]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[31],stage1_62[97],stage1_61[123],stage1_60[153]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325], stage0_60[326]},
      {stage0_61[134]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[32],stage1_62[98],stage1_61[124],stage1_60[154]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330], stage0_60[331]},
      {stage0_61[135]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[33],stage1_62[99],stage1_61[125],stage1_60[155]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335], stage0_60[336]},
      {stage0_61[136]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[34],stage1_62[100],stage1_61[126],stage1_60[156]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340], stage0_60[341]},
      {stage0_61[137]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[35],stage1_62[101],stage1_61[127],stage1_60[157]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345], stage0_60[346]},
      {stage0_61[138]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[36],stage1_62[102],stage1_61[128],stage1_60[158]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350], stage0_60[351]},
      {stage0_61[139]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[37],stage1_62[103],stage1_61[129],stage1_60[159]}
   );
   gpc615_5 gpc2364 (
      {stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355], stage0_60[356]},
      {stage0_61[140]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[38],stage1_62[104],stage1_61[130],stage1_60[160]}
   );
   gpc615_5 gpc2365 (
      {stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360], stage0_60[361]},
      {stage0_61[141]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[39],stage1_62[105],stage1_61[131],stage1_60[161]}
   );
   gpc615_5 gpc2366 (
      {stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365], stage0_60[366]},
      {stage0_61[142]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[40],stage1_62[106],stage1_61[132],stage1_60[162]}
   );
   gpc615_5 gpc2367 (
      {stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370], stage0_60[371]},
      {stage0_61[143]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[41],stage1_62[107],stage1_61[133],stage1_60[163]}
   );
   gpc615_5 gpc2368 (
      {stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375], stage0_60[376]},
      {stage0_61[144]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[42],stage1_62[108],stage1_61[134],stage1_60[164]}
   );
   gpc615_5 gpc2369 (
      {stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380], stage0_60[381]},
      {stage0_61[145]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[43],stage1_62[109],stage1_61[135],stage1_60[165]}
   );
   gpc615_5 gpc2370 (
      {stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385], stage0_60[386]},
      {stage0_61[146]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[44],stage1_62[110],stage1_61[136],stage1_60[166]}
   );
   gpc615_5 gpc2371 (
      {stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390], stage0_60[391]},
      {stage0_61[147]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[45],stage1_62[111],stage1_61[137],stage1_60[167]}
   );
   gpc615_5 gpc2372 (
      {stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395], stage0_60[396]},
      {stage0_61[148]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[46],stage1_62[112],stage1_61[138],stage1_60[168]}
   );
   gpc615_5 gpc2373 (
      {stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400], stage0_60[401]},
      {stage0_61[149]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[47],stage1_62[113],stage1_61[139],stage1_60[169]}
   );
   gpc615_5 gpc2374 (
      {stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405], stage0_60[406]},
      {stage0_61[150]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[48],stage1_62[114],stage1_61[140],stage1_60[170]}
   );
   gpc615_5 gpc2375 (
      {stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410], stage0_60[411]},
      {stage0_61[151]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[49],stage1_62[115],stage1_61[141],stage1_60[171]}
   );
   gpc615_5 gpc2376 (
      {stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415], stage0_60[416]},
      {stage0_61[152]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[50],stage1_62[116],stage1_61[142],stage1_60[172]}
   );
   gpc615_5 gpc2377 (
      {stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420], stage0_60[421]},
      {stage0_61[153]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[51],stage1_62[117],stage1_61[143],stage1_60[173]}
   );
   gpc615_5 gpc2378 (
      {stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425], stage0_60[426]},
      {stage0_61[154]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[52],stage1_62[118],stage1_61[144],stage1_60[174]}
   );
   gpc615_5 gpc2379 (
      {stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430], stage0_60[431]},
      {stage0_61[155]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[53],stage1_62[119],stage1_61[145],stage1_60[175]}
   );
   gpc615_5 gpc2380 (
      {stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435], stage0_60[436]},
      {stage0_61[156]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[54],stage1_62[120],stage1_61[146],stage1_60[176]}
   );
   gpc615_5 gpc2381 (
      {stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440], stage0_60[441]},
      {stage0_61[157]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[55],stage1_62[121],stage1_61[147],stage1_60[177]}
   );
   gpc615_5 gpc2382 (
      {stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445], stage0_60[446]},
      {stage0_61[158]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[56],stage1_62[122],stage1_61[148],stage1_60[178]}
   );
   gpc615_5 gpc2383 (
      {stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450], stage0_60[451]},
      {stage0_61[159]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[57],stage1_62[123],stage1_61[149],stage1_60[179]}
   );
   gpc615_5 gpc2384 (
      {stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455], stage0_60[456]},
      {stage0_61[160]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[58],stage1_62[124],stage1_61[150],stage1_60[180]}
   );
   gpc615_5 gpc2385 (
      {stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460], stage0_60[461]},
      {stage0_61[161]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[59],stage1_62[125],stage1_61[151],stage1_60[181]}
   );
   gpc615_5 gpc2386 (
      {stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465], stage0_60[466]},
      {stage0_61[162]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[60],stage1_62[126],stage1_61[152],stage1_60[182]}
   );
   gpc615_5 gpc2387 (
      {stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470], stage0_60[471]},
      {stage0_61[163]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[61],stage1_62[127],stage1_61[153],stage1_60[183]}
   );
   gpc615_5 gpc2388 (
      {stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475], stage0_60[476]},
      {stage0_61[164]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[62],stage1_62[128],stage1_61[154],stage1_60[184]}
   );
   gpc615_5 gpc2389 (
      {stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480], stage0_60[481]},
      {stage0_61[165]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[63],stage1_62[129],stage1_61[155],stage1_60[185]}
   );
   gpc615_5 gpc2390 (
      {stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485], stage0_60[486]},
      {stage0_61[166]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[64],stage1_62[130],stage1_61[156],stage1_60[186]}
   );
   gpc615_5 gpc2391 (
      {stage0_60[487], stage0_60[488], stage0_60[489], stage0_60[490], stage0_60[491]},
      {stage0_61[167]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[65],stage1_62[131],stage1_61[157],stage1_60[187]}
   );
   gpc615_5 gpc2392 (
      {stage0_60[492], stage0_60[493], stage0_60[494], stage0_60[495], stage0_60[496]},
      {stage0_61[168]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[66],stage1_62[132],stage1_61[158],stage1_60[188]}
   );
   gpc615_5 gpc2393 (
      {stage0_60[497], stage0_60[498], stage0_60[499], stage0_60[500], stage0_60[501]},
      {stage0_61[169]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[67],stage1_62[133],stage1_61[159],stage1_60[189]}
   );
   gpc606_5 gpc2394 (
      {stage0_61[170], stage0_61[171], stage0_61[172], stage0_61[173], stage0_61[174], stage0_61[175]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[55],stage1_63[68],stage1_62[134],stage1_61[160]}
   );
   gpc606_5 gpc2395 (
      {stage0_61[176], stage0_61[177], stage0_61[178], stage0_61[179], stage0_61[180], stage0_61[181]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[56],stage1_63[69],stage1_62[135],stage1_61[161]}
   );
   gpc606_5 gpc2396 (
      {stage0_61[182], stage0_61[183], stage0_61[184], stage0_61[185], stage0_61[186], stage0_61[187]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[57],stage1_63[70],stage1_62[136],stage1_61[162]}
   );
   gpc606_5 gpc2397 (
      {stage0_61[188], stage0_61[189], stage0_61[190], stage0_61[191], stage0_61[192], stage0_61[193]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[58],stage1_63[71],stage1_62[137],stage1_61[163]}
   );
   gpc606_5 gpc2398 (
      {stage0_61[194], stage0_61[195], stage0_61[196], stage0_61[197], stage0_61[198], stage0_61[199]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[59],stage1_63[72],stage1_62[138],stage1_61[164]}
   );
   gpc606_5 gpc2399 (
      {stage0_61[200], stage0_61[201], stage0_61[202], stage0_61[203], stage0_61[204], stage0_61[205]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[60],stage1_63[73],stage1_62[139],stage1_61[165]}
   );
   gpc606_5 gpc2400 (
      {stage0_61[206], stage0_61[207], stage0_61[208], stage0_61[209], stage0_61[210], stage0_61[211]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[61],stage1_63[74],stage1_62[140],stage1_61[166]}
   );
   gpc606_5 gpc2401 (
      {stage0_61[212], stage0_61[213], stage0_61[214], stage0_61[215], stage0_61[216], stage0_61[217]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[62],stage1_63[75],stage1_62[141],stage1_61[167]}
   );
   gpc606_5 gpc2402 (
      {stage0_61[218], stage0_61[219], stage0_61[220], stage0_61[221], stage0_61[222], stage0_61[223]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[63],stage1_63[76],stage1_62[142],stage1_61[168]}
   );
   gpc606_5 gpc2403 (
      {stage0_61[224], stage0_61[225], stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[64],stage1_63[77],stage1_62[143],stage1_61[169]}
   );
   gpc606_5 gpc2404 (
      {stage0_61[230], stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[65],stage1_63[78],stage1_62[144],stage1_61[170]}
   );
   gpc606_5 gpc2405 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240], stage0_61[241]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[66],stage1_63[79],stage1_62[145],stage1_61[171]}
   );
   gpc606_5 gpc2406 (
      {stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245], stage0_61[246], stage0_61[247]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[67],stage1_63[80],stage1_62[146],stage1_61[172]}
   );
   gpc606_5 gpc2407 (
      {stage0_61[248], stage0_61[249], stage0_61[250], stage0_61[251], stage0_61[252], stage0_61[253]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[68],stage1_63[81],stage1_62[147],stage1_61[173]}
   );
   gpc606_5 gpc2408 (
      {stage0_61[254], stage0_61[255], stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[69],stage1_63[82],stage1_62[148],stage1_61[174]}
   );
   gpc606_5 gpc2409 (
      {stage0_61[260], stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[70],stage1_63[83],stage1_62[149],stage1_61[175]}
   );
   gpc606_5 gpc2410 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270], stage0_61[271]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[71],stage1_63[84],stage1_62[150],stage1_61[176]}
   );
   gpc606_5 gpc2411 (
      {stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275], stage0_61[276], stage0_61[277]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[72],stage1_63[85],stage1_62[151],stage1_61[177]}
   );
   gpc606_5 gpc2412 (
      {stage0_61[278], stage0_61[279], stage0_61[280], stage0_61[281], stage0_61[282], stage0_61[283]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[73],stage1_63[86],stage1_62[152],stage1_61[178]}
   );
   gpc606_5 gpc2413 (
      {stage0_61[284], stage0_61[285], stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[74],stage1_63[87],stage1_62[153],stage1_61[179]}
   );
   gpc606_5 gpc2414 (
      {stage0_61[290], stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[75],stage1_63[88],stage1_62[154],stage1_61[180]}
   );
   gpc606_5 gpc2415 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300], stage0_61[301]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[76],stage1_63[89],stage1_62[155],stage1_61[181]}
   );
   gpc606_5 gpc2416 (
      {stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305], stage0_61[306], stage0_61[307]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[77],stage1_63[90],stage1_62[156],stage1_61[182]}
   );
   gpc606_5 gpc2417 (
      {stage0_61[308], stage0_61[309], stage0_61[310], stage0_61[311], stage0_61[312], stage0_61[313]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[78],stage1_63[91],stage1_62[157],stage1_61[183]}
   );
   gpc606_5 gpc2418 (
      {stage0_61[314], stage0_61[315], stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[79],stage1_63[92],stage1_62[158],stage1_61[184]}
   );
   gpc606_5 gpc2419 (
      {stage0_61[320], stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[80],stage1_63[93],stage1_62[159],stage1_61[185]}
   );
   gpc606_5 gpc2420 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330], stage0_61[331]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[81],stage1_63[94],stage1_62[160],stage1_61[186]}
   );
   gpc606_5 gpc2421 (
      {stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335], stage0_61[336], stage0_61[337]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[82],stage1_63[95],stage1_62[161],stage1_61[187]}
   );
   gpc606_5 gpc2422 (
      {stage0_61[338], stage0_61[339], stage0_61[340], stage0_61[341], stage0_61[342], stage0_61[343]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[83],stage1_63[96],stage1_62[162],stage1_61[188]}
   );
   gpc606_5 gpc2423 (
      {stage0_61[344], stage0_61[345], stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[84],stage1_63[97],stage1_62[163],stage1_61[189]}
   );
   gpc606_5 gpc2424 (
      {stage0_61[350], stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[85],stage1_63[98],stage1_62[164],stage1_61[190]}
   );
   gpc606_5 gpc2425 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360], stage0_61[361]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[86],stage1_63[99],stage1_62[165],stage1_61[191]}
   );
   gpc606_5 gpc2426 (
      {stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365], stage0_61[366], stage0_61[367]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[87],stage1_63[100],stage1_62[166],stage1_61[192]}
   );
   gpc606_5 gpc2427 (
      {stage0_61[368], stage0_61[369], stage0_61[370], stage0_61[371], stage0_61[372], stage0_61[373]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[88],stage1_63[101],stage1_62[167],stage1_61[193]}
   );
   gpc606_5 gpc2428 (
      {stage0_61[374], stage0_61[375], stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[89],stage1_63[102],stage1_62[168],stage1_61[194]}
   );
   gpc606_5 gpc2429 (
      {stage0_61[380], stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[90],stage1_63[103],stage1_62[169],stage1_61[195]}
   );
   gpc606_5 gpc2430 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390], stage0_61[391]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[91],stage1_63[104],stage1_62[170],stage1_61[196]}
   );
   gpc606_5 gpc2431 (
      {stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395], stage0_61[396], stage0_61[397]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[92],stage1_63[105],stage1_62[171],stage1_61[197]}
   );
   gpc606_5 gpc2432 (
      {stage0_61[398], stage0_61[399], stage0_61[400], stage0_61[401], stage0_61[402], stage0_61[403]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[93],stage1_63[106],stage1_62[172],stage1_61[198]}
   );
   gpc606_5 gpc2433 (
      {stage0_61[404], stage0_61[405], stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[94],stage1_63[107],stage1_62[173],stage1_61[199]}
   );
   gpc606_5 gpc2434 (
      {stage0_61[410], stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[95],stage1_63[108],stage1_62[174],stage1_61[200]}
   );
   gpc606_5 gpc2435 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420], stage0_61[421]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[96],stage1_63[109],stage1_62[175],stage1_61[201]}
   );
   gpc606_5 gpc2436 (
      {stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425], stage0_61[426], stage0_61[427]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[97],stage1_63[110],stage1_62[176],stage1_61[202]}
   );
   gpc606_5 gpc2437 (
      {stage0_61[428], stage0_61[429], stage0_61[430], stage0_61[431], stage0_61[432], stage0_61[433]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[98],stage1_63[111],stage1_62[177],stage1_61[203]}
   );
   gpc606_5 gpc2438 (
      {stage0_61[434], stage0_61[435], stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[99],stage1_63[112],stage1_62[178],stage1_61[204]}
   );
   gpc606_5 gpc2439 (
      {stage0_61[440], stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[100],stage1_63[113],stage1_62[179],stage1_61[205]}
   );
   gpc606_5 gpc2440 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450], stage0_61[451]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[101],stage1_63[114],stage1_62[180],stage1_61[206]}
   );
   gpc606_5 gpc2441 (
      {stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455], stage0_61[456], stage0_61[457]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[102],stage1_63[115],stage1_62[181],stage1_61[207]}
   );
   gpc606_5 gpc2442 (
      {stage0_61[458], stage0_61[459], stage0_61[460], stage0_61[461], stage0_61[462], stage0_61[463]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[103],stage1_63[116],stage1_62[182],stage1_61[208]}
   );
   gpc606_5 gpc2443 (
      {stage0_61[464], stage0_61[465], stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[104],stage1_63[117],stage1_62[183],stage1_61[209]}
   );
   gpc606_5 gpc2444 (
      {stage0_61[470], stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[105],stage1_63[118],stage1_62[184],stage1_61[210]}
   );
   gpc606_5 gpc2445 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480], stage0_61[481]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[106],stage1_63[119],stage1_62[185],stage1_61[211]}
   );
   gpc606_5 gpc2446 (
      {stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485], stage0_61[486], stage0_61[487]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[107],stage1_63[120],stage1_62[186],stage1_61[212]}
   );
   gpc606_5 gpc2447 (
      {stage0_61[488], stage0_61[489], stage0_61[490], stage0_61[491], stage0_61[492], stage0_61[493]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[108],stage1_63[121],stage1_62[187],stage1_61[213]}
   );
   gpc606_5 gpc2448 (
      {stage0_61[494], stage0_61[495], stage0_61[496], stage0_61[497], stage0_61[498], stage0_61[499]},
      {stage0_63[324], stage0_63[325], stage0_63[326], stage0_63[327], stage0_63[328], stage0_63[329]},
      {stage1_65[54],stage1_64[109],stage1_63[122],stage1_62[188],stage1_61[214]}
   );
   gpc606_5 gpc2449 (
      {stage0_61[500], stage0_61[501], stage0_61[502], stage0_61[503], stage0_61[504], stage0_61[505]},
      {stage0_63[330], stage0_63[331], stage0_63[332], stage0_63[333], stage0_63[334], stage0_63[335]},
      {stage1_65[55],stage1_64[110],stage1_63[123],stage1_62[189],stage1_61[215]}
   );
   gpc606_5 gpc2450 (
      {stage0_61[506], stage0_61[507], stage0_61[508], stage0_61[509], stage0_61[510], stage0_61[511]},
      {stage0_63[336], stage0_63[337], stage0_63[338], stage0_63[339], stage0_63[340], stage0_63[341]},
      {stage1_65[56],stage1_64[111],stage1_63[124],stage1_62[190],stage1_61[216]}
   );
   gpc1_1 gpc2451 (
      {stage0_1[481]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2452 (
      {stage0_1[482]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2453 (
      {stage0_1[483]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2454 (
      {stage0_1[484]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2455 (
      {stage0_1[485]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[486]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[487]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[488]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[489]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[490]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[491]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[492]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[493]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[494]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[495]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[496]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[497]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[498]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[499]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[500]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[501]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[502]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[503]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[504]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[505]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[506]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[507]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[508]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[509]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[510]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[511]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2482 (
      {stage0_2[429]},
      {stage1_2[138]}
   );
   gpc1_1 gpc2483 (
      {stage0_2[430]},
      {stage1_2[139]}
   );
   gpc1_1 gpc2484 (
      {stage0_2[431]},
      {stage1_2[140]}
   );
   gpc1_1 gpc2485 (
      {stage0_2[432]},
      {stage1_2[141]}
   );
   gpc1_1 gpc2486 (
      {stage0_2[433]},
      {stage1_2[142]}
   );
   gpc1_1 gpc2487 (
      {stage0_2[434]},
      {stage1_2[143]}
   );
   gpc1_1 gpc2488 (
      {stage0_2[435]},
      {stage1_2[144]}
   );
   gpc1_1 gpc2489 (
      {stage0_2[436]},
      {stage1_2[145]}
   );
   gpc1_1 gpc2490 (
      {stage0_2[437]},
      {stage1_2[146]}
   );
   gpc1_1 gpc2491 (
      {stage0_2[438]},
      {stage1_2[147]}
   );
   gpc1_1 gpc2492 (
      {stage0_2[439]},
      {stage1_2[148]}
   );
   gpc1_1 gpc2493 (
      {stage0_2[440]},
      {stage1_2[149]}
   );
   gpc1_1 gpc2494 (
      {stage0_2[441]},
      {stage1_2[150]}
   );
   gpc1_1 gpc2495 (
      {stage0_2[442]},
      {stage1_2[151]}
   );
   gpc1_1 gpc2496 (
      {stage0_2[443]},
      {stage1_2[152]}
   );
   gpc1_1 gpc2497 (
      {stage0_2[444]},
      {stage1_2[153]}
   );
   gpc1_1 gpc2498 (
      {stage0_2[445]},
      {stage1_2[154]}
   );
   gpc1_1 gpc2499 (
      {stage0_2[446]},
      {stage1_2[155]}
   );
   gpc1_1 gpc2500 (
      {stage0_2[447]},
      {stage1_2[156]}
   );
   gpc1_1 gpc2501 (
      {stage0_2[448]},
      {stage1_2[157]}
   );
   gpc1_1 gpc2502 (
      {stage0_2[449]},
      {stage1_2[158]}
   );
   gpc1_1 gpc2503 (
      {stage0_2[450]},
      {stage1_2[159]}
   );
   gpc1_1 gpc2504 (
      {stage0_2[451]},
      {stage1_2[160]}
   );
   gpc1_1 gpc2505 (
      {stage0_2[452]},
      {stage1_2[161]}
   );
   gpc1_1 gpc2506 (
      {stage0_2[453]},
      {stage1_2[162]}
   );
   gpc1_1 gpc2507 (
      {stage0_2[454]},
      {stage1_2[163]}
   );
   gpc1_1 gpc2508 (
      {stage0_2[455]},
      {stage1_2[164]}
   );
   gpc1_1 gpc2509 (
      {stage0_2[456]},
      {stage1_2[165]}
   );
   gpc1_1 gpc2510 (
      {stage0_2[457]},
      {stage1_2[166]}
   );
   gpc1_1 gpc2511 (
      {stage0_2[458]},
      {stage1_2[167]}
   );
   gpc1_1 gpc2512 (
      {stage0_2[459]},
      {stage1_2[168]}
   );
   gpc1_1 gpc2513 (
      {stage0_2[460]},
      {stage1_2[169]}
   );
   gpc1_1 gpc2514 (
      {stage0_2[461]},
      {stage1_2[170]}
   );
   gpc1_1 gpc2515 (
      {stage0_2[462]},
      {stage1_2[171]}
   );
   gpc1_1 gpc2516 (
      {stage0_2[463]},
      {stage1_2[172]}
   );
   gpc1_1 gpc2517 (
      {stage0_2[464]},
      {stage1_2[173]}
   );
   gpc1_1 gpc2518 (
      {stage0_2[465]},
      {stage1_2[174]}
   );
   gpc1_1 gpc2519 (
      {stage0_2[466]},
      {stage1_2[175]}
   );
   gpc1_1 gpc2520 (
      {stage0_2[467]},
      {stage1_2[176]}
   );
   gpc1_1 gpc2521 (
      {stage0_2[468]},
      {stage1_2[177]}
   );
   gpc1_1 gpc2522 (
      {stage0_2[469]},
      {stage1_2[178]}
   );
   gpc1_1 gpc2523 (
      {stage0_2[470]},
      {stage1_2[179]}
   );
   gpc1_1 gpc2524 (
      {stage0_2[471]},
      {stage1_2[180]}
   );
   gpc1_1 gpc2525 (
      {stage0_2[472]},
      {stage1_2[181]}
   );
   gpc1_1 gpc2526 (
      {stage0_2[473]},
      {stage1_2[182]}
   );
   gpc1_1 gpc2527 (
      {stage0_2[474]},
      {stage1_2[183]}
   );
   gpc1_1 gpc2528 (
      {stage0_2[475]},
      {stage1_2[184]}
   );
   gpc1_1 gpc2529 (
      {stage0_2[476]},
      {stage1_2[185]}
   );
   gpc1_1 gpc2530 (
      {stage0_2[477]},
      {stage1_2[186]}
   );
   gpc1_1 gpc2531 (
      {stage0_2[478]},
      {stage1_2[187]}
   );
   gpc1_1 gpc2532 (
      {stage0_2[479]},
      {stage1_2[188]}
   );
   gpc1_1 gpc2533 (
      {stage0_2[480]},
      {stage1_2[189]}
   );
   gpc1_1 gpc2534 (
      {stage0_2[481]},
      {stage1_2[190]}
   );
   gpc1_1 gpc2535 (
      {stage0_2[482]},
      {stage1_2[191]}
   );
   gpc1_1 gpc2536 (
      {stage0_2[483]},
      {stage1_2[192]}
   );
   gpc1_1 gpc2537 (
      {stage0_2[484]},
      {stage1_2[193]}
   );
   gpc1_1 gpc2538 (
      {stage0_2[485]},
      {stage1_2[194]}
   );
   gpc1_1 gpc2539 (
      {stage0_2[486]},
      {stage1_2[195]}
   );
   gpc1_1 gpc2540 (
      {stage0_2[487]},
      {stage1_2[196]}
   );
   gpc1_1 gpc2541 (
      {stage0_2[488]},
      {stage1_2[197]}
   );
   gpc1_1 gpc2542 (
      {stage0_2[489]},
      {stage1_2[198]}
   );
   gpc1_1 gpc2543 (
      {stage0_2[490]},
      {stage1_2[199]}
   );
   gpc1_1 gpc2544 (
      {stage0_2[491]},
      {stage1_2[200]}
   );
   gpc1_1 gpc2545 (
      {stage0_2[492]},
      {stage1_2[201]}
   );
   gpc1_1 gpc2546 (
      {stage0_2[493]},
      {stage1_2[202]}
   );
   gpc1_1 gpc2547 (
      {stage0_2[494]},
      {stage1_2[203]}
   );
   gpc1_1 gpc2548 (
      {stage0_2[495]},
      {stage1_2[204]}
   );
   gpc1_1 gpc2549 (
      {stage0_2[496]},
      {stage1_2[205]}
   );
   gpc1_1 gpc2550 (
      {stage0_2[497]},
      {stage1_2[206]}
   );
   gpc1_1 gpc2551 (
      {stage0_2[498]},
      {stage1_2[207]}
   );
   gpc1_1 gpc2552 (
      {stage0_2[499]},
      {stage1_2[208]}
   );
   gpc1_1 gpc2553 (
      {stage0_2[500]},
      {stage1_2[209]}
   );
   gpc1_1 gpc2554 (
      {stage0_2[501]},
      {stage1_2[210]}
   );
   gpc1_1 gpc2555 (
      {stage0_2[502]},
      {stage1_2[211]}
   );
   gpc1_1 gpc2556 (
      {stage0_2[503]},
      {stage1_2[212]}
   );
   gpc1_1 gpc2557 (
      {stage0_2[504]},
      {stage1_2[213]}
   );
   gpc1_1 gpc2558 (
      {stage0_2[505]},
      {stage1_2[214]}
   );
   gpc1_1 gpc2559 (
      {stage0_2[506]},
      {stage1_2[215]}
   );
   gpc1_1 gpc2560 (
      {stage0_2[507]},
      {stage1_2[216]}
   );
   gpc1_1 gpc2561 (
      {stage0_2[508]},
      {stage1_2[217]}
   );
   gpc1_1 gpc2562 (
      {stage0_2[509]},
      {stage1_2[218]}
   );
   gpc1_1 gpc2563 (
      {stage0_2[510]},
      {stage1_2[219]}
   );
   gpc1_1 gpc2564 (
      {stage0_2[511]},
      {stage1_2[220]}
   );
   gpc1_1 gpc2565 (
      {stage0_3[372]},
      {stage1_3[182]}
   );
   gpc1_1 gpc2566 (
      {stage0_3[373]},
      {stage1_3[183]}
   );
   gpc1_1 gpc2567 (
      {stage0_3[374]},
      {stage1_3[184]}
   );
   gpc1_1 gpc2568 (
      {stage0_3[375]},
      {stage1_3[185]}
   );
   gpc1_1 gpc2569 (
      {stage0_3[376]},
      {stage1_3[186]}
   );
   gpc1_1 gpc2570 (
      {stage0_3[377]},
      {stage1_3[187]}
   );
   gpc1_1 gpc2571 (
      {stage0_3[378]},
      {stage1_3[188]}
   );
   gpc1_1 gpc2572 (
      {stage0_3[379]},
      {stage1_3[189]}
   );
   gpc1_1 gpc2573 (
      {stage0_3[380]},
      {stage1_3[190]}
   );
   gpc1_1 gpc2574 (
      {stage0_3[381]},
      {stage1_3[191]}
   );
   gpc1_1 gpc2575 (
      {stage0_3[382]},
      {stage1_3[192]}
   );
   gpc1_1 gpc2576 (
      {stage0_3[383]},
      {stage1_3[193]}
   );
   gpc1_1 gpc2577 (
      {stage0_3[384]},
      {stage1_3[194]}
   );
   gpc1_1 gpc2578 (
      {stage0_3[385]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2579 (
      {stage0_3[386]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2580 (
      {stage0_3[387]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2581 (
      {stage0_3[388]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2582 (
      {stage0_3[389]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2583 (
      {stage0_3[390]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2584 (
      {stage0_3[391]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2585 (
      {stage0_3[392]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2586 (
      {stage0_3[393]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2587 (
      {stage0_3[394]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2588 (
      {stage0_3[395]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2589 (
      {stage0_3[396]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2590 (
      {stage0_3[397]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2591 (
      {stage0_3[398]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2592 (
      {stage0_3[399]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2593 (
      {stage0_3[400]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2594 (
      {stage0_3[401]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2595 (
      {stage0_3[402]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2596 (
      {stage0_3[403]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2597 (
      {stage0_3[404]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2598 (
      {stage0_3[405]},
      {stage1_3[215]}
   );
   gpc1_1 gpc2599 (
      {stage0_3[406]},
      {stage1_3[216]}
   );
   gpc1_1 gpc2600 (
      {stage0_3[407]},
      {stage1_3[217]}
   );
   gpc1_1 gpc2601 (
      {stage0_3[408]},
      {stage1_3[218]}
   );
   gpc1_1 gpc2602 (
      {stage0_3[409]},
      {stage1_3[219]}
   );
   gpc1_1 gpc2603 (
      {stage0_3[410]},
      {stage1_3[220]}
   );
   gpc1_1 gpc2604 (
      {stage0_3[411]},
      {stage1_3[221]}
   );
   gpc1_1 gpc2605 (
      {stage0_3[412]},
      {stage1_3[222]}
   );
   gpc1_1 gpc2606 (
      {stage0_3[413]},
      {stage1_3[223]}
   );
   gpc1_1 gpc2607 (
      {stage0_3[414]},
      {stage1_3[224]}
   );
   gpc1_1 gpc2608 (
      {stage0_3[415]},
      {stage1_3[225]}
   );
   gpc1_1 gpc2609 (
      {stage0_3[416]},
      {stage1_3[226]}
   );
   gpc1_1 gpc2610 (
      {stage0_3[417]},
      {stage1_3[227]}
   );
   gpc1_1 gpc2611 (
      {stage0_3[418]},
      {stage1_3[228]}
   );
   gpc1_1 gpc2612 (
      {stage0_3[419]},
      {stage1_3[229]}
   );
   gpc1_1 gpc2613 (
      {stage0_3[420]},
      {stage1_3[230]}
   );
   gpc1_1 gpc2614 (
      {stage0_3[421]},
      {stage1_3[231]}
   );
   gpc1_1 gpc2615 (
      {stage0_3[422]},
      {stage1_3[232]}
   );
   gpc1_1 gpc2616 (
      {stage0_3[423]},
      {stage1_3[233]}
   );
   gpc1_1 gpc2617 (
      {stage0_3[424]},
      {stage1_3[234]}
   );
   gpc1_1 gpc2618 (
      {stage0_3[425]},
      {stage1_3[235]}
   );
   gpc1_1 gpc2619 (
      {stage0_3[426]},
      {stage1_3[236]}
   );
   gpc1_1 gpc2620 (
      {stage0_3[427]},
      {stage1_3[237]}
   );
   gpc1_1 gpc2621 (
      {stage0_3[428]},
      {stage1_3[238]}
   );
   gpc1_1 gpc2622 (
      {stage0_3[429]},
      {stage1_3[239]}
   );
   gpc1_1 gpc2623 (
      {stage0_3[430]},
      {stage1_3[240]}
   );
   gpc1_1 gpc2624 (
      {stage0_3[431]},
      {stage1_3[241]}
   );
   gpc1_1 gpc2625 (
      {stage0_3[432]},
      {stage1_3[242]}
   );
   gpc1_1 gpc2626 (
      {stage0_3[433]},
      {stage1_3[243]}
   );
   gpc1_1 gpc2627 (
      {stage0_3[434]},
      {stage1_3[244]}
   );
   gpc1_1 gpc2628 (
      {stage0_3[435]},
      {stage1_3[245]}
   );
   gpc1_1 gpc2629 (
      {stage0_3[436]},
      {stage1_3[246]}
   );
   gpc1_1 gpc2630 (
      {stage0_3[437]},
      {stage1_3[247]}
   );
   gpc1_1 gpc2631 (
      {stage0_3[438]},
      {stage1_3[248]}
   );
   gpc1_1 gpc2632 (
      {stage0_3[439]},
      {stage1_3[249]}
   );
   gpc1_1 gpc2633 (
      {stage0_3[440]},
      {stage1_3[250]}
   );
   gpc1_1 gpc2634 (
      {stage0_3[441]},
      {stage1_3[251]}
   );
   gpc1_1 gpc2635 (
      {stage0_3[442]},
      {stage1_3[252]}
   );
   gpc1_1 gpc2636 (
      {stage0_3[443]},
      {stage1_3[253]}
   );
   gpc1_1 gpc2637 (
      {stage0_3[444]},
      {stage1_3[254]}
   );
   gpc1_1 gpc2638 (
      {stage0_3[445]},
      {stage1_3[255]}
   );
   gpc1_1 gpc2639 (
      {stage0_3[446]},
      {stage1_3[256]}
   );
   gpc1_1 gpc2640 (
      {stage0_3[447]},
      {stage1_3[257]}
   );
   gpc1_1 gpc2641 (
      {stage0_3[448]},
      {stage1_3[258]}
   );
   gpc1_1 gpc2642 (
      {stage0_3[449]},
      {stage1_3[259]}
   );
   gpc1_1 gpc2643 (
      {stage0_3[450]},
      {stage1_3[260]}
   );
   gpc1_1 gpc2644 (
      {stage0_3[451]},
      {stage1_3[261]}
   );
   gpc1_1 gpc2645 (
      {stage0_3[452]},
      {stage1_3[262]}
   );
   gpc1_1 gpc2646 (
      {stage0_3[453]},
      {stage1_3[263]}
   );
   gpc1_1 gpc2647 (
      {stage0_3[454]},
      {stage1_3[264]}
   );
   gpc1_1 gpc2648 (
      {stage0_3[455]},
      {stage1_3[265]}
   );
   gpc1_1 gpc2649 (
      {stage0_3[456]},
      {stage1_3[266]}
   );
   gpc1_1 gpc2650 (
      {stage0_3[457]},
      {stage1_3[267]}
   );
   gpc1_1 gpc2651 (
      {stage0_3[458]},
      {stage1_3[268]}
   );
   gpc1_1 gpc2652 (
      {stage0_3[459]},
      {stage1_3[269]}
   );
   gpc1_1 gpc2653 (
      {stage0_3[460]},
      {stage1_3[270]}
   );
   gpc1_1 gpc2654 (
      {stage0_3[461]},
      {stage1_3[271]}
   );
   gpc1_1 gpc2655 (
      {stage0_3[462]},
      {stage1_3[272]}
   );
   gpc1_1 gpc2656 (
      {stage0_3[463]},
      {stage1_3[273]}
   );
   gpc1_1 gpc2657 (
      {stage0_3[464]},
      {stage1_3[274]}
   );
   gpc1_1 gpc2658 (
      {stage0_3[465]},
      {stage1_3[275]}
   );
   gpc1_1 gpc2659 (
      {stage0_3[466]},
      {stage1_3[276]}
   );
   gpc1_1 gpc2660 (
      {stage0_3[467]},
      {stage1_3[277]}
   );
   gpc1_1 gpc2661 (
      {stage0_3[468]},
      {stage1_3[278]}
   );
   gpc1_1 gpc2662 (
      {stage0_3[469]},
      {stage1_3[279]}
   );
   gpc1_1 gpc2663 (
      {stage0_3[470]},
      {stage1_3[280]}
   );
   gpc1_1 gpc2664 (
      {stage0_3[471]},
      {stage1_3[281]}
   );
   gpc1_1 gpc2665 (
      {stage0_3[472]},
      {stage1_3[282]}
   );
   gpc1_1 gpc2666 (
      {stage0_3[473]},
      {stage1_3[283]}
   );
   gpc1_1 gpc2667 (
      {stage0_3[474]},
      {stage1_3[284]}
   );
   gpc1_1 gpc2668 (
      {stage0_3[475]},
      {stage1_3[285]}
   );
   gpc1_1 gpc2669 (
      {stage0_3[476]},
      {stage1_3[286]}
   );
   gpc1_1 gpc2670 (
      {stage0_3[477]},
      {stage1_3[287]}
   );
   gpc1_1 gpc2671 (
      {stage0_3[478]},
      {stage1_3[288]}
   );
   gpc1_1 gpc2672 (
      {stage0_3[479]},
      {stage1_3[289]}
   );
   gpc1_1 gpc2673 (
      {stage0_3[480]},
      {stage1_3[290]}
   );
   gpc1_1 gpc2674 (
      {stage0_3[481]},
      {stage1_3[291]}
   );
   gpc1_1 gpc2675 (
      {stage0_3[482]},
      {stage1_3[292]}
   );
   gpc1_1 gpc2676 (
      {stage0_3[483]},
      {stage1_3[293]}
   );
   gpc1_1 gpc2677 (
      {stage0_3[484]},
      {stage1_3[294]}
   );
   gpc1_1 gpc2678 (
      {stage0_3[485]},
      {stage1_3[295]}
   );
   gpc1_1 gpc2679 (
      {stage0_3[486]},
      {stage1_3[296]}
   );
   gpc1_1 gpc2680 (
      {stage0_3[487]},
      {stage1_3[297]}
   );
   gpc1_1 gpc2681 (
      {stage0_3[488]},
      {stage1_3[298]}
   );
   gpc1_1 gpc2682 (
      {stage0_3[489]},
      {stage1_3[299]}
   );
   gpc1_1 gpc2683 (
      {stage0_3[490]},
      {stage1_3[300]}
   );
   gpc1_1 gpc2684 (
      {stage0_3[491]},
      {stage1_3[301]}
   );
   gpc1_1 gpc2685 (
      {stage0_3[492]},
      {stage1_3[302]}
   );
   gpc1_1 gpc2686 (
      {stage0_3[493]},
      {stage1_3[303]}
   );
   gpc1_1 gpc2687 (
      {stage0_3[494]},
      {stage1_3[304]}
   );
   gpc1_1 gpc2688 (
      {stage0_3[495]},
      {stage1_3[305]}
   );
   gpc1_1 gpc2689 (
      {stage0_3[496]},
      {stage1_3[306]}
   );
   gpc1_1 gpc2690 (
      {stage0_3[497]},
      {stage1_3[307]}
   );
   gpc1_1 gpc2691 (
      {stage0_3[498]},
      {stage1_3[308]}
   );
   gpc1_1 gpc2692 (
      {stage0_3[499]},
      {stage1_3[309]}
   );
   gpc1_1 gpc2693 (
      {stage0_3[500]},
      {stage1_3[310]}
   );
   gpc1_1 gpc2694 (
      {stage0_3[501]},
      {stage1_3[311]}
   );
   gpc1_1 gpc2695 (
      {stage0_3[502]},
      {stage1_3[312]}
   );
   gpc1_1 gpc2696 (
      {stage0_3[503]},
      {stage1_3[313]}
   );
   gpc1_1 gpc2697 (
      {stage0_3[504]},
      {stage1_3[314]}
   );
   gpc1_1 gpc2698 (
      {stage0_3[505]},
      {stage1_3[315]}
   );
   gpc1_1 gpc2699 (
      {stage0_3[506]},
      {stage1_3[316]}
   );
   gpc1_1 gpc2700 (
      {stage0_3[507]},
      {stage1_3[317]}
   );
   gpc1_1 gpc2701 (
      {stage0_3[508]},
      {stage1_3[318]}
   );
   gpc1_1 gpc2702 (
      {stage0_3[509]},
      {stage1_3[319]}
   );
   gpc1_1 gpc2703 (
      {stage0_3[510]},
      {stage1_3[320]}
   );
   gpc1_1 gpc2704 (
      {stage0_3[511]},
      {stage1_3[321]}
   );
   gpc1_1 gpc2705 (
      {stage0_5[468]},
      {stage1_5[173]}
   );
   gpc1_1 gpc2706 (
      {stage0_5[469]},
      {stage1_5[174]}
   );
   gpc1_1 gpc2707 (
      {stage0_5[470]},
      {stage1_5[175]}
   );
   gpc1_1 gpc2708 (
      {stage0_5[471]},
      {stage1_5[176]}
   );
   gpc1_1 gpc2709 (
      {stage0_5[472]},
      {stage1_5[177]}
   );
   gpc1_1 gpc2710 (
      {stage0_5[473]},
      {stage1_5[178]}
   );
   gpc1_1 gpc2711 (
      {stage0_5[474]},
      {stage1_5[179]}
   );
   gpc1_1 gpc2712 (
      {stage0_5[475]},
      {stage1_5[180]}
   );
   gpc1_1 gpc2713 (
      {stage0_5[476]},
      {stage1_5[181]}
   );
   gpc1_1 gpc2714 (
      {stage0_5[477]},
      {stage1_5[182]}
   );
   gpc1_1 gpc2715 (
      {stage0_5[478]},
      {stage1_5[183]}
   );
   gpc1_1 gpc2716 (
      {stage0_5[479]},
      {stage1_5[184]}
   );
   gpc1_1 gpc2717 (
      {stage0_5[480]},
      {stage1_5[185]}
   );
   gpc1_1 gpc2718 (
      {stage0_5[481]},
      {stage1_5[186]}
   );
   gpc1_1 gpc2719 (
      {stage0_5[482]},
      {stage1_5[187]}
   );
   gpc1_1 gpc2720 (
      {stage0_5[483]},
      {stage1_5[188]}
   );
   gpc1_1 gpc2721 (
      {stage0_5[484]},
      {stage1_5[189]}
   );
   gpc1_1 gpc2722 (
      {stage0_5[485]},
      {stage1_5[190]}
   );
   gpc1_1 gpc2723 (
      {stage0_5[486]},
      {stage1_5[191]}
   );
   gpc1_1 gpc2724 (
      {stage0_5[487]},
      {stage1_5[192]}
   );
   gpc1_1 gpc2725 (
      {stage0_5[488]},
      {stage1_5[193]}
   );
   gpc1_1 gpc2726 (
      {stage0_5[489]},
      {stage1_5[194]}
   );
   gpc1_1 gpc2727 (
      {stage0_5[490]},
      {stage1_5[195]}
   );
   gpc1_1 gpc2728 (
      {stage0_5[491]},
      {stage1_5[196]}
   );
   gpc1_1 gpc2729 (
      {stage0_5[492]},
      {stage1_5[197]}
   );
   gpc1_1 gpc2730 (
      {stage0_5[493]},
      {stage1_5[198]}
   );
   gpc1_1 gpc2731 (
      {stage0_5[494]},
      {stage1_5[199]}
   );
   gpc1_1 gpc2732 (
      {stage0_5[495]},
      {stage1_5[200]}
   );
   gpc1_1 gpc2733 (
      {stage0_5[496]},
      {stage1_5[201]}
   );
   gpc1_1 gpc2734 (
      {stage0_5[497]},
      {stage1_5[202]}
   );
   gpc1_1 gpc2735 (
      {stage0_5[498]},
      {stage1_5[203]}
   );
   gpc1_1 gpc2736 (
      {stage0_5[499]},
      {stage1_5[204]}
   );
   gpc1_1 gpc2737 (
      {stage0_5[500]},
      {stage1_5[205]}
   );
   gpc1_1 gpc2738 (
      {stage0_5[501]},
      {stage1_5[206]}
   );
   gpc1_1 gpc2739 (
      {stage0_5[502]},
      {stage1_5[207]}
   );
   gpc1_1 gpc2740 (
      {stage0_5[503]},
      {stage1_5[208]}
   );
   gpc1_1 gpc2741 (
      {stage0_5[504]},
      {stage1_5[209]}
   );
   gpc1_1 gpc2742 (
      {stage0_5[505]},
      {stage1_5[210]}
   );
   gpc1_1 gpc2743 (
      {stage0_5[506]},
      {stage1_5[211]}
   );
   gpc1_1 gpc2744 (
      {stage0_5[507]},
      {stage1_5[212]}
   );
   gpc1_1 gpc2745 (
      {stage0_5[508]},
      {stage1_5[213]}
   );
   gpc1_1 gpc2746 (
      {stage0_5[509]},
      {stage1_5[214]}
   );
   gpc1_1 gpc2747 (
      {stage0_5[510]},
      {stage1_5[215]}
   );
   gpc1_1 gpc2748 (
      {stage0_5[511]},
      {stage1_5[216]}
   );
   gpc1_1 gpc2749 (
      {stage0_6[493]},
      {stage1_6[161]}
   );
   gpc1_1 gpc2750 (
      {stage0_6[494]},
      {stage1_6[162]}
   );
   gpc1_1 gpc2751 (
      {stage0_6[495]},
      {stage1_6[163]}
   );
   gpc1_1 gpc2752 (
      {stage0_6[496]},
      {stage1_6[164]}
   );
   gpc1_1 gpc2753 (
      {stage0_6[497]},
      {stage1_6[165]}
   );
   gpc1_1 gpc2754 (
      {stage0_6[498]},
      {stage1_6[166]}
   );
   gpc1_1 gpc2755 (
      {stage0_6[499]},
      {stage1_6[167]}
   );
   gpc1_1 gpc2756 (
      {stage0_6[500]},
      {stage1_6[168]}
   );
   gpc1_1 gpc2757 (
      {stage0_6[501]},
      {stage1_6[169]}
   );
   gpc1_1 gpc2758 (
      {stage0_6[502]},
      {stage1_6[170]}
   );
   gpc1_1 gpc2759 (
      {stage0_6[503]},
      {stage1_6[171]}
   );
   gpc1_1 gpc2760 (
      {stage0_6[504]},
      {stage1_6[172]}
   );
   gpc1_1 gpc2761 (
      {stage0_6[505]},
      {stage1_6[173]}
   );
   gpc1_1 gpc2762 (
      {stage0_6[506]},
      {stage1_6[174]}
   );
   gpc1_1 gpc2763 (
      {stage0_6[507]},
      {stage1_6[175]}
   );
   gpc1_1 gpc2764 (
      {stage0_6[508]},
      {stage1_6[176]}
   );
   gpc1_1 gpc2765 (
      {stage0_6[509]},
      {stage1_6[177]}
   );
   gpc1_1 gpc2766 (
      {stage0_6[510]},
      {stage1_6[178]}
   );
   gpc1_1 gpc2767 (
      {stage0_6[511]},
      {stage1_6[179]}
   );
   gpc1_1 gpc2768 (
      {stage0_7[364]},
      {stage1_7[192]}
   );
   gpc1_1 gpc2769 (
      {stage0_7[365]},
      {stage1_7[193]}
   );
   gpc1_1 gpc2770 (
      {stage0_7[366]},
      {stage1_7[194]}
   );
   gpc1_1 gpc2771 (
      {stage0_7[367]},
      {stage1_7[195]}
   );
   gpc1_1 gpc2772 (
      {stage0_7[368]},
      {stage1_7[196]}
   );
   gpc1_1 gpc2773 (
      {stage0_7[369]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2774 (
      {stage0_7[370]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2775 (
      {stage0_7[371]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2776 (
      {stage0_7[372]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2777 (
      {stage0_7[373]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2778 (
      {stage0_7[374]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2779 (
      {stage0_7[375]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2780 (
      {stage0_7[376]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2781 (
      {stage0_7[377]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2782 (
      {stage0_7[378]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2783 (
      {stage0_7[379]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2784 (
      {stage0_7[380]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2785 (
      {stage0_7[381]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2786 (
      {stage0_7[382]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2787 (
      {stage0_7[383]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2788 (
      {stage0_7[384]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2789 (
      {stage0_7[385]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2790 (
      {stage0_7[386]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2791 (
      {stage0_7[387]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2792 (
      {stage0_7[388]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2793 (
      {stage0_7[389]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2794 (
      {stage0_7[390]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2795 (
      {stage0_7[391]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2796 (
      {stage0_7[392]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2797 (
      {stage0_7[393]},
      {stage1_7[221]}
   );
   gpc1_1 gpc2798 (
      {stage0_7[394]},
      {stage1_7[222]}
   );
   gpc1_1 gpc2799 (
      {stage0_7[395]},
      {stage1_7[223]}
   );
   gpc1_1 gpc2800 (
      {stage0_7[396]},
      {stage1_7[224]}
   );
   gpc1_1 gpc2801 (
      {stage0_7[397]},
      {stage1_7[225]}
   );
   gpc1_1 gpc2802 (
      {stage0_7[398]},
      {stage1_7[226]}
   );
   gpc1_1 gpc2803 (
      {stage0_7[399]},
      {stage1_7[227]}
   );
   gpc1_1 gpc2804 (
      {stage0_7[400]},
      {stage1_7[228]}
   );
   gpc1_1 gpc2805 (
      {stage0_7[401]},
      {stage1_7[229]}
   );
   gpc1_1 gpc2806 (
      {stage0_7[402]},
      {stage1_7[230]}
   );
   gpc1_1 gpc2807 (
      {stage0_7[403]},
      {stage1_7[231]}
   );
   gpc1_1 gpc2808 (
      {stage0_7[404]},
      {stage1_7[232]}
   );
   gpc1_1 gpc2809 (
      {stage0_7[405]},
      {stage1_7[233]}
   );
   gpc1_1 gpc2810 (
      {stage0_7[406]},
      {stage1_7[234]}
   );
   gpc1_1 gpc2811 (
      {stage0_7[407]},
      {stage1_7[235]}
   );
   gpc1_1 gpc2812 (
      {stage0_7[408]},
      {stage1_7[236]}
   );
   gpc1_1 gpc2813 (
      {stage0_7[409]},
      {stage1_7[237]}
   );
   gpc1_1 gpc2814 (
      {stage0_7[410]},
      {stage1_7[238]}
   );
   gpc1_1 gpc2815 (
      {stage0_7[411]},
      {stage1_7[239]}
   );
   gpc1_1 gpc2816 (
      {stage0_7[412]},
      {stage1_7[240]}
   );
   gpc1_1 gpc2817 (
      {stage0_7[413]},
      {stage1_7[241]}
   );
   gpc1_1 gpc2818 (
      {stage0_7[414]},
      {stage1_7[242]}
   );
   gpc1_1 gpc2819 (
      {stage0_7[415]},
      {stage1_7[243]}
   );
   gpc1_1 gpc2820 (
      {stage0_7[416]},
      {stage1_7[244]}
   );
   gpc1_1 gpc2821 (
      {stage0_7[417]},
      {stage1_7[245]}
   );
   gpc1_1 gpc2822 (
      {stage0_7[418]},
      {stage1_7[246]}
   );
   gpc1_1 gpc2823 (
      {stage0_7[419]},
      {stage1_7[247]}
   );
   gpc1_1 gpc2824 (
      {stage0_7[420]},
      {stage1_7[248]}
   );
   gpc1_1 gpc2825 (
      {stage0_7[421]},
      {stage1_7[249]}
   );
   gpc1_1 gpc2826 (
      {stage0_7[422]},
      {stage1_7[250]}
   );
   gpc1_1 gpc2827 (
      {stage0_7[423]},
      {stage1_7[251]}
   );
   gpc1_1 gpc2828 (
      {stage0_7[424]},
      {stage1_7[252]}
   );
   gpc1_1 gpc2829 (
      {stage0_7[425]},
      {stage1_7[253]}
   );
   gpc1_1 gpc2830 (
      {stage0_7[426]},
      {stage1_7[254]}
   );
   gpc1_1 gpc2831 (
      {stage0_7[427]},
      {stage1_7[255]}
   );
   gpc1_1 gpc2832 (
      {stage0_7[428]},
      {stage1_7[256]}
   );
   gpc1_1 gpc2833 (
      {stage0_7[429]},
      {stage1_7[257]}
   );
   gpc1_1 gpc2834 (
      {stage0_7[430]},
      {stage1_7[258]}
   );
   gpc1_1 gpc2835 (
      {stage0_7[431]},
      {stage1_7[259]}
   );
   gpc1_1 gpc2836 (
      {stage0_7[432]},
      {stage1_7[260]}
   );
   gpc1_1 gpc2837 (
      {stage0_7[433]},
      {stage1_7[261]}
   );
   gpc1_1 gpc2838 (
      {stage0_7[434]},
      {stage1_7[262]}
   );
   gpc1_1 gpc2839 (
      {stage0_7[435]},
      {stage1_7[263]}
   );
   gpc1_1 gpc2840 (
      {stage0_7[436]},
      {stage1_7[264]}
   );
   gpc1_1 gpc2841 (
      {stage0_7[437]},
      {stage1_7[265]}
   );
   gpc1_1 gpc2842 (
      {stage0_7[438]},
      {stage1_7[266]}
   );
   gpc1_1 gpc2843 (
      {stage0_7[439]},
      {stage1_7[267]}
   );
   gpc1_1 gpc2844 (
      {stage0_7[440]},
      {stage1_7[268]}
   );
   gpc1_1 gpc2845 (
      {stage0_7[441]},
      {stage1_7[269]}
   );
   gpc1_1 gpc2846 (
      {stage0_7[442]},
      {stage1_7[270]}
   );
   gpc1_1 gpc2847 (
      {stage0_7[443]},
      {stage1_7[271]}
   );
   gpc1_1 gpc2848 (
      {stage0_7[444]},
      {stage1_7[272]}
   );
   gpc1_1 gpc2849 (
      {stage0_7[445]},
      {stage1_7[273]}
   );
   gpc1_1 gpc2850 (
      {stage0_7[446]},
      {stage1_7[274]}
   );
   gpc1_1 gpc2851 (
      {stage0_7[447]},
      {stage1_7[275]}
   );
   gpc1_1 gpc2852 (
      {stage0_7[448]},
      {stage1_7[276]}
   );
   gpc1_1 gpc2853 (
      {stage0_7[449]},
      {stage1_7[277]}
   );
   gpc1_1 gpc2854 (
      {stage0_7[450]},
      {stage1_7[278]}
   );
   gpc1_1 gpc2855 (
      {stage0_7[451]},
      {stage1_7[279]}
   );
   gpc1_1 gpc2856 (
      {stage0_7[452]},
      {stage1_7[280]}
   );
   gpc1_1 gpc2857 (
      {stage0_7[453]},
      {stage1_7[281]}
   );
   gpc1_1 gpc2858 (
      {stage0_7[454]},
      {stage1_7[282]}
   );
   gpc1_1 gpc2859 (
      {stage0_7[455]},
      {stage1_7[283]}
   );
   gpc1_1 gpc2860 (
      {stage0_7[456]},
      {stage1_7[284]}
   );
   gpc1_1 gpc2861 (
      {stage0_7[457]},
      {stage1_7[285]}
   );
   gpc1_1 gpc2862 (
      {stage0_7[458]},
      {stage1_7[286]}
   );
   gpc1_1 gpc2863 (
      {stage0_7[459]},
      {stage1_7[287]}
   );
   gpc1_1 gpc2864 (
      {stage0_7[460]},
      {stage1_7[288]}
   );
   gpc1_1 gpc2865 (
      {stage0_7[461]},
      {stage1_7[289]}
   );
   gpc1_1 gpc2866 (
      {stage0_7[462]},
      {stage1_7[290]}
   );
   gpc1_1 gpc2867 (
      {stage0_7[463]},
      {stage1_7[291]}
   );
   gpc1_1 gpc2868 (
      {stage0_7[464]},
      {stage1_7[292]}
   );
   gpc1_1 gpc2869 (
      {stage0_7[465]},
      {stage1_7[293]}
   );
   gpc1_1 gpc2870 (
      {stage0_7[466]},
      {stage1_7[294]}
   );
   gpc1_1 gpc2871 (
      {stage0_7[467]},
      {stage1_7[295]}
   );
   gpc1_1 gpc2872 (
      {stage0_7[468]},
      {stage1_7[296]}
   );
   gpc1_1 gpc2873 (
      {stage0_7[469]},
      {stage1_7[297]}
   );
   gpc1_1 gpc2874 (
      {stage0_7[470]},
      {stage1_7[298]}
   );
   gpc1_1 gpc2875 (
      {stage0_7[471]},
      {stage1_7[299]}
   );
   gpc1_1 gpc2876 (
      {stage0_7[472]},
      {stage1_7[300]}
   );
   gpc1_1 gpc2877 (
      {stage0_7[473]},
      {stage1_7[301]}
   );
   gpc1_1 gpc2878 (
      {stage0_7[474]},
      {stage1_7[302]}
   );
   gpc1_1 gpc2879 (
      {stage0_7[475]},
      {stage1_7[303]}
   );
   gpc1_1 gpc2880 (
      {stage0_7[476]},
      {stage1_7[304]}
   );
   gpc1_1 gpc2881 (
      {stage0_7[477]},
      {stage1_7[305]}
   );
   gpc1_1 gpc2882 (
      {stage0_7[478]},
      {stage1_7[306]}
   );
   gpc1_1 gpc2883 (
      {stage0_7[479]},
      {stage1_7[307]}
   );
   gpc1_1 gpc2884 (
      {stage0_7[480]},
      {stage1_7[308]}
   );
   gpc1_1 gpc2885 (
      {stage0_7[481]},
      {stage1_7[309]}
   );
   gpc1_1 gpc2886 (
      {stage0_7[482]},
      {stage1_7[310]}
   );
   gpc1_1 gpc2887 (
      {stage0_7[483]},
      {stage1_7[311]}
   );
   gpc1_1 gpc2888 (
      {stage0_7[484]},
      {stage1_7[312]}
   );
   gpc1_1 gpc2889 (
      {stage0_7[485]},
      {stage1_7[313]}
   );
   gpc1_1 gpc2890 (
      {stage0_7[486]},
      {stage1_7[314]}
   );
   gpc1_1 gpc2891 (
      {stage0_7[487]},
      {stage1_7[315]}
   );
   gpc1_1 gpc2892 (
      {stage0_7[488]},
      {stage1_7[316]}
   );
   gpc1_1 gpc2893 (
      {stage0_7[489]},
      {stage1_7[317]}
   );
   gpc1_1 gpc2894 (
      {stage0_7[490]},
      {stage1_7[318]}
   );
   gpc1_1 gpc2895 (
      {stage0_7[491]},
      {stage1_7[319]}
   );
   gpc1_1 gpc2896 (
      {stage0_7[492]},
      {stage1_7[320]}
   );
   gpc1_1 gpc2897 (
      {stage0_7[493]},
      {stage1_7[321]}
   );
   gpc1_1 gpc2898 (
      {stage0_7[494]},
      {stage1_7[322]}
   );
   gpc1_1 gpc2899 (
      {stage0_7[495]},
      {stage1_7[323]}
   );
   gpc1_1 gpc2900 (
      {stage0_7[496]},
      {stage1_7[324]}
   );
   gpc1_1 gpc2901 (
      {stage0_7[497]},
      {stage1_7[325]}
   );
   gpc1_1 gpc2902 (
      {stage0_7[498]},
      {stage1_7[326]}
   );
   gpc1_1 gpc2903 (
      {stage0_7[499]},
      {stage1_7[327]}
   );
   gpc1_1 gpc2904 (
      {stage0_7[500]},
      {stage1_7[328]}
   );
   gpc1_1 gpc2905 (
      {stage0_7[501]},
      {stage1_7[329]}
   );
   gpc1_1 gpc2906 (
      {stage0_7[502]},
      {stage1_7[330]}
   );
   gpc1_1 gpc2907 (
      {stage0_7[503]},
      {stage1_7[331]}
   );
   gpc1_1 gpc2908 (
      {stage0_7[504]},
      {stage1_7[332]}
   );
   gpc1_1 gpc2909 (
      {stage0_7[505]},
      {stage1_7[333]}
   );
   gpc1_1 gpc2910 (
      {stage0_7[506]},
      {stage1_7[334]}
   );
   gpc1_1 gpc2911 (
      {stage0_7[507]},
      {stage1_7[335]}
   );
   gpc1_1 gpc2912 (
      {stage0_7[508]},
      {stage1_7[336]}
   );
   gpc1_1 gpc2913 (
      {stage0_7[509]},
      {stage1_7[337]}
   );
   gpc1_1 gpc2914 (
      {stage0_7[510]},
      {stage1_7[338]}
   );
   gpc1_1 gpc2915 (
      {stage0_7[511]},
      {stage1_7[339]}
   );
   gpc1_1 gpc2916 (
      {stage0_8[493]},
      {stage1_8[220]}
   );
   gpc1_1 gpc2917 (
      {stage0_8[494]},
      {stage1_8[221]}
   );
   gpc1_1 gpc2918 (
      {stage0_8[495]},
      {stage1_8[222]}
   );
   gpc1_1 gpc2919 (
      {stage0_8[496]},
      {stage1_8[223]}
   );
   gpc1_1 gpc2920 (
      {stage0_8[497]},
      {stage1_8[224]}
   );
   gpc1_1 gpc2921 (
      {stage0_8[498]},
      {stage1_8[225]}
   );
   gpc1_1 gpc2922 (
      {stage0_8[499]},
      {stage1_8[226]}
   );
   gpc1_1 gpc2923 (
      {stage0_8[500]},
      {stage1_8[227]}
   );
   gpc1_1 gpc2924 (
      {stage0_8[501]},
      {stage1_8[228]}
   );
   gpc1_1 gpc2925 (
      {stage0_8[502]},
      {stage1_8[229]}
   );
   gpc1_1 gpc2926 (
      {stage0_8[503]},
      {stage1_8[230]}
   );
   gpc1_1 gpc2927 (
      {stage0_8[504]},
      {stage1_8[231]}
   );
   gpc1_1 gpc2928 (
      {stage0_8[505]},
      {stage1_8[232]}
   );
   gpc1_1 gpc2929 (
      {stage0_8[506]},
      {stage1_8[233]}
   );
   gpc1_1 gpc2930 (
      {stage0_8[507]},
      {stage1_8[234]}
   );
   gpc1_1 gpc2931 (
      {stage0_8[508]},
      {stage1_8[235]}
   );
   gpc1_1 gpc2932 (
      {stage0_8[509]},
      {stage1_8[236]}
   );
   gpc1_1 gpc2933 (
      {stage0_8[510]},
      {stage1_8[237]}
   );
   gpc1_1 gpc2934 (
      {stage0_8[511]},
      {stage1_8[238]}
   );
   gpc1_1 gpc2935 (
      {stage0_9[312]},
      {stage1_9[163]}
   );
   gpc1_1 gpc2936 (
      {stage0_9[313]},
      {stage1_9[164]}
   );
   gpc1_1 gpc2937 (
      {stage0_9[314]},
      {stage1_9[165]}
   );
   gpc1_1 gpc2938 (
      {stage0_9[315]},
      {stage1_9[166]}
   );
   gpc1_1 gpc2939 (
      {stage0_9[316]},
      {stage1_9[167]}
   );
   gpc1_1 gpc2940 (
      {stage0_9[317]},
      {stage1_9[168]}
   );
   gpc1_1 gpc2941 (
      {stage0_9[318]},
      {stage1_9[169]}
   );
   gpc1_1 gpc2942 (
      {stage0_9[319]},
      {stage1_9[170]}
   );
   gpc1_1 gpc2943 (
      {stage0_9[320]},
      {stage1_9[171]}
   );
   gpc1_1 gpc2944 (
      {stage0_9[321]},
      {stage1_9[172]}
   );
   gpc1_1 gpc2945 (
      {stage0_9[322]},
      {stage1_9[173]}
   );
   gpc1_1 gpc2946 (
      {stage0_9[323]},
      {stage1_9[174]}
   );
   gpc1_1 gpc2947 (
      {stage0_9[324]},
      {stage1_9[175]}
   );
   gpc1_1 gpc2948 (
      {stage0_9[325]},
      {stage1_9[176]}
   );
   gpc1_1 gpc2949 (
      {stage0_9[326]},
      {stage1_9[177]}
   );
   gpc1_1 gpc2950 (
      {stage0_9[327]},
      {stage1_9[178]}
   );
   gpc1_1 gpc2951 (
      {stage0_9[328]},
      {stage1_9[179]}
   );
   gpc1_1 gpc2952 (
      {stage0_9[329]},
      {stage1_9[180]}
   );
   gpc1_1 gpc2953 (
      {stage0_9[330]},
      {stage1_9[181]}
   );
   gpc1_1 gpc2954 (
      {stage0_9[331]},
      {stage1_9[182]}
   );
   gpc1_1 gpc2955 (
      {stage0_9[332]},
      {stage1_9[183]}
   );
   gpc1_1 gpc2956 (
      {stage0_9[333]},
      {stage1_9[184]}
   );
   gpc1_1 gpc2957 (
      {stage0_9[334]},
      {stage1_9[185]}
   );
   gpc1_1 gpc2958 (
      {stage0_9[335]},
      {stage1_9[186]}
   );
   gpc1_1 gpc2959 (
      {stage0_9[336]},
      {stage1_9[187]}
   );
   gpc1_1 gpc2960 (
      {stage0_9[337]},
      {stage1_9[188]}
   );
   gpc1_1 gpc2961 (
      {stage0_9[338]},
      {stage1_9[189]}
   );
   gpc1_1 gpc2962 (
      {stage0_9[339]},
      {stage1_9[190]}
   );
   gpc1_1 gpc2963 (
      {stage0_9[340]},
      {stage1_9[191]}
   );
   gpc1_1 gpc2964 (
      {stage0_9[341]},
      {stage1_9[192]}
   );
   gpc1_1 gpc2965 (
      {stage0_9[342]},
      {stage1_9[193]}
   );
   gpc1_1 gpc2966 (
      {stage0_9[343]},
      {stage1_9[194]}
   );
   gpc1_1 gpc2967 (
      {stage0_9[344]},
      {stage1_9[195]}
   );
   gpc1_1 gpc2968 (
      {stage0_9[345]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2969 (
      {stage0_9[346]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2970 (
      {stage0_9[347]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2971 (
      {stage0_9[348]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2972 (
      {stage0_9[349]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2973 (
      {stage0_9[350]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2974 (
      {stage0_9[351]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2975 (
      {stage0_9[352]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2976 (
      {stage0_9[353]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2977 (
      {stage0_9[354]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2978 (
      {stage0_9[355]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2979 (
      {stage0_9[356]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2980 (
      {stage0_9[357]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2981 (
      {stage0_9[358]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2982 (
      {stage0_9[359]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2983 (
      {stage0_9[360]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2984 (
      {stage0_9[361]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2985 (
      {stage0_9[362]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2986 (
      {stage0_9[363]},
      {stage1_9[214]}
   );
   gpc1_1 gpc2987 (
      {stage0_9[364]},
      {stage1_9[215]}
   );
   gpc1_1 gpc2988 (
      {stage0_9[365]},
      {stage1_9[216]}
   );
   gpc1_1 gpc2989 (
      {stage0_9[366]},
      {stage1_9[217]}
   );
   gpc1_1 gpc2990 (
      {stage0_9[367]},
      {stage1_9[218]}
   );
   gpc1_1 gpc2991 (
      {stage0_9[368]},
      {stage1_9[219]}
   );
   gpc1_1 gpc2992 (
      {stage0_9[369]},
      {stage1_9[220]}
   );
   gpc1_1 gpc2993 (
      {stage0_9[370]},
      {stage1_9[221]}
   );
   gpc1_1 gpc2994 (
      {stage0_9[371]},
      {stage1_9[222]}
   );
   gpc1_1 gpc2995 (
      {stage0_9[372]},
      {stage1_9[223]}
   );
   gpc1_1 gpc2996 (
      {stage0_9[373]},
      {stage1_9[224]}
   );
   gpc1_1 gpc2997 (
      {stage0_9[374]},
      {stage1_9[225]}
   );
   gpc1_1 gpc2998 (
      {stage0_9[375]},
      {stage1_9[226]}
   );
   gpc1_1 gpc2999 (
      {stage0_9[376]},
      {stage1_9[227]}
   );
   gpc1_1 gpc3000 (
      {stage0_9[377]},
      {stage1_9[228]}
   );
   gpc1_1 gpc3001 (
      {stage0_9[378]},
      {stage1_9[229]}
   );
   gpc1_1 gpc3002 (
      {stage0_9[379]},
      {stage1_9[230]}
   );
   gpc1_1 gpc3003 (
      {stage0_9[380]},
      {stage1_9[231]}
   );
   gpc1_1 gpc3004 (
      {stage0_9[381]},
      {stage1_9[232]}
   );
   gpc1_1 gpc3005 (
      {stage0_9[382]},
      {stage1_9[233]}
   );
   gpc1_1 gpc3006 (
      {stage0_9[383]},
      {stage1_9[234]}
   );
   gpc1_1 gpc3007 (
      {stage0_9[384]},
      {stage1_9[235]}
   );
   gpc1_1 gpc3008 (
      {stage0_9[385]},
      {stage1_9[236]}
   );
   gpc1_1 gpc3009 (
      {stage0_9[386]},
      {stage1_9[237]}
   );
   gpc1_1 gpc3010 (
      {stage0_9[387]},
      {stage1_9[238]}
   );
   gpc1_1 gpc3011 (
      {stage0_9[388]},
      {stage1_9[239]}
   );
   gpc1_1 gpc3012 (
      {stage0_9[389]},
      {stage1_9[240]}
   );
   gpc1_1 gpc3013 (
      {stage0_9[390]},
      {stage1_9[241]}
   );
   gpc1_1 gpc3014 (
      {stage0_9[391]},
      {stage1_9[242]}
   );
   gpc1_1 gpc3015 (
      {stage0_9[392]},
      {stage1_9[243]}
   );
   gpc1_1 gpc3016 (
      {stage0_9[393]},
      {stage1_9[244]}
   );
   gpc1_1 gpc3017 (
      {stage0_9[394]},
      {stage1_9[245]}
   );
   gpc1_1 gpc3018 (
      {stage0_9[395]},
      {stage1_9[246]}
   );
   gpc1_1 gpc3019 (
      {stage0_9[396]},
      {stage1_9[247]}
   );
   gpc1_1 gpc3020 (
      {stage0_9[397]},
      {stage1_9[248]}
   );
   gpc1_1 gpc3021 (
      {stage0_9[398]},
      {stage1_9[249]}
   );
   gpc1_1 gpc3022 (
      {stage0_9[399]},
      {stage1_9[250]}
   );
   gpc1_1 gpc3023 (
      {stage0_9[400]},
      {stage1_9[251]}
   );
   gpc1_1 gpc3024 (
      {stage0_9[401]},
      {stage1_9[252]}
   );
   gpc1_1 gpc3025 (
      {stage0_9[402]},
      {stage1_9[253]}
   );
   gpc1_1 gpc3026 (
      {stage0_9[403]},
      {stage1_9[254]}
   );
   gpc1_1 gpc3027 (
      {stage0_9[404]},
      {stage1_9[255]}
   );
   gpc1_1 gpc3028 (
      {stage0_9[405]},
      {stage1_9[256]}
   );
   gpc1_1 gpc3029 (
      {stage0_9[406]},
      {stage1_9[257]}
   );
   gpc1_1 gpc3030 (
      {stage0_9[407]},
      {stage1_9[258]}
   );
   gpc1_1 gpc3031 (
      {stage0_9[408]},
      {stage1_9[259]}
   );
   gpc1_1 gpc3032 (
      {stage0_9[409]},
      {stage1_9[260]}
   );
   gpc1_1 gpc3033 (
      {stage0_9[410]},
      {stage1_9[261]}
   );
   gpc1_1 gpc3034 (
      {stage0_9[411]},
      {stage1_9[262]}
   );
   gpc1_1 gpc3035 (
      {stage0_9[412]},
      {stage1_9[263]}
   );
   gpc1_1 gpc3036 (
      {stage0_9[413]},
      {stage1_9[264]}
   );
   gpc1_1 gpc3037 (
      {stage0_9[414]},
      {stage1_9[265]}
   );
   gpc1_1 gpc3038 (
      {stage0_9[415]},
      {stage1_9[266]}
   );
   gpc1_1 gpc3039 (
      {stage0_9[416]},
      {stage1_9[267]}
   );
   gpc1_1 gpc3040 (
      {stage0_9[417]},
      {stage1_9[268]}
   );
   gpc1_1 gpc3041 (
      {stage0_9[418]},
      {stage1_9[269]}
   );
   gpc1_1 gpc3042 (
      {stage0_9[419]},
      {stage1_9[270]}
   );
   gpc1_1 gpc3043 (
      {stage0_9[420]},
      {stage1_9[271]}
   );
   gpc1_1 gpc3044 (
      {stage0_9[421]},
      {stage1_9[272]}
   );
   gpc1_1 gpc3045 (
      {stage0_9[422]},
      {stage1_9[273]}
   );
   gpc1_1 gpc3046 (
      {stage0_9[423]},
      {stage1_9[274]}
   );
   gpc1_1 gpc3047 (
      {stage0_9[424]},
      {stage1_9[275]}
   );
   gpc1_1 gpc3048 (
      {stage0_9[425]},
      {stage1_9[276]}
   );
   gpc1_1 gpc3049 (
      {stage0_9[426]},
      {stage1_9[277]}
   );
   gpc1_1 gpc3050 (
      {stage0_9[427]},
      {stage1_9[278]}
   );
   gpc1_1 gpc3051 (
      {stage0_9[428]},
      {stage1_9[279]}
   );
   gpc1_1 gpc3052 (
      {stage0_9[429]},
      {stage1_9[280]}
   );
   gpc1_1 gpc3053 (
      {stage0_9[430]},
      {stage1_9[281]}
   );
   gpc1_1 gpc3054 (
      {stage0_9[431]},
      {stage1_9[282]}
   );
   gpc1_1 gpc3055 (
      {stage0_9[432]},
      {stage1_9[283]}
   );
   gpc1_1 gpc3056 (
      {stage0_9[433]},
      {stage1_9[284]}
   );
   gpc1_1 gpc3057 (
      {stage0_9[434]},
      {stage1_9[285]}
   );
   gpc1_1 gpc3058 (
      {stage0_9[435]},
      {stage1_9[286]}
   );
   gpc1_1 gpc3059 (
      {stage0_9[436]},
      {stage1_9[287]}
   );
   gpc1_1 gpc3060 (
      {stage0_9[437]},
      {stage1_9[288]}
   );
   gpc1_1 gpc3061 (
      {stage0_9[438]},
      {stage1_9[289]}
   );
   gpc1_1 gpc3062 (
      {stage0_9[439]},
      {stage1_9[290]}
   );
   gpc1_1 gpc3063 (
      {stage0_9[440]},
      {stage1_9[291]}
   );
   gpc1_1 gpc3064 (
      {stage0_9[441]},
      {stage1_9[292]}
   );
   gpc1_1 gpc3065 (
      {stage0_9[442]},
      {stage1_9[293]}
   );
   gpc1_1 gpc3066 (
      {stage0_9[443]},
      {stage1_9[294]}
   );
   gpc1_1 gpc3067 (
      {stage0_9[444]},
      {stage1_9[295]}
   );
   gpc1_1 gpc3068 (
      {stage0_9[445]},
      {stage1_9[296]}
   );
   gpc1_1 gpc3069 (
      {stage0_9[446]},
      {stage1_9[297]}
   );
   gpc1_1 gpc3070 (
      {stage0_9[447]},
      {stage1_9[298]}
   );
   gpc1_1 gpc3071 (
      {stage0_9[448]},
      {stage1_9[299]}
   );
   gpc1_1 gpc3072 (
      {stage0_9[449]},
      {stage1_9[300]}
   );
   gpc1_1 gpc3073 (
      {stage0_9[450]},
      {stage1_9[301]}
   );
   gpc1_1 gpc3074 (
      {stage0_9[451]},
      {stage1_9[302]}
   );
   gpc1_1 gpc3075 (
      {stage0_9[452]},
      {stage1_9[303]}
   );
   gpc1_1 gpc3076 (
      {stage0_9[453]},
      {stage1_9[304]}
   );
   gpc1_1 gpc3077 (
      {stage0_9[454]},
      {stage1_9[305]}
   );
   gpc1_1 gpc3078 (
      {stage0_9[455]},
      {stage1_9[306]}
   );
   gpc1_1 gpc3079 (
      {stage0_9[456]},
      {stage1_9[307]}
   );
   gpc1_1 gpc3080 (
      {stage0_9[457]},
      {stage1_9[308]}
   );
   gpc1_1 gpc3081 (
      {stage0_9[458]},
      {stage1_9[309]}
   );
   gpc1_1 gpc3082 (
      {stage0_9[459]},
      {stage1_9[310]}
   );
   gpc1_1 gpc3083 (
      {stage0_9[460]},
      {stage1_9[311]}
   );
   gpc1_1 gpc3084 (
      {stage0_9[461]},
      {stage1_9[312]}
   );
   gpc1_1 gpc3085 (
      {stage0_9[462]},
      {stage1_9[313]}
   );
   gpc1_1 gpc3086 (
      {stage0_9[463]},
      {stage1_9[314]}
   );
   gpc1_1 gpc3087 (
      {stage0_9[464]},
      {stage1_9[315]}
   );
   gpc1_1 gpc3088 (
      {stage0_9[465]},
      {stage1_9[316]}
   );
   gpc1_1 gpc3089 (
      {stage0_9[466]},
      {stage1_9[317]}
   );
   gpc1_1 gpc3090 (
      {stage0_9[467]},
      {stage1_9[318]}
   );
   gpc1_1 gpc3091 (
      {stage0_9[468]},
      {stage1_9[319]}
   );
   gpc1_1 gpc3092 (
      {stage0_9[469]},
      {stage1_9[320]}
   );
   gpc1_1 gpc3093 (
      {stage0_9[470]},
      {stage1_9[321]}
   );
   gpc1_1 gpc3094 (
      {stage0_9[471]},
      {stage1_9[322]}
   );
   gpc1_1 gpc3095 (
      {stage0_9[472]},
      {stage1_9[323]}
   );
   gpc1_1 gpc3096 (
      {stage0_9[473]},
      {stage1_9[324]}
   );
   gpc1_1 gpc3097 (
      {stage0_9[474]},
      {stage1_9[325]}
   );
   gpc1_1 gpc3098 (
      {stage0_9[475]},
      {stage1_9[326]}
   );
   gpc1_1 gpc3099 (
      {stage0_9[476]},
      {stage1_9[327]}
   );
   gpc1_1 gpc3100 (
      {stage0_9[477]},
      {stage1_9[328]}
   );
   gpc1_1 gpc3101 (
      {stage0_9[478]},
      {stage1_9[329]}
   );
   gpc1_1 gpc3102 (
      {stage0_9[479]},
      {stage1_9[330]}
   );
   gpc1_1 gpc3103 (
      {stage0_9[480]},
      {stage1_9[331]}
   );
   gpc1_1 gpc3104 (
      {stage0_9[481]},
      {stage1_9[332]}
   );
   gpc1_1 gpc3105 (
      {stage0_9[482]},
      {stage1_9[333]}
   );
   gpc1_1 gpc3106 (
      {stage0_9[483]},
      {stage1_9[334]}
   );
   gpc1_1 gpc3107 (
      {stage0_9[484]},
      {stage1_9[335]}
   );
   gpc1_1 gpc3108 (
      {stage0_9[485]},
      {stage1_9[336]}
   );
   gpc1_1 gpc3109 (
      {stage0_9[486]},
      {stage1_9[337]}
   );
   gpc1_1 gpc3110 (
      {stage0_9[487]},
      {stage1_9[338]}
   );
   gpc1_1 gpc3111 (
      {stage0_9[488]},
      {stage1_9[339]}
   );
   gpc1_1 gpc3112 (
      {stage0_9[489]},
      {stage1_9[340]}
   );
   gpc1_1 gpc3113 (
      {stage0_9[490]},
      {stage1_9[341]}
   );
   gpc1_1 gpc3114 (
      {stage0_9[491]},
      {stage1_9[342]}
   );
   gpc1_1 gpc3115 (
      {stage0_9[492]},
      {stage1_9[343]}
   );
   gpc1_1 gpc3116 (
      {stage0_9[493]},
      {stage1_9[344]}
   );
   gpc1_1 gpc3117 (
      {stage0_9[494]},
      {stage1_9[345]}
   );
   gpc1_1 gpc3118 (
      {stage0_9[495]},
      {stage1_9[346]}
   );
   gpc1_1 gpc3119 (
      {stage0_9[496]},
      {stage1_9[347]}
   );
   gpc1_1 gpc3120 (
      {stage0_9[497]},
      {stage1_9[348]}
   );
   gpc1_1 gpc3121 (
      {stage0_9[498]},
      {stage1_9[349]}
   );
   gpc1_1 gpc3122 (
      {stage0_9[499]},
      {stage1_9[350]}
   );
   gpc1_1 gpc3123 (
      {stage0_9[500]},
      {stage1_9[351]}
   );
   gpc1_1 gpc3124 (
      {stage0_9[501]},
      {stage1_9[352]}
   );
   gpc1_1 gpc3125 (
      {stage0_9[502]},
      {stage1_9[353]}
   );
   gpc1_1 gpc3126 (
      {stage0_9[503]},
      {stage1_9[354]}
   );
   gpc1_1 gpc3127 (
      {stage0_9[504]},
      {stage1_9[355]}
   );
   gpc1_1 gpc3128 (
      {stage0_9[505]},
      {stage1_9[356]}
   );
   gpc1_1 gpc3129 (
      {stage0_9[506]},
      {stage1_9[357]}
   );
   gpc1_1 gpc3130 (
      {stage0_9[507]},
      {stage1_9[358]}
   );
   gpc1_1 gpc3131 (
      {stage0_9[508]},
      {stage1_9[359]}
   );
   gpc1_1 gpc3132 (
      {stage0_9[509]},
      {stage1_9[360]}
   );
   gpc1_1 gpc3133 (
      {stage0_9[510]},
      {stage1_9[361]}
   );
   gpc1_1 gpc3134 (
      {stage0_9[511]},
      {stage1_9[362]}
   );
   gpc1_1 gpc3135 (
      {stage0_10[502]},
      {stage1_10[143]}
   );
   gpc1_1 gpc3136 (
      {stage0_10[503]},
      {stage1_10[144]}
   );
   gpc1_1 gpc3137 (
      {stage0_10[504]},
      {stage1_10[145]}
   );
   gpc1_1 gpc3138 (
      {stage0_10[505]},
      {stage1_10[146]}
   );
   gpc1_1 gpc3139 (
      {stage0_10[506]},
      {stage1_10[147]}
   );
   gpc1_1 gpc3140 (
      {stage0_10[507]},
      {stage1_10[148]}
   );
   gpc1_1 gpc3141 (
      {stage0_10[508]},
      {stage1_10[149]}
   );
   gpc1_1 gpc3142 (
      {stage0_10[509]},
      {stage1_10[150]}
   );
   gpc1_1 gpc3143 (
      {stage0_10[510]},
      {stage1_10[151]}
   );
   gpc1_1 gpc3144 (
      {stage0_10[511]},
      {stage1_10[152]}
   );
   gpc1_1 gpc3145 (
      {stage0_11[380]},
      {stage1_11[186]}
   );
   gpc1_1 gpc3146 (
      {stage0_11[381]},
      {stage1_11[187]}
   );
   gpc1_1 gpc3147 (
      {stage0_11[382]},
      {stage1_11[188]}
   );
   gpc1_1 gpc3148 (
      {stage0_11[383]},
      {stage1_11[189]}
   );
   gpc1_1 gpc3149 (
      {stage0_11[384]},
      {stage1_11[190]}
   );
   gpc1_1 gpc3150 (
      {stage0_11[385]},
      {stage1_11[191]}
   );
   gpc1_1 gpc3151 (
      {stage0_11[386]},
      {stage1_11[192]}
   );
   gpc1_1 gpc3152 (
      {stage0_11[387]},
      {stage1_11[193]}
   );
   gpc1_1 gpc3153 (
      {stage0_11[388]},
      {stage1_11[194]}
   );
   gpc1_1 gpc3154 (
      {stage0_11[389]},
      {stage1_11[195]}
   );
   gpc1_1 gpc3155 (
      {stage0_11[390]},
      {stage1_11[196]}
   );
   gpc1_1 gpc3156 (
      {stage0_11[391]},
      {stage1_11[197]}
   );
   gpc1_1 gpc3157 (
      {stage0_11[392]},
      {stage1_11[198]}
   );
   gpc1_1 gpc3158 (
      {stage0_11[393]},
      {stage1_11[199]}
   );
   gpc1_1 gpc3159 (
      {stage0_11[394]},
      {stage1_11[200]}
   );
   gpc1_1 gpc3160 (
      {stage0_11[395]},
      {stage1_11[201]}
   );
   gpc1_1 gpc3161 (
      {stage0_11[396]},
      {stage1_11[202]}
   );
   gpc1_1 gpc3162 (
      {stage0_11[397]},
      {stage1_11[203]}
   );
   gpc1_1 gpc3163 (
      {stage0_11[398]},
      {stage1_11[204]}
   );
   gpc1_1 gpc3164 (
      {stage0_11[399]},
      {stage1_11[205]}
   );
   gpc1_1 gpc3165 (
      {stage0_11[400]},
      {stage1_11[206]}
   );
   gpc1_1 gpc3166 (
      {stage0_11[401]},
      {stage1_11[207]}
   );
   gpc1_1 gpc3167 (
      {stage0_11[402]},
      {stage1_11[208]}
   );
   gpc1_1 gpc3168 (
      {stage0_11[403]},
      {stage1_11[209]}
   );
   gpc1_1 gpc3169 (
      {stage0_11[404]},
      {stage1_11[210]}
   );
   gpc1_1 gpc3170 (
      {stage0_11[405]},
      {stage1_11[211]}
   );
   gpc1_1 gpc3171 (
      {stage0_11[406]},
      {stage1_11[212]}
   );
   gpc1_1 gpc3172 (
      {stage0_11[407]},
      {stage1_11[213]}
   );
   gpc1_1 gpc3173 (
      {stage0_11[408]},
      {stage1_11[214]}
   );
   gpc1_1 gpc3174 (
      {stage0_11[409]},
      {stage1_11[215]}
   );
   gpc1_1 gpc3175 (
      {stage0_11[410]},
      {stage1_11[216]}
   );
   gpc1_1 gpc3176 (
      {stage0_11[411]},
      {stage1_11[217]}
   );
   gpc1_1 gpc3177 (
      {stage0_11[412]},
      {stage1_11[218]}
   );
   gpc1_1 gpc3178 (
      {stage0_11[413]},
      {stage1_11[219]}
   );
   gpc1_1 gpc3179 (
      {stage0_11[414]},
      {stage1_11[220]}
   );
   gpc1_1 gpc3180 (
      {stage0_11[415]},
      {stage1_11[221]}
   );
   gpc1_1 gpc3181 (
      {stage0_11[416]},
      {stage1_11[222]}
   );
   gpc1_1 gpc3182 (
      {stage0_11[417]},
      {stage1_11[223]}
   );
   gpc1_1 gpc3183 (
      {stage0_11[418]},
      {stage1_11[224]}
   );
   gpc1_1 gpc3184 (
      {stage0_11[419]},
      {stage1_11[225]}
   );
   gpc1_1 gpc3185 (
      {stage0_11[420]},
      {stage1_11[226]}
   );
   gpc1_1 gpc3186 (
      {stage0_11[421]},
      {stage1_11[227]}
   );
   gpc1_1 gpc3187 (
      {stage0_11[422]},
      {stage1_11[228]}
   );
   gpc1_1 gpc3188 (
      {stage0_11[423]},
      {stage1_11[229]}
   );
   gpc1_1 gpc3189 (
      {stage0_11[424]},
      {stage1_11[230]}
   );
   gpc1_1 gpc3190 (
      {stage0_11[425]},
      {stage1_11[231]}
   );
   gpc1_1 gpc3191 (
      {stage0_11[426]},
      {stage1_11[232]}
   );
   gpc1_1 gpc3192 (
      {stage0_11[427]},
      {stage1_11[233]}
   );
   gpc1_1 gpc3193 (
      {stage0_11[428]},
      {stage1_11[234]}
   );
   gpc1_1 gpc3194 (
      {stage0_11[429]},
      {stage1_11[235]}
   );
   gpc1_1 gpc3195 (
      {stage0_11[430]},
      {stage1_11[236]}
   );
   gpc1_1 gpc3196 (
      {stage0_11[431]},
      {stage1_11[237]}
   );
   gpc1_1 gpc3197 (
      {stage0_11[432]},
      {stage1_11[238]}
   );
   gpc1_1 gpc3198 (
      {stage0_11[433]},
      {stage1_11[239]}
   );
   gpc1_1 gpc3199 (
      {stage0_11[434]},
      {stage1_11[240]}
   );
   gpc1_1 gpc3200 (
      {stage0_11[435]},
      {stage1_11[241]}
   );
   gpc1_1 gpc3201 (
      {stage0_11[436]},
      {stage1_11[242]}
   );
   gpc1_1 gpc3202 (
      {stage0_11[437]},
      {stage1_11[243]}
   );
   gpc1_1 gpc3203 (
      {stage0_11[438]},
      {stage1_11[244]}
   );
   gpc1_1 gpc3204 (
      {stage0_11[439]},
      {stage1_11[245]}
   );
   gpc1_1 gpc3205 (
      {stage0_11[440]},
      {stage1_11[246]}
   );
   gpc1_1 gpc3206 (
      {stage0_11[441]},
      {stage1_11[247]}
   );
   gpc1_1 gpc3207 (
      {stage0_11[442]},
      {stage1_11[248]}
   );
   gpc1_1 gpc3208 (
      {stage0_11[443]},
      {stage1_11[249]}
   );
   gpc1_1 gpc3209 (
      {stage0_11[444]},
      {stage1_11[250]}
   );
   gpc1_1 gpc3210 (
      {stage0_11[445]},
      {stage1_11[251]}
   );
   gpc1_1 gpc3211 (
      {stage0_11[446]},
      {stage1_11[252]}
   );
   gpc1_1 gpc3212 (
      {stage0_11[447]},
      {stage1_11[253]}
   );
   gpc1_1 gpc3213 (
      {stage0_11[448]},
      {stage1_11[254]}
   );
   gpc1_1 gpc3214 (
      {stage0_11[449]},
      {stage1_11[255]}
   );
   gpc1_1 gpc3215 (
      {stage0_11[450]},
      {stage1_11[256]}
   );
   gpc1_1 gpc3216 (
      {stage0_11[451]},
      {stage1_11[257]}
   );
   gpc1_1 gpc3217 (
      {stage0_11[452]},
      {stage1_11[258]}
   );
   gpc1_1 gpc3218 (
      {stage0_11[453]},
      {stage1_11[259]}
   );
   gpc1_1 gpc3219 (
      {stage0_11[454]},
      {stage1_11[260]}
   );
   gpc1_1 gpc3220 (
      {stage0_11[455]},
      {stage1_11[261]}
   );
   gpc1_1 gpc3221 (
      {stage0_11[456]},
      {stage1_11[262]}
   );
   gpc1_1 gpc3222 (
      {stage0_11[457]},
      {stage1_11[263]}
   );
   gpc1_1 gpc3223 (
      {stage0_11[458]},
      {stage1_11[264]}
   );
   gpc1_1 gpc3224 (
      {stage0_11[459]},
      {stage1_11[265]}
   );
   gpc1_1 gpc3225 (
      {stage0_11[460]},
      {stage1_11[266]}
   );
   gpc1_1 gpc3226 (
      {stage0_11[461]},
      {stage1_11[267]}
   );
   gpc1_1 gpc3227 (
      {stage0_11[462]},
      {stage1_11[268]}
   );
   gpc1_1 gpc3228 (
      {stage0_11[463]},
      {stage1_11[269]}
   );
   gpc1_1 gpc3229 (
      {stage0_11[464]},
      {stage1_11[270]}
   );
   gpc1_1 gpc3230 (
      {stage0_11[465]},
      {stage1_11[271]}
   );
   gpc1_1 gpc3231 (
      {stage0_11[466]},
      {stage1_11[272]}
   );
   gpc1_1 gpc3232 (
      {stage0_11[467]},
      {stage1_11[273]}
   );
   gpc1_1 gpc3233 (
      {stage0_11[468]},
      {stage1_11[274]}
   );
   gpc1_1 gpc3234 (
      {stage0_11[469]},
      {stage1_11[275]}
   );
   gpc1_1 gpc3235 (
      {stage0_11[470]},
      {stage1_11[276]}
   );
   gpc1_1 gpc3236 (
      {stage0_11[471]},
      {stage1_11[277]}
   );
   gpc1_1 gpc3237 (
      {stage0_11[472]},
      {stage1_11[278]}
   );
   gpc1_1 gpc3238 (
      {stage0_11[473]},
      {stage1_11[279]}
   );
   gpc1_1 gpc3239 (
      {stage0_11[474]},
      {stage1_11[280]}
   );
   gpc1_1 gpc3240 (
      {stage0_11[475]},
      {stage1_11[281]}
   );
   gpc1_1 gpc3241 (
      {stage0_11[476]},
      {stage1_11[282]}
   );
   gpc1_1 gpc3242 (
      {stage0_11[477]},
      {stage1_11[283]}
   );
   gpc1_1 gpc3243 (
      {stage0_11[478]},
      {stage1_11[284]}
   );
   gpc1_1 gpc3244 (
      {stage0_11[479]},
      {stage1_11[285]}
   );
   gpc1_1 gpc3245 (
      {stage0_11[480]},
      {stage1_11[286]}
   );
   gpc1_1 gpc3246 (
      {stage0_11[481]},
      {stage1_11[287]}
   );
   gpc1_1 gpc3247 (
      {stage0_11[482]},
      {stage1_11[288]}
   );
   gpc1_1 gpc3248 (
      {stage0_11[483]},
      {stage1_11[289]}
   );
   gpc1_1 gpc3249 (
      {stage0_11[484]},
      {stage1_11[290]}
   );
   gpc1_1 gpc3250 (
      {stage0_11[485]},
      {stage1_11[291]}
   );
   gpc1_1 gpc3251 (
      {stage0_11[486]},
      {stage1_11[292]}
   );
   gpc1_1 gpc3252 (
      {stage0_11[487]},
      {stage1_11[293]}
   );
   gpc1_1 gpc3253 (
      {stage0_11[488]},
      {stage1_11[294]}
   );
   gpc1_1 gpc3254 (
      {stage0_11[489]},
      {stage1_11[295]}
   );
   gpc1_1 gpc3255 (
      {stage0_11[490]},
      {stage1_11[296]}
   );
   gpc1_1 gpc3256 (
      {stage0_11[491]},
      {stage1_11[297]}
   );
   gpc1_1 gpc3257 (
      {stage0_11[492]},
      {stage1_11[298]}
   );
   gpc1_1 gpc3258 (
      {stage0_11[493]},
      {stage1_11[299]}
   );
   gpc1_1 gpc3259 (
      {stage0_11[494]},
      {stage1_11[300]}
   );
   gpc1_1 gpc3260 (
      {stage0_11[495]},
      {stage1_11[301]}
   );
   gpc1_1 gpc3261 (
      {stage0_11[496]},
      {stage1_11[302]}
   );
   gpc1_1 gpc3262 (
      {stage0_11[497]},
      {stage1_11[303]}
   );
   gpc1_1 gpc3263 (
      {stage0_11[498]},
      {stage1_11[304]}
   );
   gpc1_1 gpc3264 (
      {stage0_11[499]},
      {stage1_11[305]}
   );
   gpc1_1 gpc3265 (
      {stage0_11[500]},
      {stage1_11[306]}
   );
   gpc1_1 gpc3266 (
      {stage0_11[501]},
      {stage1_11[307]}
   );
   gpc1_1 gpc3267 (
      {stage0_11[502]},
      {stage1_11[308]}
   );
   gpc1_1 gpc3268 (
      {stage0_11[503]},
      {stage1_11[309]}
   );
   gpc1_1 gpc3269 (
      {stage0_11[504]},
      {stage1_11[310]}
   );
   gpc1_1 gpc3270 (
      {stage0_11[505]},
      {stage1_11[311]}
   );
   gpc1_1 gpc3271 (
      {stage0_11[506]},
      {stage1_11[312]}
   );
   gpc1_1 gpc3272 (
      {stage0_11[507]},
      {stage1_11[313]}
   );
   gpc1_1 gpc3273 (
      {stage0_11[508]},
      {stage1_11[314]}
   );
   gpc1_1 gpc3274 (
      {stage0_11[509]},
      {stage1_11[315]}
   );
   gpc1_1 gpc3275 (
      {stage0_11[510]},
      {stage1_11[316]}
   );
   gpc1_1 gpc3276 (
      {stage0_11[511]},
      {stage1_11[317]}
   );
   gpc1_1 gpc3277 (
      {stage0_14[429]},
      {stage1_14[173]}
   );
   gpc1_1 gpc3278 (
      {stage0_14[430]},
      {stage1_14[174]}
   );
   gpc1_1 gpc3279 (
      {stage0_14[431]},
      {stage1_14[175]}
   );
   gpc1_1 gpc3280 (
      {stage0_14[432]},
      {stage1_14[176]}
   );
   gpc1_1 gpc3281 (
      {stage0_14[433]},
      {stage1_14[177]}
   );
   gpc1_1 gpc3282 (
      {stage0_14[434]},
      {stage1_14[178]}
   );
   gpc1_1 gpc3283 (
      {stage0_14[435]},
      {stage1_14[179]}
   );
   gpc1_1 gpc3284 (
      {stage0_14[436]},
      {stage1_14[180]}
   );
   gpc1_1 gpc3285 (
      {stage0_14[437]},
      {stage1_14[181]}
   );
   gpc1_1 gpc3286 (
      {stage0_14[438]},
      {stage1_14[182]}
   );
   gpc1_1 gpc3287 (
      {stage0_14[439]},
      {stage1_14[183]}
   );
   gpc1_1 gpc3288 (
      {stage0_14[440]},
      {stage1_14[184]}
   );
   gpc1_1 gpc3289 (
      {stage0_14[441]},
      {stage1_14[185]}
   );
   gpc1_1 gpc3290 (
      {stage0_14[442]},
      {stage1_14[186]}
   );
   gpc1_1 gpc3291 (
      {stage0_14[443]},
      {stage1_14[187]}
   );
   gpc1_1 gpc3292 (
      {stage0_14[444]},
      {stage1_14[188]}
   );
   gpc1_1 gpc3293 (
      {stage0_14[445]},
      {stage1_14[189]}
   );
   gpc1_1 gpc3294 (
      {stage0_14[446]},
      {stage1_14[190]}
   );
   gpc1_1 gpc3295 (
      {stage0_14[447]},
      {stage1_14[191]}
   );
   gpc1_1 gpc3296 (
      {stage0_14[448]},
      {stage1_14[192]}
   );
   gpc1_1 gpc3297 (
      {stage0_14[449]},
      {stage1_14[193]}
   );
   gpc1_1 gpc3298 (
      {stage0_14[450]},
      {stage1_14[194]}
   );
   gpc1_1 gpc3299 (
      {stage0_14[451]},
      {stage1_14[195]}
   );
   gpc1_1 gpc3300 (
      {stage0_14[452]},
      {stage1_14[196]}
   );
   gpc1_1 gpc3301 (
      {stage0_14[453]},
      {stage1_14[197]}
   );
   gpc1_1 gpc3302 (
      {stage0_14[454]},
      {stage1_14[198]}
   );
   gpc1_1 gpc3303 (
      {stage0_14[455]},
      {stage1_14[199]}
   );
   gpc1_1 gpc3304 (
      {stage0_14[456]},
      {stage1_14[200]}
   );
   gpc1_1 gpc3305 (
      {stage0_14[457]},
      {stage1_14[201]}
   );
   gpc1_1 gpc3306 (
      {stage0_14[458]},
      {stage1_14[202]}
   );
   gpc1_1 gpc3307 (
      {stage0_14[459]},
      {stage1_14[203]}
   );
   gpc1_1 gpc3308 (
      {stage0_14[460]},
      {stage1_14[204]}
   );
   gpc1_1 gpc3309 (
      {stage0_14[461]},
      {stage1_14[205]}
   );
   gpc1_1 gpc3310 (
      {stage0_14[462]},
      {stage1_14[206]}
   );
   gpc1_1 gpc3311 (
      {stage0_14[463]},
      {stage1_14[207]}
   );
   gpc1_1 gpc3312 (
      {stage0_14[464]},
      {stage1_14[208]}
   );
   gpc1_1 gpc3313 (
      {stage0_14[465]},
      {stage1_14[209]}
   );
   gpc1_1 gpc3314 (
      {stage0_14[466]},
      {stage1_14[210]}
   );
   gpc1_1 gpc3315 (
      {stage0_14[467]},
      {stage1_14[211]}
   );
   gpc1_1 gpc3316 (
      {stage0_14[468]},
      {stage1_14[212]}
   );
   gpc1_1 gpc3317 (
      {stage0_14[469]},
      {stage1_14[213]}
   );
   gpc1_1 gpc3318 (
      {stage0_14[470]},
      {stage1_14[214]}
   );
   gpc1_1 gpc3319 (
      {stage0_14[471]},
      {stage1_14[215]}
   );
   gpc1_1 gpc3320 (
      {stage0_14[472]},
      {stage1_14[216]}
   );
   gpc1_1 gpc3321 (
      {stage0_14[473]},
      {stage1_14[217]}
   );
   gpc1_1 gpc3322 (
      {stage0_14[474]},
      {stage1_14[218]}
   );
   gpc1_1 gpc3323 (
      {stage0_14[475]},
      {stage1_14[219]}
   );
   gpc1_1 gpc3324 (
      {stage0_14[476]},
      {stage1_14[220]}
   );
   gpc1_1 gpc3325 (
      {stage0_14[477]},
      {stage1_14[221]}
   );
   gpc1_1 gpc3326 (
      {stage0_14[478]},
      {stage1_14[222]}
   );
   gpc1_1 gpc3327 (
      {stage0_14[479]},
      {stage1_14[223]}
   );
   gpc1_1 gpc3328 (
      {stage0_14[480]},
      {stage1_14[224]}
   );
   gpc1_1 gpc3329 (
      {stage0_14[481]},
      {stage1_14[225]}
   );
   gpc1_1 gpc3330 (
      {stage0_14[482]},
      {stage1_14[226]}
   );
   gpc1_1 gpc3331 (
      {stage0_14[483]},
      {stage1_14[227]}
   );
   gpc1_1 gpc3332 (
      {stage0_14[484]},
      {stage1_14[228]}
   );
   gpc1_1 gpc3333 (
      {stage0_14[485]},
      {stage1_14[229]}
   );
   gpc1_1 gpc3334 (
      {stage0_14[486]},
      {stage1_14[230]}
   );
   gpc1_1 gpc3335 (
      {stage0_14[487]},
      {stage1_14[231]}
   );
   gpc1_1 gpc3336 (
      {stage0_14[488]},
      {stage1_14[232]}
   );
   gpc1_1 gpc3337 (
      {stage0_14[489]},
      {stage1_14[233]}
   );
   gpc1_1 gpc3338 (
      {stage0_14[490]},
      {stage1_14[234]}
   );
   gpc1_1 gpc3339 (
      {stage0_14[491]},
      {stage1_14[235]}
   );
   gpc1_1 gpc3340 (
      {stage0_14[492]},
      {stage1_14[236]}
   );
   gpc1_1 gpc3341 (
      {stage0_14[493]},
      {stage1_14[237]}
   );
   gpc1_1 gpc3342 (
      {stage0_14[494]},
      {stage1_14[238]}
   );
   gpc1_1 gpc3343 (
      {stage0_14[495]},
      {stage1_14[239]}
   );
   gpc1_1 gpc3344 (
      {stage0_14[496]},
      {stage1_14[240]}
   );
   gpc1_1 gpc3345 (
      {stage0_14[497]},
      {stage1_14[241]}
   );
   gpc1_1 gpc3346 (
      {stage0_14[498]},
      {stage1_14[242]}
   );
   gpc1_1 gpc3347 (
      {stage0_14[499]},
      {stage1_14[243]}
   );
   gpc1_1 gpc3348 (
      {stage0_14[500]},
      {stage1_14[244]}
   );
   gpc1_1 gpc3349 (
      {stage0_14[501]},
      {stage1_14[245]}
   );
   gpc1_1 gpc3350 (
      {stage0_14[502]},
      {stage1_14[246]}
   );
   gpc1_1 gpc3351 (
      {stage0_14[503]},
      {stage1_14[247]}
   );
   gpc1_1 gpc3352 (
      {stage0_14[504]},
      {stage1_14[248]}
   );
   gpc1_1 gpc3353 (
      {stage0_14[505]},
      {stage1_14[249]}
   );
   gpc1_1 gpc3354 (
      {stage0_14[506]},
      {stage1_14[250]}
   );
   gpc1_1 gpc3355 (
      {stage0_14[507]},
      {stage1_14[251]}
   );
   gpc1_1 gpc3356 (
      {stage0_14[508]},
      {stage1_14[252]}
   );
   gpc1_1 gpc3357 (
      {stage0_14[509]},
      {stage1_14[253]}
   );
   gpc1_1 gpc3358 (
      {stage0_14[510]},
      {stage1_14[254]}
   );
   gpc1_1 gpc3359 (
      {stage0_14[511]},
      {stage1_14[255]}
   );
   gpc1_1 gpc3360 (
      {stage0_15[457]},
      {stage1_15[203]}
   );
   gpc1_1 gpc3361 (
      {stage0_15[458]},
      {stage1_15[204]}
   );
   gpc1_1 gpc3362 (
      {stage0_15[459]},
      {stage1_15[205]}
   );
   gpc1_1 gpc3363 (
      {stage0_15[460]},
      {stage1_15[206]}
   );
   gpc1_1 gpc3364 (
      {stage0_15[461]},
      {stage1_15[207]}
   );
   gpc1_1 gpc3365 (
      {stage0_15[462]},
      {stage1_15[208]}
   );
   gpc1_1 gpc3366 (
      {stage0_15[463]},
      {stage1_15[209]}
   );
   gpc1_1 gpc3367 (
      {stage0_15[464]},
      {stage1_15[210]}
   );
   gpc1_1 gpc3368 (
      {stage0_15[465]},
      {stage1_15[211]}
   );
   gpc1_1 gpc3369 (
      {stage0_15[466]},
      {stage1_15[212]}
   );
   gpc1_1 gpc3370 (
      {stage0_15[467]},
      {stage1_15[213]}
   );
   gpc1_1 gpc3371 (
      {stage0_15[468]},
      {stage1_15[214]}
   );
   gpc1_1 gpc3372 (
      {stage0_15[469]},
      {stage1_15[215]}
   );
   gpc1_1 gpc3373 (
      {stage0_15[470]},
      {stage1_15[216]}
   );
   gpc1_1 gpc3374 (
      {stage0_15[471]},
      {stage1_15[217]}
   );
   gpc1_1 gpc3375 (
      {stage0_15[472]},
      {stage1_15[218]}
   );
   gpc1_1 gpc3376 (
      {stage0_15[473]},
      {stage1_15[219]}
   );
   gpc1_1 gpc3377 (
      {stage0_15[474]},
      {stage1_15[220]}
   );
   gpc1_1 gpc3378 (
      {stage0_15[475]},
      {stage1_15[221]}
   );
   gpc1_1 gpc3379 (
      {stage0_15[476]},
      {stage1_15[222]}
   );
   gpc1_1 gpc3380 (
      {stage0_15[477]},
      {stage1_15[223]}
   );
   gpc1_1 gpc3381 (
      {stage0_15[478]},
      {stage1_15[224]}
   );
   gpc1_1 gpc3382 (
      {stage0_15[479]},
      {stage1_15[225]}
   );
   gpc1_1 gpc3383 (
      {stage0_15[480]},
      {stage1_15[226]}
   );
   gpc1_1 gpc3384 (
      {stage0_15[481]},
      {stage1_15[227]}
   );
   gpc1_1 gpc3385 (
      {stage0_15[482]},
      {stage1_15[228]}
   );
   gpc1_1 gpc3386 (
      {stage0_15[483]},
      {stage1_15[229]}
   );
   gpc1_1 gpc3387 (
      {stage0_15[484]},
      {stage1_15[230]}
   );
   gpc1_1 gpc3388 (
      {stage0_15[485]},
      {stage1_15[231]}
   );
   gpc1_1 gpc3389 (
      {stage0_15[486]},
      {stage1_15[232]}
   );
   gpc1_1 gpc3390 (
      {stage0_15[487]},
      {stage1_15[233]}
   );
   gpc1_1 gpc3391 (
      {stage0_15[488]},
      {stage1_15[234]}
   );
   gpc1_1 gpc3392 (
      {stage0_15[489]},
      {stage1_15[235]}
   );
   gpc1_1 gpc3393 (
      {stage0_15[490]},
      {stage1_15[236]}
   );
   gpc1_1 gpc3394 (
      {stage0_15[491]},
      {stage1_15[237]}
   );
   gpc1_1 gpc3395 (
      {stage0_15[492]},
      {stage1_15[238]}
   );
   gpc1_1 gpc3396 (
      {stage0_15[493]},
      {stage1_15[239]}
   );
   gpc1_1 gpc3397 (
      {stage0_15[494]},
      {stage1_15[240]}
   );
   gpc1_1 gpc3398 (
      {stage0_15[495]},
      {stage1_15[241]}
   );
   gpc1_1 gpc3399 (
      {stage0_15[496]},
      {stage1_15[242]}
   );
   gpc1_1 gpc3400 (
      {stage0_15[497]},
      {stage1_15[243]}
   );
   gpc1_1 gpc3401 (
      {stage0_15[498]},
      {stage1_15[244]}
   );
   gpc1_1 gpc3402 (
      {stage0_15[499]},
      {stage1_15[245]}
   );
   gpc1_1 gpc3403 (
      {stage0_15[500]},
      {stage1_15[246]}
   );
   gpc1_1 gpc3404 (
      {stage0_15[501]},
      {stage1_15[247]}
   );
   gpc1_1 gpc3405 (
      {stage0_15[502]},
      {stage1_15[248]}
   );
   gpc1_1 gpc3406 (
      {stage0_15[503]},
      {stage1_15[249]}
   );
   gpc1_1 gpc3407 (
      {stage0_15[504]},
      {stage1_15[250]}
   );
   gpc1_1 gpc3408 (
      {stage0_15[505]},
      {stage1_15[251]}
   );
   gpc1_1 gpc3409 (
      {stage0_15[506]},
      {stage1_15[252]}
   );
   gpc1_1 gpc3410 (
      {stage0_15[507]},
      {stage1_15[253]}
   );
   gpc1_1 gpc3411 (
      {stage0_15[508]},
      {stage1_15[254]}
   );
   gpc1_1 gpc3412 (
      {stage0_15[509]},
      {stage1_15[255]}
   );
   gpc1_1 gpc3413 (
      {stage0_15[510]},
      {stage1_15[256]}
   );
   gpc1_1 gpc3414 (
      {stage0_15[511]},
      {stage1_15[257]}
   );
   gpc1_1 gpc3415 (
      {stage0_17[492]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3416 (
      {stage0_17[493]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3417 (
      {stage0_17[494]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3418 (
      {stage0_17[495]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3419 (
      {stage0_17[496]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3420 (
      {stage0_17[497]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3421 (
      {stage0_17[498]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3422 (
      {stage0_17[499]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3423 (
      {stage0_17[500]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3424 (
      {stage0_17[501]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3425 (
      {stage0_17[502]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3426 (
      {stage0_17[503]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3427 (
      {stage0_17[504]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3428 (
      {stage0_17[505]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3429 (
      {stage0_17[506]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3430 (
      {stage0_17[507]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3431 (
      {stage0_17[508]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3432 (
      {stage0_17[509]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3433 (
      {stage0_17[510]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3434 (
      {stage0_17[511]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3435 (
      {stage0_18[434]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3436 (
      {stage0_18[435]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3437 (
      {stage0_18[436]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3438 (
      {stage0_18[437]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3439 (
      {stage0_18[438]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3440 (
      {stage0_18[439]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3441 (
      {stage0_18[440]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3442 (
      {stage0_18[441]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3443 (
      {stage0_18[442]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3444 (
      {stage0_18[443]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3445 (
      {stage0_18[444]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3446 (
      {stage0_18[445]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3447 (
      {stage0_18[446]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3448 (
      {stage0_18[447]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3449 (
      {stage0_18[448]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3450 (
      {stage0_18[449]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3451 (
      {stage0_18[450]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3452 (
      {stage0_18[451]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3453 (
      {stage0_18[452]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3454 (
      {stage0_18[453]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3455 (
      {stage0_18[454]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3456 (
      {stage0_18[455]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3457 (
      {stage0_18[456]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3458 (
      {stage0_18[457]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3459 (
      {stage0_18[458]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3460 (
      {stage0_18[459]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3461 (
      {stage0_18[460]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3462 (
      {stage0_18[461]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3463 (
      {stage0_18[462]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3464 (
      {stage0_18[463]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3465 (
      {stage0_18[464]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3466 (
      {stage0_18[465]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3467 (
      {stage0_18[466]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3468 (
      {stage0_18[467]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3469 (
      {stage0_18[468]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3470 (
      {stage0_18[469]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3471 (
      {stage0_18[470]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3472 (
      {stage0_18[471]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3473 (
      {stage0_18[472]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3474 (
      {stage0_18[473]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3475 (
      {stage0_18[474]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3476 (
      {stage0_18[475]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3477 (
      {stage0_18[476]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3478 (
      {stage0_18[477]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3479 (
      {stage0_18[478]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3480 (
      {stage0_18[479]},
      {stage1_18[209]}
   );
   gpc1_1 gpc3481 (
      {stage0_18[480]},
      {stage1_18[210]}
   );
   gpc1_1 gpc3482 (
      {stage0_18[481]},
      {stage1_18[211]}
   );
   gpc1_1 gpc3483 (
      {stage0_18[482]},
      {stage1_18[212]}
   );
   gpc1_1 gpc3484 (
      {stage0_18[483]},
      {stage1_18[213]}
   );
   gpc1_1 gpc3485 (
      {stage0_18[484]},
      {stage1_18[214]}
   );
   gpc1_1 gpc3486 (
      {stage0_18[485]},
      {stage1_18[215]}
   );
   gpc1_1 gpc3487 (
      {stage0_18[486]},
      {stage1_18[216]}
   );
   gpc1_1 gpc3488 (
      {stage0_18[487]},
      {stage1_18[217]}
   );
   gpc1_1 gpc3489 (
      {stage0_18[488]},
      {stage1_18[218]}
   );
   gpc1_1 gpc3490 (
      {stage0_18[489]},
      {stage1_18[219]}
   );
   gpc1_1 gpc3491 (
      {stage0_18[490]},
      {stage1_18[220]}
   );
   gpc1_1 gpc3492 (
      {stage0_18[491]},
      {stage1_18[221]}
   );
   gpc1_1 gpc3493 (
      {stage0_18[492]},
      {stage1_18[222]}
   );
   gpc1_1 gpc3494 (
      {stage0_18[493]},
      {stage1_18[223]}
   );
   gpc1_1 gpc3495 (
      {stage0_18[494]},
      {stage1_18[224]}
   );
   gpc1_1 gpc3496 (
      {stage0_18[495]},
      {stage1_18[225]}
   );
   gpc1_1 gpc3497 (
      {stage0_18[496]},
      {stage1_18[226]}
   );
   gpc1_1 gpc3498 (
      {stage0_18[497]},
      {stage1_18[227]}
   );
   gpc1_1 gpc3499 (
      {stage0_18[498]},
      {stage1_18[228]}
   );
   gpc1_1 gpc3500 (
      {stage0_18[499]},
      {stage1_18[229]}
   );
   gpc1_1 gpc3501 (
      {stage0_18[500]},
      {stage1_18[230]}
   );
   gpc1_1 gpc3502 (
      {stage0_18[501]},
      {stage1_18[231]}
   );
   gpc1_1 gpc3503 (
      {stage0_18[502]},
      {stage1_18[232]}
   );
   gpc1_1 gpc3504 (
      {stage0_18[503]},
      {stage1_18[233]}
   );
   gpc1_1 gpc3505 (
      {stage0_18[504]},
      {stage1_18[234]}
   );
   gpc1_1 gpc3506 (
      {stage0_18[505]},
      {stage1_18[235]}
   );
   gpc1_1 gpc3507 (
      {stage0_18[506]},
      {stage1_18[236]}
   );
   gpc1_1 gpc3508 (
      {stage0_18[507]},
      {stage1_18[237]}
   );
   gpc1_1 gpc3509 (
      {stage0_18[508]},
      {stage1_18[238]}
   );
   gpc1_1 gpc3510 (
      {stage0_18[509]},
      {stage1_18[239]}
   );
   gpc1_1 gpc3511 (
      {stage0_18[510]},
      {stage1_18[240]}
   );
   gpc1_1 gpc3512 (
      {stage0_18[511]},
      {stage1_18[241]}
   );
   gpc1_1 gpc3513 (
      {stage0_19[502]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3514 (
      {stage0_19[503]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3515 (
      {stage0_19[504]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3516 (
      {stage0_19[505]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3517 (
      {stage0_19[506]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3518 (
      {stage0_19[507]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3519 (
      {stage0_19[508]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3520 (
      {stage0_19[509]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3521 (
      {stage0_19[510]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3522 (
      {stage0_19[511]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3523 (
      {stage0_20[504]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3524 (
      {stage0_20[505]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3525 (
      {stage0_20[506]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3526 (
      {stage0_20[507]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3527 (
      {stage0_20[508]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3528 (
      {stage0_20[509]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3529 (
      {stage0_20[510]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3530 (
      {stage0_20[511]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3531 (
      {stage0_21[504]},
      {stage1_21[197]}
   );
   gpc1_1 gpc3532 (
      {stage0_21[505]},
      {stage1_21[198]}
   );
   gpc1_1 gpc3533 (
      {stage0_21[506]},
      {stage1_21[199]}
   );
   gpc1_1 gpc3534 (
      {stage0_21[507]},
      {stage1_21[200]}
   );
   gpc1_1 gpc3535 (
      {stage0_21[508]},
      {stage1_21[201]}
   );
   gpc1_1 gpc3536 (
      {stage0_21[509]},
      {stage1_21[202]}
   );
   gpc1_1 gpc3537 (
      {stage0_21[510]},
      {stage1_21[203]}
   );
   gpc1_1 gpc3538 (
      {stage0_21[511]},
      {stage1_21[204]}
   );
   gpc1_1 gpc3539 (
      {stage0_22[481]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3540 (
      {stage0_22[482]},
      {stage1_22[171]}
   );
   gpc1_1 gpc3541 (
      {stage0_22[483]},
      {stage1_22[172]}
   );
   gpc1_1 gpc3542 (
      {stage0_22[484]},
      {stage1_22[173]}
   );
   gpc1_1 gpc3543 (
      {stage0_22[485]},
      {stage1_22[174]}
   );
   gpc1_1 gpc3544 (
      {stage0_22[486]},
      {stage1_22[175]}
   );
   gpc1_1 gpc3545 (
      {stage0_22[487]},
      {stage1_22[176]}
   );
   gpc1_1 gpc3546 (
      {stage0_22[488]},
      {stage1_22[177]}
   );
   gpc1_1 gpc3547 (
      {stage0_22[489]},
      {stage1_22[178]}
   );
   gpc1_1 gpc3548 (
      {stage0_22[490]},
      {stage1_22[179]}
   );
   gpc1_1 gpc3549 (
      {stage0_22[491]},
      {stage1_22[180]}
   );
   gpc1_1 gpc3550 (
      {stage0_22[492]},
      {stage1_22[181]}
   );
   gpc1_1 gpc3551 (
      {stage0_22[493]},
      {stage1_22[182]}
   );
   gpc1_1 gpc3552 (
      {stage0_22[494]},
      {stage1_22[183]}
   );
   gpc1_1 gpc3553 (
      {stage0_22[495]},
      {stage1_22[184]}
   );
   gpc1_1 gpc3554 (
      {stage0_22[496]},
      {stage1_22[185]}
   );
   gpc1_1 gpc3555 (
      {stage0_22[497]},
      {stage1_22[186]}
   );
   gpc1_1 gpc3556 (
      {stage0_22[498]},
      {stage1_22[187]}
   );
   gpc1_1 gpc3557 (
      {stage0_22[499]},
      {stage1_22[188]}
   );
   gpc1_1 gpc3558 (
      {stage0_22[500]},
      {stage1_22[189]}
   );
   gpc1_1 gpc3559 (
      {stage0_22[501]},
      {stage1_22[190]}
   );
   gpc1_1 gpc3560 (
      {stage0_22[502]},
      {stage1_22[191]}
   );
   gpc1_1 gpc3561 (
      {stage0_22[503]},
      {stage1_22[192]}
   );
   gpc1_1 gpc3562 (
      {stage0_22[504]},
      {stage1_22[193]}
   );
   gpc1_1 gpc3563 (
      {stage0_22[505]},
      {stage1_22[194]}
   );
   gpc1_1 gpc3564 (
      {stage0_22[506]},
      {stage1_22[195]}
   );
   gpc1_1 gpc3565 (
      {stage0_22[507]},
      {stage1_22[196]}
   );
   gpc1_1 gpc3566 (
      {stage0_22[508]},
      {stage1_22[197]}
   );
   gpc1_1 gpc3567 (
      {stage0_22[509]},
      {stage1_22[198]}
   );
   gpc1_1 gpc3568 (
      {stage0_22[510]},
      {stage1_22[199]}
   );
   gpc1_1 gpc3569 (
      {stage0_22[511]},
      {stage1_22[200]}
   );
   gpc1_1 gpc3570 (
      {stage0_23[418]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3571 (
      {stage0_23[419]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3572 (
      {stage0_23[420]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3573 (
      {stage0_23[421]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3574 (
      {stage0_23[422]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3575 (
      {stage0_23[423]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3576 (
      {stage0_23[424]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3577 (
      {stage0_23[425]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3578 (
      {stage0_23[426]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3579 (
      {stage0_23[427]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3580 (
      {stage0_23[428]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3581 (
      {stage0_23[429]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3582 (
      {stage0_23[430]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3583 (
      {stage0_23[431]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3584 (
      {stage0_23[432]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3585 (
      {stage0_23[433]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3586 (
      {stage0_23[434]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3587 (
      {stage0_23[435]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3588 (
      {stage0_23[436]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3589 (
      {stage0_23[437]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3590 (
      {stage0_23[438]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3591 (
      {stage0_23[439]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3592 (
      {stage0_23[440]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3593 (
      {stage0_23[441]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3594 (
      {stage0_23[442]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3595 (
      {stage0_23[443]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3596 (
      {stage0_23[444]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3597 (
      {stage0_23[445]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3598 (
      {stage0_23[446]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3599 (
      {stage0_23[447]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3600 (
      {stage0_23[448]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3601 (
      {stage0_23[449]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3602 (
      {stage0_23[450]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3603 (
      {stage0_23[451]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3604 (
      {stage0_23[452]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3605 (
      {stage0_23[453]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3606 (
      {stage0_23[454]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3607 (
      {stage0_23[455]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3608 (
      {stage0_23[456]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3609 (
      {stage0_23[457]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3610 (
      {stage0_23[458]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3611 (
      {stage0_23[459]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3612 (
      {stage0_23[460]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3613 (
      {stage0_23[461]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3614 (
      {stage0_23[462]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3615 (
      {stage0_23[463]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3616 (
      {stage0_23[464]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3617 (
      {stage0_23[465]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3618 (
      {stage0_23[466]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3619 (
      {stage0_23[467]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3620 (
      {stage0_23[468]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3621 (
      {stage0_23[469]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3622 (
      {stage0_23[470]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3623 (
      {stage0_23[471]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3624 (
      {stage0_23[472]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3625 (
      {stage0_23[473]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3626 (
      {stage0_23[474]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3627 (
      {stage0_23[475]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3628 (
      {stage0_23[476]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3629 (
      {stage0_23[477]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3630 (
      {stage0_23[478]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3631 (
      {stage0_23[479]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3632 (
      {stage0_23[480]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3633 (
      {stage0_23[481]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3634 (
      {stage0_23[482]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3635 (
      {stage0_23[483]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3636 (
      {stage0_23[484]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3637 (
      {stage0_23[485]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3638 (
      {stage0_23[486]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3639 (
      {stage0_23[487]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3640 (
      {stage0_23[488]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3641 (
      {stage0_23[489]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3642 (
      {stage0_23[490]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3643 (
      {stage0_23[491]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3644 (
      {stage0_23[492]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3645 (
      {stage0_23[493]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3646 (
      {stage0_23[494]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3647 (
      {stage0_23[495]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3648 (
      {stage0_23[496]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3649 (
      {stage0_23[497]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3650 (
      {stage0_23[498]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3651 (
      {stage0_23[499]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3652 (
      {stage0_23[500]},
      {stage1_23[287]}
   );
   gpc1_1 gpc3653 (
      {stage0_23[501]},
      {stage1_23[288]}
   );
   gpc1_1 gpc3654 (
      {stage0_23[502]},
      {stage1_23[289]}
   );
   gpc1_1 gpc3655 (
      {stage0_23[503]},
      {stage1_23[290]}
   );
   gpc1_1 gpc3656 (
      {stage0_23[504]},
      {stage1_23[291]}
   );
   gpc1_1 gpc3657 (
      {stage0_23[505]},
      {stage1_23[292]}
   );
   gpc1_1 gpc3658 (
      {stage0_23[506]},
      {stage1_23[293]}
   );
   gpc1_1 gpc3659 (
      {stage0_23[507]},
      {stage1_23[294]}
   );
   gpc1_1 gpc3660 (
      {stage0_23[508]},
      {stage1_23[295]}
   );
   gpc1_1 gpc3661 (
      {stage0_23[509]},
      {stage1_23[296]}
   );
   gpc1_1 gpc3662 (
      {stage0_23[510]},
      {stage1_23[297]}
   );
   gpc1_1 gpc3663 (
      {stage0_23[511]},
      {stage1_23[298]}
   );
   gpc1_1 gpc3664 (
      {stage0_24[499]},
      {stage1_24[222]}
   );
   gpc1_1 gpc3665 (
      {stage0_24[500]},
      {stage1_24[223]}
   );
   gpc1_1 gpc3666 (
      {stage0_24[501]},
      {stage1_24[224]}
   );
   gpc1_1 gpc3667 (
      {stage0_24[502]},
      {stage1_24[225]}
   );
   gpc1_1 gpc3668 (
      {stage0_24[503]},
      {stage1_24[226]}
   );
   gpc1_1 gpc3669 (
      {stage0_24[504]},
      {stage1_24[227]}
   );
   gpc1_1 gpc3670 (
      {stage0_24[505]},
      {stage1_24[228]}
   );
   gpc1_1 gpc3671 (
      {stage0_24[506]},
      {stage1_24[229]}
   );
   gpc1_1 gpc3672 (
      {stage0_24[507]},
      {stage1_24[230]}
   );
   gpc1_1 gpc3673 (
      {stage0_24[508]},
      {stage1_24[231]}
   );
   gpc1_1 gpc3674 (
      {stage0_24[509]},
      {stage1_24[232]}
   );
   gpc1_1 gpc3675 (
      {stage0_24[510]},
      {stage1_24[233]}
   );
   gpc1_1 gpc3676 (
      {stage0_24[511]},
      {stage1_24[234]}
   );
   gpc1_1 gpc3677 (
      {stage0_25[506]},
      {stage1_25[205]}
   );
   gpc1_1 gpc3678 (
      {stage0_25[507]},
      {stage1_25[206]}
   );
   gpc1_1 gpc3679 (
      {stage0_25[508]},
      {stage1_25[207]}
   );
   gpc1_1 gpc3680 (
      {stage0_25[509]},
      {stage1_25[208]}
   );
   gpc1_1 gpc3681 (
      {stage0_25[510]},
      {stage1_25[209]}
   );
   gpc1_1 gpc3682 (
      {stage0_25[511]},
      {stage1_25[210]}
   );
   gpc1_1 gpc3683 (
      {stage0_26[503]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3684 (
      {stage0_26[504]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3685 (
      {stage0_26[505]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3686 (
      {stage0_26[506]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3687 (
      {stage0_26[507]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3688 (
      {stage0_26[508]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3689 (
      {stage0_26[509]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3690 (
      {stage0_26[510]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3691 (
      {stage0_26[511]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3692 (
      {stage0_27[503]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3693 (
      {stage0_27[504]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3694 (
      {stage0_27[505]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3695 (
      {stage0_27[506]},
      {stage1_27[206]}
   );
   gpc1_1 gpc3696 (
      {stage0_27[507]},
      {stage1_27[207]}
   );
   gpc1_1 gpc3697 (
      {stage0_27[508]},
      {stage1_27[208]}
   );
   gpc1_1 gpc3698 (
      {stage0_27[509]},
      {stage1_27[209]}
   );
   gpc1_1 gpc3699 (
      {stage0_27[510]},
      {stage1_27[210]}
   );
   gpc1_1 gpc3700 (
      {stage0_27[511]},
      {stage1_27[211]}
   );
   gpc1_1 gpc3701 (
      {stage0_28[500]},
      {stage1_28[237]}
   );
   gpc1_1 gpc3702 (
      {stage0_28[501]},
      {stage1_28[238]}
   );
   gpc1_1 gpc3703 (
      {stage0_28[502]},
      {stage1_28[239]}
   );
   gpc1_1 gpc3704 (
      {stage0_28[503]},
      {stage1_28[240]}
   );
   gpc1_1 gpc3705 (
      {stage0_28[504]},
      {stage1_28[241]}
   );
   gpc1_1 gpc3706 (
      {stage0_28[505]},
      {stage1_28[242]}
   );
   gpc1_1 gpc3707 (
      {stage0_28[506]},
      {stage1_28[243]}
   );
   gpc1_1 gpc3708 (
      {stage0_28[507]},
      {stage1_28[244]}
   );
   gpc1_1 gpc3709 (
      {stage0_28[508]},
      {stage1_28[245]}
   );
   gpc1_1 gpc3710 (
      {stage0_28[509]},
      {stage1_28[246]}
   );
   gpc1_1 gpc3711 (
      {stage0_28[510]},
      {stage1_28[247]}
   );
   gpc1_1 gpc3712 (
      {stage0_28[511]},
      {stage1_28[248]}
   );
   gpc1_1 gpc3713 (
      {stage0_29[510]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3714 (
      {stage0_29[511]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3715 (
      {stage0_30[443]},
      {stage1_30[164]}
   );
   gpc1_1 gpc3716 (
      {stage0_30[444]},
      {stage1_30[165]}
   );
   gpc1_1 gpc3717 (
      {stage0_30[445]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3718 (
      {stage0_30[446]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3719 (
      {stage0_30[447]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3720 (
      {stage0_30[448]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3721 (
      {stage0_30[449]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3722 (
      {stage0_30[450]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3723 (
      {stage0_30[451]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3724 (
      {stage0_30[452]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3725 (
      {stage0_30[453]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3726 (
      {stage0_30[454]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3727 (
      {stage0_30[455]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3728 (
      {stage0_30[456]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3729 (
      {stage0_30[457]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3730 (
      {stage0_30[458]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3731 (
      {stage0_30[459]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3732 (
      {stage0_30[460]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3733 (
      {stage0_30[461]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3734 (
      {stage0_30[462]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3735 (
      {stage0_30[463]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3736 (
      {stage0_30[464]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3737 (
      {stage0_30[465]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3738 (
      {stage0_30[466]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3739 (
      {stage0_30[467]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3740 (
      {stage0_30[468]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3741 (
      {stage0_30[469]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3742 (
      {stage0_30[470]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3743 (
      {stage0_30[471]},
      {stage1_30[192]}
   );
   gpc1_1 gpc3744 (
      {stage0_30[472]},
      {stage1_30[193]}
   );
   gpc1_1 gpc3745 (
      {stage0_30[473]},
      {stage1_30[194]}
   );
   gpc1_1 gpc3746 (
      {stage0_30[474]},
      {stage1_30[195]}
   );
   gpc1_1 gpc3747 (
      {stage0_30[475]},
      {stage1_30[196]}
   );
   gpc1_1 gpc3748 (
      {stage0_30[476]},
      {stage1_30[197]}
   );
   gpc1_1 gpc3749 (
      {stage0_30[477]},
      {stage1_30[198]}
   );
   gpc1_1 gpc3750 (
      {stage0_30[478]},
      {stage1_30[199]}
   );
   gpc1_1 gpc3751 (
      {stage0_30[479]},
      {stage1_30[200]}
   );
   gpc1_1 gpc3752 (
      {stage0_30[480]},
      {stage1_30[201]}
   );
   gpc1_1 gpc3753 (
      {stage0_30[481]},
      {stage1_30[202]}
   );
   gpc1_1 gpc3754 (
      {stage0_30[482]},
      {stage1_30[203]}
   );
   gpc1_1 gpc3755 (
      {stage0_30[483]},
      {stage1_30[204]}
   );
   gpc1_1 gpc3756 (
      {stage0_30[484]},
      {stage1_30[205]}
   );
   gpc1_1 gpc3757 (
      {stage0_30[485]},
      {stage1_30[206]}
   );
   gpc1_1 gpc3758 (
      {stage0_30[486]},
      {stage1_30[207]}
   );
   gpc1_1 gpc3759 (
      {stage0_30[487]},
      {stage1_30[208]}
   );
   gpc1_1 gpc3760 (
      {stage0_30[488]},
      {stage1_30[209]}
   );
   gpc1_1 gpc3761 (
      {stage0_30[489]},
      {stage1_30[210]}
   );
   gpc1_1 gpc3762 (
      {stage0_30[490]},
      {stage1_30[211]}
   );
   gpc1_1 gpc3763 (
      {stage0_30[491]},
      {stage1_30[212]}
   );
   gpc1_1 gpc3764 (
      {stage0_30[492]},
      {stage1_30[213]}
   );
   gpc1_1 gpc3765 (
      {stage0_30[493]},
      {stage1_30[214]}
   );
   gpc1_1 gpc3766 (
      {stage0_30[494]},
      {stage1_30[215]}
   );
   gpc1_1 gpc3767 (
      {stage0_30[495]},
      {stage1_30[216]}
   );
   gpc1_1 gpc3768 (
      {stage0_30[496]},
      {stage1_30[217]}
   );
   gpc1_1 gpc3769 (
      {stage0_30[497]},
      {stage1_30[218]}
   );
   gpc1_1 gpc3770 (
      {stage0_30[498]},
      {stage1_30[219]}
   );
   gpc1_1 gpc3771 (
      {stage0_30[499]},
      {stage1_30[220]}
   );
   gpc1_1 gpc3772 (
      {stage0_30[500]},
      {stage1_30[221]}
   );
   gpc1_1 gpc3773 (
      {stage0_30[501]},
      {stage1_30[222]}
   );
   gpc1_1 gpc3774 (
      {stage0_30[502]},
      {stage1_30[223]}
   );
   gpc1_1 gpc3775 (
      {stage0_30[503]},
      {stage1_30[224]}
   );
   gpc1_1 gpc3776 (
      {stage0_30[504]},
      {stage1_30[225]}
   );
   gpc1_1 gpc3777 (
      {stage0_30[505]},
      {stage1_30[226]}
   );
   gpc1_1 gpc3778 (
      {stage0_30[506]},
      {stage1_30[227]}
   );
   gpc1_1 gpc3779 (
      {stage0_30[507]},
      {stage1_30[228]}
   );
   gpc1_1 gpc3780 (
      {stage0_30[508]},
      {stage1_30[229]}
   );
   gpc1_1 gpc3781 (
      {stage0_30[509]},
      {stage1_30[230]}
   );
   gpc1_1 gpc3782 (
      {stage0_30[510]},
      {stage1_30[231]}
   );
   gpc1_1 gpc3783 (
      {stage0_30[511]},
      {stage1_30[232]}
   );
   gpc1_1 gpc3784 (
      {stage0_31[494]},
      {stage1_31[194]}
   );
   gpc1_1 gpc3785 (
      {stage0_31[495]},
      {stage1_31[195]}
   );
   gpc1_1 gpc3786 (
      {stage0_31[496]},
      {stage1_31[196]}
   );
   gpc1_1 gpc3787 (
      {stage0_31[497]},
      {stage1_31[197]}
   );
   gpc1_1 gpc3788 (
      {stage0_31[498]},
      {stage1_31[198]}
   );
   gpc1_1 gpc3789 (
      {stage0_31[499]},
      {stage1_31[199]}
   );
   gpc1_1 gpc3790 (
      {stage0_31[500]},
      {stage1_31[200]}
   );
   gpc1_1 gpc3791 (
      {stage0_31[501]},
      {stage1_31[201]}
   );
   gpc1_1 gpc3792 (
      {stage0_31[502]},
      {stage1_31[202]}
   );
   gpc1_1 gpc3793 (
      {stage0_31[503]},
      {stage1_31[203]}
   );
   gpc1_1 gpc3794 (
      {stage0_31[504]},
      {stage1_31[204]}
   );
   gpc1_1 gpc3795 (
      {stage0_31[505]},
      {stage1_31[205]}
   );
   gpc1_1 gpc3796 (
      {stage0_31[506]},
      {stage1_31[206]}
   );
   gpc1_1 gpc3797 (
      {stage0_31[507]},
      {stage1_31[207]}
   );
   gpc1_1 gpc3798 (
      {stage0_31[508]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3799 (
      {stage0_31[509]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3800 (
      {stage0_31[510]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3801 (
      {stage0_31[511]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3802 (
      {stage0_32[303]},
      {stage1_32[206]}
   );
   gpc1_1 gpc3803 (
      {stage0_32[304]},
      {stage1_32[207]}
   );
   gpc1_1 gpc3804 (
      {stage0_32[305]},
      {stage1_32[208]}
   );
   gpc1_1 gpc3805 (
      {stage0_32[306]},
      {stage1_32[209]}
   );
   gpc1_1 gpc3806 (
      {stage0_32[307]},
      {stage1_32[210]}
   );
   gpc1_1 gpc3807 (
      {stage0_32[308]},
      {stage1_32[211]}
   );
   gpc1_1 gpc3808 (
      {stage0_32[309]},
      {stage1_32[212]}
   );
   gpc1_1 gpc3809 (
      {stage0_32[310]},
      {stage1_32[213]}
   );
   gpc1_1 gpc3810 (
      {stage0_32[311]},
      {stage1_32[214]}
   );
   gpc1_1 gpc3811 (
      {stage0_32[312]},
      {stage1_32[215]}
   );
   gpc1_1 gpc3812 (
      {stage0_32[313]},
      {stage1_32[216]}
   );
   gpc1_1 gpc3813 (
      {stage0_32[314]},
      {stage1_32[217]}
   );
   gpc1_1 gpc3814 (
      {stage0_32[315]},
      {stage1_32[218]}
   );
   gpc1_1 gpc3815 (
      {stage0_32[316]},
      {stage1_32[219]}
   );
   gpc1_1 gpc3816 (
      {stage0_32[317]},
      {stage1_32[220]}
   );
   gpc1_1 gpc3817 (
      {stage0_32[318]},
      {stage1_32[221]}
   );
   gpc1_1 gpc3818 (
      {stage0_32[319]},
      {stage1_32[222]}
   );
   gpc1_1 gpc3819 (
      {stage0_32[320]},
      {stage1_32[223]}
   );
   gpc1_1 gpc3820 (
      {stage0_32[321]},
      {stage1_32[224]}
   );
   gpc1_1 gpc3821 (
      {stage0_32[322]},
      {stage1_32[225]}
   );
   gpc1_1 gpc3822 (
      {stage0_32[323]},
      {stage1_32[226]}
   );
   gpc1_1 gpc3823 (
      {stage0_32[324]},
      {stage1_32[227]}
   );
   gpc1_1 gpc3824 (
      {stage0_32[325]},
      {stage1_32[228]}
   );
   gpc1_1 gpc3825 (
      {stage0_32[326]},
      {stage1_32[229]}
   );
   gpc1_1 gpc3826 (
      {stage0_32[327]},
      {stage1_32[230]}
   );
   gpc1_1 gpc3827 (
      {stage0_32[328]},
      {stage1_32[231]}
   );
   gpc1_1 gpc3828 (
      {stage0_32[329]},
      {stage1_32[232]}
   );
   gpc1_1 gpc3829 (
      {stage0_32[330]},
      {stage1_32[233]}
   );
   gpc1_1 gpc3830 (
      {stage0_32[331]},
      {stage1_32[234]}
   );
   gpc1_1 gpc3831 (
      {stage0_32[332]},
      {stage1_32[235]}
   );
   gpc1_1 gpc3832 (
      {stage0_32[333]},
      {stage1_32[236]}
   );
   gpc1_1 gpc3833 (
      {stage0_32[334]},
      {stage1_32[237]}
   );
   gpc1_1 gpc3834 (
      {stage0_32[335]},
      {stage1_32[238]}
   );
   gpc1_1 gpc3835 (
      {stage0_32[336]},
      {stage1_32[239]}
   );
   gpc1_1 gpc3836 (
      {stage0_32[337]},
      {stage1_32[240]}
   );
   gpc1_1 gpc3837 (
      {stage0_32[338]},
      {stage1_32[241]}
   );
   gpc1_1 gpc3838 (
      {stage0_32[339]},
      {stage1_32[242]}
   );
   gpc1_1 gpc3839 (
      {stage0_32[340]},
      {stage1_32[243]}
   );
   gpc1_1 gpc3840 (
      {stage0_32[341]},
      {stage1_32[244]}
   );
   gpc1_1 gpc3841 (
      {stage0_32[342]},
      {stage1_32[245]}
   );
   gpc1_1 gpc3842 (
      {stage0_32[343]},
      {stage1_32[246]}
   );
   gpc1_1 gpc3843 (
      {stage0_32[344]},
      {stage1_32[247]}
   );
   gpc1_1 gpc3844 (
      {stage0_32[345]},
      {stage1_32[248]}
   );
   gpc1_1 gpc3845 (
      {stage0_32[346]},
      {stage1_32[249]}
   );
   gpc1_1 gpc3846 (
      {stage0_32[347]},
      {stage1_32[250]}
   );
   gpc1_1 gpc3847 (
      {stage0_32[348]},
      {stage1_32[251]}
   );
   gpc1_1 gpc3848 (
      {stage0_32[349]},
      {stage1_32[252]}
   );
   gpc1_1 gpc3849 (
      {stage0_32[350]},
      {stage1_32[253]}
   );
   gpc1_1 gpc3850 (
      {stage0_32[351]},
      {stage1_32[254]}
   );
   gpc1_1 gpc3851 (
      {stage0_32[352]},
      {stage1_32[255]}
   );
   gpc1_1 gpc3852 (
      {stage0_32[353]},
      {stage1_32[256]}
   );
   gpc1_1 gpc3853 (
      {stage0_32[354]},
      {stage1_32[257]}
   );
   gpc1_1 gpc3854 (
      {stage0_32[355]},
      {stage1_32[258]}
   );
   gpc1_1 gpc3855 (
      {stage0_32[356]},
      {stage1_32[259]}
   );
   gpc1_1 gpc3856 (
      {stage0_32[357]},
      {stage1_32[260]}
   );
   gpc1_1 gpc3857 (
      {stage0_32[358]},
      {stage1_32[261]}
   );
   gpc1_1 gpc3858 (
      {stage0_32[359]},
      {stage1_32[262]}
   );
   gpc1_1 gpc3859 (
      {stage0_32[360]},
      {stage1_32[263]}
   );
   gpc1_1 gpc3860 (
      {stage0_32[361]},
      {stage1_32[264]}
   );
   gpc1_1 gpc3861 (
      {stage0_32[362]},
      {stage1_32[265]}
   );
   gpc1_1 gpc3862 (
      {stage0_32[363]},
      {stage1_32[266]}
   );
   gpc1_1 gpc3863 (
      {stage0_32[364]},
      {stage1_32[267]}
   );
   gpc1_1 gpc3864 (
      {stage0_32[365]},
      {stage1_32[268]}
   );
   gpc1_1 gpc3865 (
      {stage0_32[366]},
      {stage1_32[269]}
   );
   gpc1_1 gpc3866 (
      {stage0_32[367]},
      {stage1_32[270]}
   );
   gpc1_1 gpc3867 (
      {stage0_32[368]},
      {stage1_32[271]}
   );
   gpc1_1 gpc3868 (
      {stage0_32[369]},
      {stage1_32[272]}
   );
   gpc1_1 gpc3869 (
      {stage0_32[370]},
      {stage1_32[273]}
   );
   gpc1_1 gpc3870 (
      {stage0_32[371]},
      {stage1_32[274]}
   );
   gpc1_1 gpc3871 (
      {stage0_32[372]},
      {stage1_32[275]}
   );
   gpc1_1 gpc3872 (
      {stage0_32[373]},
      {stage1_32[276]}
   );
   gpc1_1 gpc3873 (
      {stage0_32[374]},
      {stage1_32[277]}
   );
   gpc1_1 gpc3874 (
      {stage0_32[375]},
      {stage1_32[278]}
   );
   gpc1_1 gpc3875 (
      {stage0_32[376]},
      {stage1_32[279]}
   );
   gpc1_1 gpc3876 (
      {stage0_32[377]},
      {stage1_32[280]}
   );
   gpc1_1 gpc3877 (
      {stage0_32[378]},
      {stage1_32[281]}
   );
   gpc1_1 gpc3878 (
      {stage0_32[379]},
      {stage1_32[282]}
   );
   gpc1_1 gpc3879 (
      {stage0_32[380]},
      {stage1_32[283]}
   );
   gpc1_1 gpc3880 (
      {stage0_32[381]},
      {stage1_32[284]}
   );
   gpc1_1 gpc3881 (
      {stage0_32[382]},
      {stage1_32[285]}
   );
   gpc1_1 gpc3882 (
      {stage0_32[383]},
      {stage1_32[286]}
   );
   gpc1_1 gpc3883 (
      {stage0_32[384]},
      {stage1_32[287]}
   );
   gpc1_1 gpc3884 (
      {stage0_32[385]},
      {stage1_32[288]}
   );
   gpc1_1 gpc3885 (
      {stage0_32[386]},
      {stage1_32[289]}
   );
   gpc1_1 gpc3886 (
      {stage0_32[387]},
      {stage1_32[290]}
   );
   gpc1_1 gpc3887 (
      {stage0_32[388]},
      {stage1_32[291]}
   );
   gpc1_1 gpc3888 (
      {stage0_32[389]},
      {stage1_32[292]}
   );
   gpc1_1 gpc3889 (
      {stage0_32[390]},
      {stage1_32[293]}
   );
   gpc1_1 gpc3890 (
      {stage0_32[391]},
      {stage1_32[294]}
   );
   gpc1_1 gpc3891 (
      {stage0_32[392]},
      {stage1_32[295]}
   );
   gpc1_1 gpc3892 (
      {stage0_32[393]},
      {stage1_32[296]}
   );
   gpc1_1 gpc3893 (
      {stage0_32[394]},
      {stage1_32[297]}
   );
   gpc1_1 gpc3894 (
      {stage0_32[395]},
      {stage1_32[298]}
   );
   gpc1_1 gpc3895 (
      {stage0_32[396]},
      {stage1_32[299]}
   );
   gpc1_1 gpc3896 (
      {stage0_32[397]},
      {stage1_32[300]}
   );
   gpc1_1 gpc3897 (
      {stage0_32[398]},
      {stage1_32[301]}
   );
   gpc1_1 gpc3898 (
      {stage0_32[399]},
      {stage1_32[302]}
   );
   gpc1_1 gpc3899 (
      {stage0_32[400]},
      {stage1_32[303]}
   );
   gpc1_1 gpc3900 (
      {stage0_32[401]},
      {stage1_32[304]}
   );
   gpc1_1 gpc3901 (
      {stage0_32[402]},
      {stage1_32[305]}
   );
   gpc1_1 gpc3902 (
      {stage0_32[403]},
      {stage1_32[306]}
   );
   gpc1_1 gpc3903 (
      {stage0_32[404]},
      {stage1_32[307]}
   );
   gpc1_1 gpc3904 (
      {stage0_32[405]},
      {stage1_32[308]}
   );
   gpc1_1 gpc3905 (
      {stage0_32[406]},
      {stage1_32[309]}
   );
   gpc1_1 gpc3906 (
      {stage0_32[407]},
      {stage1_32[310]}
   );
   gpc1_1 gpc3907 (
      {stage0_32[408]},
      {stage1_32[311]}
   );
   gpc1_1 gpc3908 (
      {stage0_32[409]},
      {stage1_32[312]}
   );
   gpc1_1 gpc3909 (
      {stage0_32[410]},
      {stage1_32[313]}
   );
   gpc1_1 gpc3910 (
      {stage0_32[411]},
      {stage1_32[314]}
   );
   gpc1_1 gpc3911 (
      {stage0_32[412]},
      {stage1_32[315]}
   );
   gpc1_1 gpc3912 (
      {stage0_32[413]},
      {stage1_32[316]}
   );
   gpc1_1 gpc3913 (
      {stage0_32[414]},
      {stage1_32[317]}
   );
   gpc1_1 gpc3914 (
      {stage0_32[415]},
      {stage1_32[318]}
   );
   gpc1_1 gpc3915 (
      {stage0_32[416]},
      {stage1_32[319]}
   );
   gpc1_1 gpc3916 (
      {stage0_32[417]},
      {stage1_32[320]}
   );
   gpc1_1 gpc3917 (
      {stage0_32[418]},
      {stage1_32[321]}
   );
   gpc1_1 gpc3918 (
      {stage0_32[419]},
      {stage1_32[322]}
   );
   gpc1_1 gpc3919 (
      {stage0_32[420]},
      {stage1_32[323]}
   );
   gpc1_1 gpc3920 (
      {stage0_32[421]},
      {stage1_32[324]}
   );
   gpc1_1 gpc3921 (
      {stage0_32[422]},
      {stage1_32[325]}
   );
   gpc1_1 gpc3922 (
      {stage0_32[423]},
      {stage1_32[326]}
   );
   gpc1_1 gpc3923 (
      {stage0_32[424]},
      {stage1_32[327]}
   );
   gpc1_1 gpc3924 (
      {stage0_32[425]},
      {stage1_32[328]}
   );
   gpc1_1 gpc3925 (
      {stage0_32[426]},
      {stage1_32[329]}
   );
   gpc1_1 gpc3926 (
      {stage0_32[427]},
      {stage1_32[330]}
   );
   gpc1_1 gpc3927 (
      {stage0_32[428]},
      {stage1_32[331]}
   );
   gpc1_1 gpc3928 (
      {stage0_32[429]},
      {stage1_32[332]}
   );
   gpc1_1 gpc3929 (
      {stage0_32[430]},
      {stage1_32[333]}
   );
   gpc1_1 gpc3930 (
      {stage0_32[431]},
      {stage1_32[334]}
   );
   gpc1_1 gpc3931 (
      {stage0_32[432]},
      {stage1_32[335]}
   );
   gpc1_1 gpc3932 (
      {stage0_32[433]},
      {stage1_32[336]}
   );
   gpc1_1 gpc3933 (
      {stage0_32[434]},
      {stage1_32[337]}
   );
   gpc1_1 gpc3934 (
      {stage0_32[435]},
      {stage1_32[338]}
   );
   gpc1_1 gpc3935 (
      {stage0_32[436]},
      {stage1_32[339]}
   );
   gpc1_1 gpc3936 (
      {stage0_32[437]},
      {stage1_32[340]}
   );
   gpc1_1 gpc3937 (
      {stage0_32[438]},
      {stage1_32[341]}
   );
   gpc1_1 gpc3938 (
      {stage0_32[439]},
      {stage1_32[342]}
   );
   gpc1_1 gpc3939 (
      {stage0_32[440]},
      {stage1_32[343]}
   );
   gpc1_1 gpc3940 (
      {stage0_32[441]},
      {stage1_32[344]}
   );
   gpc1_1 gpc3941 (
      {stage0_32[442]},
      {stage1_32[345]}
   );
   gpc1_1 gpc3942 (
      {stage0_32[443]},
      {stage1_32[346]}
   );
   gpc1_1 gpc3943 (
      {stage0_32[444]},
      {stage1_32[347]}
   );
   gpc1_1 gpc3944 (
      {stage0_32[445]},
      {stage1_32[348]}
   );
   gpc1_1 gpc3945 (
      {stage0_32[446]},
      {stage1_32[349]}
   );
   gpc1_1 gpc3946 (
      {stage0_32[447]},
      {stage1_32[350]}
   );
   gpc1_1 gpc3947 (
      {stage0_32[448]},
      {stage1_32[351]}
   );
   gpc1_1 gpc3948 (
      {stage0_32[449]},
      {stage1_32[352]}
   );
   gpc1_1 gpc3949 (
      {stage0_32[450]},
      {stage1_32[353]}
   );
   gpc1_1 gpc3950 (
      {stage0_32[451]},
      {stage1_32[354]}
   );
   gpc1_1 gpc3951 (
      {stage0_32[452]},
      {stage1_32[355]}
   );
   gpc1_1 gpc3952 (
      {stage0_32[453]},
      {stage1_32[356]}
   );
   gpc1_1 gpc3953 (
      {stage0_32[454]},
      {stage1_32[357]}
   );
   gpc1_1 gpc3954 (
      {stage0_32[455]},
      {stage1_32[358]}
   );
   gpc1_1 gpc3955 (
      {stage0_32[456]},
      {stage1_32[359]}
   );
   gpc1_1 gpc3956 (
      {stage0_32[457]},
      {stage1_32[360]}
   );
   gpc1_1 gpc3957 (
      {stage0_32[458]},
      {stage1_32[361]}
   );
   gpc1_1 gpc3958 (
      {stage0_32[459]},
      {stage1_32[362]}
   );
   gpc1_1 gpc3959 (
      {stage0_32[460]},
      {stage1_32[363]}
   );
   gpc1_1 gpc3960 (
      {stage0_32[461]},
      {stage1_32[364]}
   );
   gpc1_1 gpc3961 (
      {stage0_32[462]},
      {stage1_32[365]}
   );
   gpc1_1 gpc3962 (
      {stage0_32[463]},
      {stage1_32[366]}
   );
   gpc1_1 gpc3963 (
      {stage0_32[464]},
      {stage1_32[367]}
   );
   gpc1_1 gpc3964 (
      {stage0_32[465]},
      {stage1_32[368]}
   );
   gpc1_1 gpc3965 (
      {stage0_32[466]},
      {stage1_32[369]}
   );
   gpc1_1 gpc3966 (
      {stage0_32[467]},
      {stage1_32[370]}
   );
   gpc1_1 gpc3967 (
      {stage0_32[468]},
      {stage1_32[371]}
   );
   gpc1_1 gpc3968 (
      {stage0_32[469]},
      {stage1_32[372]}
   );
   gpc1_1 gpc3969 (
      {stage0_32[470]},
      {stage1_32[373]}
   );
   gpc1_1 gpc3970 (
      {stage0_32[471]},
      {stage1_32[374]}
   );
   gpc1_1 gpc3971 (
      {stage0_32[472]},
      {stage1_32[375]}
   );
   gpc1_1 gpc3972 (
      {stage0_32[473]},
      {stage1_32[376]}
   );
   gpc1_1 gpc3973 (
      {stage0_32[474]},
      {stage1_32[377]}
   );
   gpc1_1 gpc3974 (
      {stage0_32[475]},
      {stage1_32[378]}
   );
   gpc1_1 gpc3975 (
      {stage0_32[476]},
      {stage1_32[379]}
   );
   gpc1_1 gpc3976 (
      {stage0_32[477]},
      {stage1_32[380]}
   );
   gpc1_1 gpc3977 (
      {stage0_32[478]},
      {stage1_32[381]}
   );
   gpc1_1 gpc3978 (
      {stage0_32[479]},
      {stage1_32[382]}
   );
   gpc1_1 gpc3979 (
      {stage0_32[480]},
      {stage1_32[383]}
   );
   gpc1_1 gpc3980 (
      {stage0_32[481]},
      {stage1_32[384]}
   );
   gpc1_1 gpc3981 (
      {stage0_32[482]},
      {stage1_32[385]}
   );
   gpc1_1 gpc3982 (
      {stage0_32[483]},
      {stage1_32[386]}
   );
   gpc1_1 gpc3983 (
      {stage0_32[484]},
      {stage1_32[387]}
   );
   gpc1_1 gpc3984 (
      {stage0_32[485]},
      {stage1_32[388]}
   );
   gpc1_1 gpc3985 (
      {stage0_32[486]},
      {stage1_32[389]}
   );
   gpc1_1 gpc3986 (
      {stage0_32[487]},
      {stage1_32[390]}
   );
   gpc1_1 gpc3987 (
      {stage0_32[488]},
      {stage1_32[391]}
   );
   gpc1_1 gpc3988 (
      {stage0_32[489]},
      {stage1_32[392]}
   );
   gpc1_1 gpc3989 (
      {stage0_32[490]},
      {stage1_32[393]}
   );
   gpc1_1 gpc3990 (
      {stage0_32[491]},
      {stage1_32[394]}
   );
   gpc1_1 gpc3991 (
      {stage0_32[492]},
      {stage1_32[395]}
   );
   gpc1_1 gpc3992 (
      {stage0_32[493]},
      {stage1_32[396]}
   );
   gpc1_1 gpc3993 (
      {stage0_32[494]},
      {stage1_32[397]}
   );
   gpc1_1 gpc3994 (
      {stage0_32[495]},
      {stage1_32[398]}
   );
   gpc1_1 gpc3995 (
      {stage0_32[496]},
      {stage1_32[399]}
   );
   gpc1_1 gpc3996 (
      {stage0_32[497]},
      {stage1_32[400]}
   );
   gpc1_1 gpc3997 (
      {stage0_32[498]},
      {stage1_32[401]}
   );
   gpc1_1 gpc3998 (
      {stage0_32[499]},
      {stage1_32[402]}
   );
   gpc1_1 gpc3999 (
      {stage0_32[500]},
      {stage1_32[403]}
   );
   gpc1_1 gpc4000 (
      {stage0_32[501]},
      {stage1_32[404]}
   );
   gpc1_1 gpc4001 (
      {stage0_32[502]},
      {stage1_32[405]}
   );
   gpc1_1 gpc4002 (
      {stage0_32[503]},
      {stage1_32[406]}
   );
   gpc1_1 gpc4003 (
      {stage0_32[504]},
      {stage1_32[407]}
   );
   gpc1_1 gpc4004 (
      {stage0_32[505]},
      {stage1_32[408]}
   );
   gpc1_1 gpc4005 (
      {stage0_32[506]},
      {stage1_32[409]}
   );
   gpc1_1 gpc4006 (
      {stage0_32[507]},
      {stage1_32[410]}
   );
   gpc1_1 gpc4007 (
      {stage0_32[508]},
      {stage1_32[411]}
   );
   gpc1_1 gpc4008 (
      {stage0_32[509]},
      {stage1_32[412]}
   );
   gpc1_1 gpc4009 (
      {stage0_32[510]},
      {stage1_32[413]}
   );
   gpc1_1 gpc4010 (
      {stage0_32[511]},
      {stage1_32[414]}
   );
   gpc1_1 gpc4011 (
      {stage0_33[491]},
      {stage1_33[189]}
   );
   gpc1_1 gpc4012 (
      {stage0_33[492]},
      {stage1_33[190]}
   );
   gpc1_1 gpc4013 (
      {stage0_33[493]},
      {stage1_33[191]}
   );
   gpc1_1 gpc4014 (
      {stage0_33[494]},
      {stage1_33[192]}
   );
   gpc1_1 gpc4015 (
      {stage0_33[495]},
      {stage1_33[193]}
   );
   gpc1_1 gpc4016 (
      {stage0_33[496]},
      {stage1_33[194]}
   );
   gpc1_1 gpc4017 (
      {stage0_33[497]},
      {stage1_33[195]}
   );
   gpc1_1 gpc4018 (
      {stage0_33[498]},
      {stage1_33[196]}
   );
   gpc1_1 gpc4019 (
      {stage0_33[499]},
      {stage1_33[197]}
   );
   gpc1_1 gpc4020 (
      {stage0_33[500]},
      {stage1_33[198]}
   );
   gpc1_1 gpc4021 (
      {stage0_33[501]},
      {stage1_33[199]}
   );
   gpc1_1 gpc4022 (
      {stage0_33[502]},
      {stage1_33[200]}
   );
   gpc1_1 gpc4023 (
      {stage0_33[503]},
      {stage1_33[201]}
   );
   gpc1_1 gpc4024 (
      {stage0_33[504]},
      {stage1_33[202]}
   );
   gpc1_1 gpc4025 (
      {stage0_33[505]},
      {stage1_33[203]}
   );
   gpc1_1 gpc4026 (
      {stage0_33[506]},
      {stage1_33[204]}
   );
   gpc1_1 gpc4027 (
      {stage0_33[507]},
      {stage1_33[205]}
   );
   gpc1_1 gpc4028 (
      {stage0_33[508]},
      {stage1_33[206]}
   );
   gpc1_1 gpc4029 (
      {stage0_33[509]},
      {stage1_33[207]}
   );
   gpc1_1 gpc4030 (
      {stage0_33[510]},
      {stage1_33[208]}
   );
   gpc1_1 gpc4031 (
      {stage0_33[511]},
      {stage1_33[209]}
   );
   gpc1_1 gpc4032 (
      {stage0_34[396]},
      {stage1_34[152]}
   );
   gpc1_1 gpc4033 (
      {stage0_34[397]},
      {stage1_34[153]}
   );
   gpc1_1 gpc4034 (
      {stage0_34[398]},
      {stage1_34[154]}
   );
   gpc1_1 gpc4035 (
      {stage0_34[399]},
      {stage1_34[155]}
   );
   gpc1_1 gpc4036 (
      {stage0_34[400]},
      {stage1_34[156]}
   );
   gpc1_1 gpc4037 (
      {stage0_34[401]},
      {stage1_34[157]}
   );
   gpc1_1 gpc4038 (
      {stage0_34[402]},
      {stage1_34[158]}
   );
   gpc1_1 gpc4039 (
      {stage0_34[403]},
      {stage1_34[159]}
   );
   gpc1_1 gpc4040 (
      {stage0_34[404]},
      {stage1_34[160]}
   );
   gpc1_1 gpc4041 (
      {stage0_34[405]},
      {stage1_34[161]}
   );
   gpc1_1 gpc4042 (
      {stage0_34[406]},
      {stage1_34[162]}
   );
   gpc1_1 gpc4043 (
      {stage0_34[407]},
      {stage1_34[163]}
   );
   gpc1_1 gpc4044 (
      {stage0_34[408]},
      {stage1_34[164]}
   );
   gpc1_1 gpc4045 (
      {stage0_34[409]},
      {stage1_34[165]}
   );
   gpc1_1 gpc4046 (
      {stage0_34[410]},
      {stage1_34[166]}
   );
   gpc1_1 gpc4047 (
      {stage0_34[411]},
      {stage1_34[167]}
   );
   gpc1_1 gpc4048 (
      {stage0_34[412]},
      {stage1_34[168]}
   );
   gpc1_1 gpc4049 (
      {stage0_34[413]},
      {stage1_34[169]}
   );
   gpc1_1 gpc4050 (
      {stage0_34[414]},
      {stage1_34[170]}
   );
   gpc1_1 gpc4051 (
      {stage0_34[415]},
      {stage1_34[171]}
   );
   gpc1_1 gpc4052 (
      {stage0_34[416]},
      {stage1_34[172]}
   );
   gpc1_1 gpc4053 (
      {stage0_34[417]},
      {stage1_34[173]}
   );
   gpc1_1 gpc4054 (
      {stage0_34[418]},
      {stage1_34[174]}
   );
   gpc1_1 gpc4055 (
      {stage0_34[419]},
      {stage1_34[175]}
   );
   gpc1_1 gpc4056 (
      {stage0_34[420]},
      {stage1_34[176]}
   );
   gpc1_1 gpc4057 (
      {stage0_34[421]},
      {stage1_34[177]}
   );
   gpc1_1 gpc4058 (
      {stage0_34[422]},
      {stage1_34[178]}
   );
   gpc1_1 gpc4059 (
      {stage0_34[423]},
      {stage1_34[179]}
   );
   gpc1_1 gpc4060 (
      {stage0_34[424]},
      {stage1_34[180]}
   );
   gpc1_1 gpc4061 (
      {stage0_34[425]},
      {stage1_34[181]}
   );
   gpc1_1 gpc4062 (
      {stage0_34[426]},
      {stage1_34[182]}
   );
   gpc1_1 gpc4063 (
      {stage0_34[427]},
      {stage1_34[183]}
   );
   gpc1_1 gpc4064 (
      {stage0_34[428]},
      {stage1_34[184]}
   );
   gpc1_1 gpc4065 (
      {stage0_34[429]},
      {stage1_34[185]}
   );
   gpc1_1 gpc4066 (
      {stage0_34[430]},
      {stage1_34[186]}
   );
   gpc1_1 gpc4067 (
      {stage0_34[431]},
      {stage1_34[187]}
   );
   gpc1_1 gpc4068 (
      {stage0_34[432]},
      {stage1_34[188]}
   );
   gpc1_1 gpc4069 (
      {stage0_34[433]},
      {stage1_34[189]}
   );
   gpc1_1 gpc4070 (
      {stage0_34[434]},
      {stage1_34[190]}
   );
   gpc1_1 gpc4071 (
      {stage0_34[435]},
      {stage1_34[191]}
   );
   gpc1_1 gpc4072 (
      {stage0_34[436]},
      {stage1_34[192]}
   );
   gpc1_1 gpc4073 (
      {stage0_34[437]},
      {stage1_34[193]}
   );
   gpc1_1 gpc4074 (
      {stage0_34[438]},
      {stage1_34[194]}
   );
   gpc1_1 gpc4075 (
      {stage0_34[439]},
      {stage1_34[195]}
   );
   gpc1_1 gpc4076 (
      {stage0_34[440]},
      {stage1_34[196]}
   );
   gpc1_1 gpc4077 (
      {stage0_34[441]},
      {stage1_34[197]}
   );
   gpc1_1 gpc4078 (
      {stage0_34[442]},
      {stage1_34[198]}
   );
   gpc1_1 gpc4079 (
      {stage0_34[443]},
      {stage1_34[199]}
   );
   gpc1_1 gpc4080 (
      {stage0_34[444]},
      {stage1_34[200]}
   );
   gpc1_1 gpc4081 (
      {stage0_34[445]},
      {stage1_34[201]}
   );
   gpc1_1 gpc4082 (
      {stage0_34[446]},
      {stage1_34[202]}
   );
   gpc1_1 gpc4083 (
      {stage0_34[447]},
      {stage1_34[203]}
   );
   gpc1_1 gpc4084 (
      {stage0_34[448]},
      {stage1_34[204]}
   );
   gpc1_1 gpc4085 (
      {stage0_34[449]},
      {stage1_34[205]}
   );
   gpc1_1 gpc4086 (
      {stage0_34[450]},
      {stage1_34[206]}
   );
   gpc1_1 gpc4087 (
      {stage0_34[451]},
      {stage1_34[207]}
   );
   gpc1_1 gpc4088 (
      {stage0_34[452]},
      {stage1_34[208]}
   );
   gpc1_1 gpc4089 (
      {stage0_34[453]},
      {stage1_34[209]}
   );
   gpc1_1 gpc4090 (
      {stage0_34[454]},
      {stage1_34[210]}
   );
   gpc1_1 gpc4091 (
      {stage0_34[455]},
      {stage1_34[211]}
   );
   gpc1_1 gpc4092 (
      {stage0_34[456]},
      {stage1_34[212]}
   );
   gpc1_1 gpc4093 (
      {stage0_34[457]},
      {stage1_34[213]}
   );
   gpc1_1 gpc4094 (
      {stage0_34[458]},
      {stage1_34[214]}
   );
   gpc1_1 gpc4095 (
      {stage0_34[459]},
      {stage1_34[215]}
   );
   gpc1_1 gpc4096 (
      {stage0_34[460]},
      {stage1_34[216]}
   );
   gpc1_1 gpc4097 (
      {stage0_34[461]},
      {stage1_34[217]}
   );
   gpc1_1 gpc4098 (
      {stage0_34[462]},
      {stage1_34[218]}
   );
   gpc1_1 gpc4099 (
      {stage0_34[463]},
      {stage1_34[219]}
   );
   gpc1_1 gpc4100 (
      {stage0_34[464]},
      {stage1_34[220]}
   );
   gpc1_1 gpc4101 (
      {stage0_34[465]},
      {stage1_34[221]}
   );
   gpc1_1 gpc4102 (
      {stage0_34[466]},
      {stage1_34[222]}
   );
   gpc1_1 gpc4103 (
      {stage0_34[467]},
      {stage1_34[223]}
   );
   gpc1_1 gpc4104 (
      {stage0_34[468]},
      {stage1_34[224]}
   );
   gpc1_1 gpc4105 (
      {stage0_34[469]},
      {stage1_34[225]}
   );
   gpc1_1 gpc4106 (
      {stage0_34[470]},
      {stage1_34[226]}
   );
   gpc1_1 gpc4107 (
      {stage0_34[471]},
      {stage1_34[227]}
   );
   gpc1_1 gpc4108 (
      {stage0_34[472]},
      {stage1_34[228]}
   );
   gpc1_1 gpc4109 (
      {stage0_34[473]},
      {stage1_34[229]}
   );
   gpc1_1 gpc4110 (
      {stage0_34[474]},
      {stage1_34[230]}
   );
   gpc1_1 gpc4111 (
      {stage0_34[475]},
      {stage1_34[231]}
   );
   gpc1_1 gpc4112 (
      {stage0_34[476]},
      {stage1_34[232]}
   );
   gpc1_1 gpc4113 (
      {stage0_34[477]},
      {stage1_34[233]}
   );
   gpc1_1 gpc4114 (
      {stage0_34[478]},
      {stage1_34[234]}
   );
   gpc1_1 gpc4115 (
      {stage0_34[479]},
      {stage1_34[235]}
   );
   gpc1_1 gpc4116 (
      {stage0_34[480]},
      {stage1_34[236]}
   );
   gpc1_1 gpc4117 (
      {stage0_34[481]},
      {stage1_34[237]}
   );
   gpc1_1 gpc4118 (
      {stage0_34[482]},
      {stage1_34[238]}
   );
   gpc1_1 gpc4119 (
      {stage0_34[483]},
      {stage1_34[239]}
   );
   gpc1_1 gpc4120 (
      {stage0_34[484]},
      {stage1_34[240]}
   );
   gpc1_1 gpc4121 (
      {stage0_34[485]},
      {stage1_34[241]}
   );
   gpc1_1 gpc4122 (
      {stage0_34[486]},
      {stage1_34[242]}
   );
   gpc1_1 gpc4123 (
      {stage0_34[487]},
      {stage1_34[243]}
   );
   gpc1_1 gpc4124 (
      {stage0_34[488]},
      {stage1_34[244]}
   );
   gpc1_1 gpc4125 (
      {stage0_34[489]},
      {stage1_34[245]}
   );
   gpc1_1 gpc4126 (
      {stage0_34[490]},
      {stage1_34[246]}
   );
   gpc1_1 gpc4127 (
      {stage0_34[491]},
      {stage1_34[247]}
   );
   gpc1_1 gpc4128 (
      {stage0_34[492]},
      {stage1_34[248]}
   );
   gpc1_1 gpc4129 (
      {stage0_34[493]},
      {stage1_34[249]}
   );
   gpc1_1 gpc4130 (
      {stage0_34[494]},
      {stage1_34[250]}
   );
   gpc1_1 gpc4131 (
      {stage0_34[495]},
      {stage1_34[251]}
   );
   gpc1_1 gpc4132 (
      {stage0_34[496]},
      {stage1_34[252]}
   );
   gpc1_1 gpc4133 (
      {stage0_34[497]},
      {stage1_34[253]}
   );
   gpc1_1 gpc4134 (
      {stage0_34[498]},
      {stage1_34[254]}
   );
   gpc1_1 gpc4135 (
      {stage0_34[499]},
      {stage1_34[255]}
   );
   gpc1_1 gpc4136 (
      {stage0_34[500]},
      {stage1_34[256]}
   );
   gpc1_1 gpc4137 (
      {stage0_34[501]},
      {stage1_34[257]}
   );
   gpc1_1 gpc4138 (
      {stage0_34[502]},
      {stage1_34[258]}
   );
   gpc1_1 gpc4139 (
      {stage0_34[503]},
      {stage1_34[259]}
   );
   gpc1_1 gpc4140 (
      {stage0_34[504]},
      {stage1_34[260]}
   );
   gpc1_1 gpc4141 (
      {stage0_34[505]},
      {stage1_34[261]}
   );
   gpc1_1 gpc4142 (
      {stage0_34[506]},
      {stage1_34[262]}
   );
   gpc1_1 gpc4143 (
      {stage0_34[507]},
      {stage1_34[263]}
   );
   gpc1_1 gpc4144 (
      {stage0_34[508]},
      {stage1_34[264]}
   );
   gpc1_1 gpc4145 (
      {stage0_34[509]},
      {stage1_34[265]}
   );
   gpc1_1 gpc4146 (
      {stage0_34[510]},
      {stage1_34[266]}
   );
   gpc1_1 gpc4147 (
      {stage0_34[511]},
      {stage1_34[267]}
   );
   gpc1_1 gpc4148 (
      {stage0_35[495]},
      {stage1_35[174]}
   );
   gpc1_1 gpc4149 (
      {stage0_35[496]},
      {stage1_35[175]}
   );
   gpc1_1 gpc4150 (
      {stage0_35[497]},
      {stage1_35[176]}
   );
   gpc1_1 gpc4151 (
      {stage0_35[498]},
      {stage1_35[177]}
   );
   gpc1_1 gpc4152 (
      {stage0_35[499]},
      {stage1_35[178]}
   );
   gpc1_1 gpc4153 (
      {stage0_35[500]},
      {stage1_35[179]}
   );
   gpc1_1 gpc4154 (
      {stage0_35[501]},
      {stage1_35[180]}
   );
   gpc1_1 gpc4155 (
      {stage0_35[502]},
      {stage1_35[181]}
   );
   gpc1_1 gpc4156 (
      {stage0_35[503]},
      {stage1_35[182]}
   );
   gpc1_1 gpc4157 (
      {stage0_35[504]},
      {stage1_35[183]}
   );
   gpc1_1 gpc4158 (
      {stage0_35[505]},
      {stage1_35[184]}
   );
   gpc1_1 gpc4159 (
      {stage0_35[506]},
      {stage1_35[185]}
   );
   gpc1_1 gpc4160 (
      {stage0_35[507]},
      {stage1_35[186]}
   );
   gpc1_1 gpc4161 (
      {stage0_35[508]},
      {stage1_35[187]}
   );
   gpc1_1 gpc4162 (
      {stage0_35[509]},
      {stage1_35[188]}
   );
   gpc1_1 gpc4163 (
      {stage0_35[510]},
      {stage1_35[189]}
   );
   gpc1_1 gpc4164 (
      {stage0_35[511]},
      {stage1_35[190]}
   );
   gpc1_1 gpc4165 (
      {stage0_36[367]},
      {stage1_36[186]}
   );
   gpc1_1 gpc4166 (
      {stage0_36[368]},
      {stage1_36[187]}
   );
   gpc1_1 gpc4167 (
      {stage0_36[369]},
      {stage1_36[188]}
   );
   gpc1_1 gpc4168 (
      {stage0_36[370]},
      {stage1_36[189]}
   );
   gpc1_1 gpc4169 (
      {stage0_36[371]},
      {stage1_36[190]}
   );
   gpc1_1 gpc4170 (
      {stage0_36[372]},
      {stage1_36[191]}
   );
   gpc1_1 gpc4171 (
      {stage0_36[373]},
      {stage1_36[192]}
   );
   gpc1_1 gpc4172 (
      {stage0_36[374]},
      {stage1_36[193]}
   );
   gpc1_1 gpc4173 (
      {stage0_36[375]},
      {stage1_36[194]}
   );
   gpc1_1 gpc4174 (
      {stage0_36[376]},
      {stage1_36[195]}
   );
   gpc1_1 gpc4175 (
      {stage0_36[377]},
      {stage1_36[196]}
   );
   gpc1_1 gpc4176 (
      {stage0_36[378]},
      {stage1_36[197]}
   );
   gpc1_1 gpc4177 (
      {stage0_36[379]},
      {stage1_36[198]}
   );
   gpc1_1 gpc4178 (
      {stage0_36[380]},
      {stage1_36[199]}
   );
   gpc1_1 gpc4179 (
      {stage0_36[381]},
      {stage1_36[200]}
   );
   gpc1_1 gpc4180 (
      {stage0_36[382]},
      {stage1_36[201]}
   );
   gpc1_1 gpc4181 (
      {stage0_36[383]},
      {stage1_36[202]}
   );
   gpc1_1 gpc4182 (
      {stage0_36[384]},
      {stage1_36[203]}
   );
   gpc1_1 gpc4183 (
      {stage0_36[385]},
      {stage1_36[204]}
   );
   gpc1_1 gpc4184 (
      {stage0_36[386]},
      {stage1_36[205]}
   );
   gpc1_1 gpc4185 (
      {stage0_36[387]},
      {stage1_36[206]}
   );
   gpc1_1 gpc4186 (
      {stage0_36[388]},
      {stage1_36[207]}
   );
   gpc1_1 gpc4187 (
      {stage0_36[389]},
      {stage1_36[208]}
   );
   gpc1_1 gpc4188 (
      {stage0_36[390]},
      {stage1_36[209]}
   );
   gpc1_1 gpc4189 (
      {stage0_36[391]},
      {stage1_36[210]}
   );
   gpc1_1 gpc4190 (
      {stage0_36[392]},
      {stage1_36[211]}
   );
   gpc1_1 gpc4191 (
      {stage0_36[393]},
      {stage1_36[212]}
   );
   gpc1_1 gpc4192 (
      {stage0_36[394]},
      {stage1_36[213]}
   );
   gpc1_1 gpc4193 (
      {stage0_36[395]},
      {stage1_36[214]}
   );
   gpc1_1 gpc4194 (
      {stage0_36[396]},
      {stage1_36[215]}
   );
   gpc1_1 gpc4195 (
      {stage0_36[397]},
      {stage1_36[216]}
   );
   gpc1_1 gpc4196 (
      {stage0_36[398]},
      {stage1_36[217]}
   );
   gpc1_1 gpc4197 (
      {stage0_36[399]},
      {stage1_36[218]}
   );
   gpc1_1 gpc4198 (
      {stage0_36[400]},
      {stage1_36[219]}
   );
   gpc1_1 gpc4199 (
      {stage0_36[401]},
      {stage1_36[220]}
   );
   gpc1_1 gpc4200 (
      {stage0_36[402]},
      {stage1_36[221]}
   );
   gpc1_1 gpc4201 (
      {stage0_36[403]},
      {stage1_36[222]}
   );
   gpc1_1 gpc4202 (
      {stage0_36[404]},
      {stage1_36[223]}
   );
   gpc1_1 gpc4203 (
      {stage0_36[405]},
      {stage1_36[224]}
   );
   gpc1_1 gpc4204 (
      {stage0_36[406]},
      {stage1_36[225]}
   );
   gpc1_1 gpc4205 (
      {stage0_36[407]},
      {stage1_36[226]}
   );
   gpc1_1 gpc4206 (
      {stage0_36[408]},
      {stage1_36[227]}
   );
   gpc1_1 gpc4207 (
      {stage0_36[409]},
      {stage1_36[228]}
   );
   gpc1_1 gpc4208 (
      {stage0_36[410]},
      {stage1_36[229]}
   );
   gpc1_1 gpc4209 (
      {stage0_36[411]},
      {stage1_36[230]}
   );
   gpc1_1 gpc4210 (
      {stage0_36[412]},
      {stage1_36[231]}
   );
   gpc1_1 gpc4211 (
      {stage0_36[413]},
      {stage1_36[232]}
   );
   gpc1_1 gpc4212 (
      {stage0_36[414]},
      {stage1_36[233]}
   );
   gpc1_1 gpc4213 (
      {stage0_36[415]},
      {stage1_36[234]}
   );
   gpc1_1 gpc4214 (
      {stage0_36[416]},
      {stage1_36[235]}
   );
   gpc1_1 gpc4215 (
      {stage0_36[417]},
      {stage1_36[236]}
   );
   gpc1_1 gpc4216 (
      {stage0_36[418]},
      {stage1_36[237]}
   );
   gpc1_1 gpc4217 (
      {stage0_36[419]},
      {stage1_36[238]}
   );
   gpc1_1 gpc4218 (
      {stage0_36[420]},
      {stage1_36[239]}
   );
   gpc1_1 gpc4219 (
      {stage0_36[421]},
      {stage1_36[240]}
   );
   gpc1_1 gpc4220 (
      {stage0_36[422]},
      {stage1_36[241]}
   );
   gpc1_1 gpc4221 (
      {stage0_36[423]},
      {stage1_36[242]}
   );
   gpc1_1 gpc4222 (
      {stage0_36[424]},
      {stage1_36[243]}
   );
   gpc1_1 gpc4223 (
      {stage0_36[425]},
      {stage1_36[244]}
   );
   gpc1_1 gpc4224 (
      {stage0_36[426]},
      {stage1_36[245]}
   );
   gpc1_1 gpc4225 (
      {stage0_36[427]},
      {stage1_36[246]}
   );
   gpc1_1 gpc4226 (
      {stage0_36[428]},
      {stage1_36[247]}
   );
   gpc1_1 gpc4227 (
      {stage0_36[429]},
      {stage1_36[248]}
   );
   gpc1_1 gpc4228 (
      {stage0_36[430]},
      {stage1_36[249]}
   );
   gpc1_1 gpc4229 (
      {stage0_36[431]},
      {stage1_36[250]}
   );
   gpc1_1 gpc4230 (
      {stage0_36[432]},
      {stage1_36[251]}
   );
   gpc1_1 gpc4231 (
      {stage0_36[433]},
      {stage1_36[252]}
   );
   gpc1_1 gpc4232 (
      {stage0_36[434]},
      {stage1_36[253]}
   );
   gpc1_1 gpc4233 (
      {stage0_36[435]},
      {stage1_36[254]}
   );
   gpc1_1 gpc4234 (
      {stage0_36[436]},
      {stage1_36[255]}
   );
   gpc1_1 gpc4235 (
      {stage0_36[437]},
      {stage1_36[256]}
   );
   gpc1_1 gpc4236 (
      {stage0_36[438]},
      {stage1_36[257]}
   );
   gpc1_1 gpc4237 (
      {stage0_36[439]},
      {stage1_36[258]}
   );
   gpc1_1 gpc4238 (
      {stage0_36[440]},
      {stage1_36[259]}
   );
   gpc1_1 gpc4239 (
      {stage0_36[441]},
      {stage1_36[260]}
   );
   gpc1_1 gpc4240 (
      {stage0_36[442]},
      {stage1_36[261]}
   );
   gpc1_1 gpc4241 (
      {stage0_36[443]},
      {stage1_36[262]}
   );
   gpc1_1 gpc4242 (
      {stage0_36[444]},
      {stage1_36[263]}
   );
   gpc1_1 gpc4243 (
      {stage0_36[445]},
      {stage1_36[264]}
   );
   gpc1_1 gpc4244 (
      {stage0_36[446]},
      {stage1_36[265]}
   );
   gpc1_1 gpc4245 (
      {stage0_36[447]},
      {stage1_36[266]}
   );
   gpc1_1 gpc4246 (
      {stage0_36[448]},
      {stage1_36[267]}
   );
   gpc1_1 gpc4247 (
      {stage0_36[449]},
      {stage1_36[268]}
   );
   gpc1_1 gpc4248 (
      {stage0_36[450]},
      {stage1_36[269]}
   );
   gpc1_1 gpc4249 (
      {stage0_36[451]},
      {stage1_36[270]}
   );
   gpc1_1 gpc4250 (
      {stage0_36[452]},
      {stage1_36[271]}
   );
   gpc1_1 gpc4251 (
      {stage0_36[453]},
      {stage1_36[272]}
   );
   gpc1_1 gpc4252 (
      {stage0_36[454]},
      {stage1_36[273]}
   );
   gpc1_1 gpc4253 (
      {stage0_36[455]},
      {stage1_36[274]}
   );
   gpc1_1 gpc4254 (
      {stage0_36[456]},
      {stage1_36[275]}
   );
   gpc1_1 gpc4255 (
      {stage0_36[457]},
      {stage1_36[276]}
   );
   gpc1_1 gpc4256 (
      {stage0_36[458]},
      {stage1_36[277]}
   );
   gpc1_1 gpc4257 (
      {stage0_36[459]},
      {stage1_36[278]}
   );
   gpc1_1 gpc4258 (
      {stage0_36[460]},
      {stage1_36[279]}
   );
   gpc1_1 gpc4259 (
      {stage0_36[461]},
      {stage1_36[280]}
   );
   gpc1_1 gpc4260 (
      {stage0_36[462]},
      {stage1_36[281]}
   );
   gpc1_1 gpc4261 (
      {stage0_36[463]},
      {stage1_36[282]}
   );
   gpc1_1 gpc4262 (
      {stage0_36[464]},
      {stage1_36[283]}
   );
   gpc1_1 gpc4263 (
      {stage0_36[465]},
      {stage1_36[284]}
   );
   gpc1_1 gpc4264 (
      {stage0_36[466]},
      {stage1_36[285]}
   );
   gpc1_1 gpc4265 (
      {stage0_36[467]},
      {stage1_36[286]}
   );
   gpc1_1 gpc4266 (
      {stage0_36[468]},
      {stage1_36[287]}
   );
   gpc1_1 gpc4267 (
      {stage0_36[469]},
      {stage1_36[288]}
   );
   gpc1_1 gpc4268 (
      {stage0_36[470]},
      {stage1_36[289]}
   );
   gpc1_1 gpc4269 (
      {stage0_36[471]},
      {stage1_36[290]}
   );
   gpc1_1 gpc4270 (
      {stage0_36[472]},
      {stage1_36[291]}
   );
   gpc1_1 gpc4271 (
      {stage0_36[473]},
      {stage1_36[292]}
   );
   gpc1_1 gpc4272 (
      {stage0_36[474]},
      {stage1_36[293]}
   );
   gpc1_1 gpc4273 (
      {stage0_36[475]},
      {stage1_36[294]}
   );
   gpc1_1 gpc4274 (
      {stage0_36[476]},
      {stage1_36[295]}
   );
   gpc1_1 gpc4275 (
      {stage0_36[477]},
      {stage1_36[296]}
   );
   gpc1_1 gpc4276 (
      {stage0_36[478]},
      {stage1_36[297]}
   );
   gpc1_1 gpc4277 (
      {stage0_36[479]},
      {stage1_36[298]}
   );
   gpc1_1 gpc4278 (
      {stage0_36[480]},
      {stage1_36[299]}
   );
   gpc1_1 gpc4279 (
      {stage0_36[481]},
      {stage1_36[300]}
   );
   gpc1_1 gpc4280 (
      {stage0_36[482]},
      {stage1_36[301]}
   );
   gpc1_1 gpc4281 (
      {stage0_36[483]},
      {stage1_36[302]}
   );
   gpc1_1 gpc4282 (
      {stage0_36[484]},
      {stage1_36[303]}
   );
   gpc1_1 gpc4283 (
      {stage0_36[485]},
      {stage1_36[304]}
   );
   gpc1_1 gpc4284 (
      {stage0_36[486]},
      {stage1_36[305]}
   );
   gpc1_1 gpc4285 (
      {stage0_36[487]},
      {stage1_36[306]}
   );
   gpc1_1 gpc4286 (
      {stage0_36[488]},
      {stage1_36[307]}
   );
   gpc1_1 gpc4287 (
      {stage0_36[489]},
      {stage1_36[308]}
   );
   gpc1_1 gpc4288 (
      {stage0_36[490]},
      {stage1_36[309]}
   );
   gpc1_1 gpc4289 (
      {stage0_36[491]},
      {stage1_36[310]}
   );
   gpc1_1 gpc4290 (
      {stage0_36[492]},
      {stage1_36[311]}
   );
   gpc1_1 gpc4291 (
      {stage0_36[493]},
      {stage1_36[312]}
   );
   gpc1_1 gpc4292 (
      {stage0_36[494]},
      {stage1_36[313]}
   );
   gpc1_1 gpc4293 (
      {stage0_36[495]},
      {stage1_36[314]}
   );
   gpc1_1 gpc4294 (
      {stage0_36[496]},
      {stage1_36[315]}
   );
   gpc1_1 gpc4295 (
      {stage0_36[497]},
      {stage1_36[316]}
   );
   gpc1_1 gpc4296 (
      {stage0_36[498]},
      {stage1_36[317]}
   );
   gpc1_1 gpc4297 (
      {stage0_36[499]},
      {stage1_36[318]}
   );
   gpc1_1 gpc4298 (
      {stage0_36[500]},
      {stage1_36[319]}
   );
   gpc1_1 gpc4299 (
      {stage0_36[501]},
      {stage1_36[320]}
   );
   gpc1_1 gpc4300 (
      {stage0_36[502]},
      {stage1_36[321]}
   );
   gpc1_1 gpc4301 (
      {stage0_36[503]},
      {stage1_36[322]}
   );
   gpc1_1 gpc4302 (
      {stage0_36[504]},
      {stage1_36[323]}
   );
   gpc1_1 gpc4303 (
      {stage0_36[505]},
      {stage1_36[324]}
   );
   gpc1_1 gpc4304 (
      {stage0_36[506]},
      {stage1_36[325]}
   );
   gpc1_1 gpc4305 (
      {stage0_36[507]},
      {stage1_36[326]}
   );
   gpc1_1 gpc4306 (
      {stage0_36[508]},
      {stage1_36[327]}
   );
   gpc1_1 gpc4307 (
      {stage0_36[509]},
      {stage1_36[328]}
   );
   gpc1_1 gpc4308 (
      {stage0_36[510]},
      {stage1_36[329]}
   );
   gpc1_1 gpc4309 (
      {stage0_36[511]},
      {stage1_36[330]}
   );
   gpc1_1 gpc4310 (
      {stage0_37[392]},
      {stage1_37[183]}
   );
   gpc1_1 gpc4311 (
      {stage0_37[393]},
      {stage1_37[184]}
   );
   gpc1_1 gpc4312 (
      {stage0_37[394]},
      {stage1_37[185]}
   );
   gpc1_1 gpc4313 (
      {stage0_37[395]},
      {stage1_37[186]}
   );
   gpc1_1 gpc4314 (
      {stage0_37[396]},
      {stage1_37[187]}
   );
   gpc1_1 gpc4315 (
      {stage0_37[397]},
      {stage1_37[188]}
   );
   gpc1_1 gpc4316 (
      {stage0_37[398]},
      {stage1_37[189]}
   );
   gpc1_1 gpc4317 (
      {stage0_37[399]},
      {stage1_37[190]}
   );
   gpc1_1 gpc4318 (
      {stage0_37[400]},
      {stage1_37[191]}
   );
   gpc1_1 gpc4319 (
      {stage0_37[401]},
      {stage1_37[192]}
   );
   gpc1_1 gpc4320 (
      {stage0_37[402]},
      {stage1_37[193]}
   );
   gpc1_1 gpc4321 (
      {stage0_37[403]},
      {stage1_37[194]}
   );
   gpc1_1 gpc4322 (
      {stage0_37[404]},
      {stage1_37[195]}
   );
   gpc1_1 gpc4323 (
      {stage0_37[405]},
      {stage1_37[196]}
   );
   gpc1_1 gpc4324 (
      {stage0_37[406]},
      {stage1_37[197]}
   );
   gpc1_1 gpc4325 (
      {stage0_37[407]},
      {stage1_37[198]}
   );
   gpc1_1 gpc4326 (
      {stage0_37[408]},
      {stage1_37[199]}
   );
   gpc1_1 gpc4327 (
      {stage0_37[409]},
      {stage1_37[200]}
   );
   gpc1_1 gpc4328 (
      {stage0_37[410]},
      {stage1_37[201]}
   );
   gpc1_1 gpc4329 (
      {stage0_37[411]},
      {stage1_37[202]}
   );
   gpc1_1 gpc4330 (
      {stage0_37[412]},
      {stage1_37[203]}
   );
   gpc1_1 gpc4331 (
      {stage0_37[413]},
      {stage1_37[204]}
   );
   gpc1_1 gpc4332 (
      {stage0_37[414]},
      {stage1_37[205]}
   );
   gpc1_1 gpc4333 (
      {stage0_37[415]},
      {stage1_37[206]}
   );
   gpc1_1 gpc4334 (
      {stage0_37[416]},
      {stage1_37[207]}
   );
   gpc1_1 gpc4335 (
      {stage0_37[417]},
      {stage1_37[208]}
   );
   gpc1_1 gpc4336 (
      {stage0_37[418]},
      {stage1_37[209]}
   );
   gpc1_1 gpc4337 (
      {stage0_37[419]},
      {stage1_37[210]}
   );
   gpc1_1 gpc4338 (
      {stage0_37[420]},
      {stage1_37[211]}
   );
   gpc1_1 gpc4339 (
      {stage0_37[421]},
      {stage1_37[212]}
   );
   gpc1_1 gpc4340 (
      {stage0_37[422]},
      {stage1_37[213]}
   );
   gpc1_1 gpc4341 (
      {stage0_37[423]},
      {stage1_37[214]}
   );
   gpc1_1 gpc4342 (
      {stage0_37[424]},
      {stage1_37[215]}
   );
   gpc1_1 gpc4343 (
      {stage0_37[425]},
      {stage1_37[216]}
   );
   gpc1_1 gpc4344 (
      {stage0_37[426]},
      {stage1_37[217]}
   );
   gpc1_1 gpc4345 (
      {stage0_37[427]},
      {stage1_37[218]}
   );
   gpc1_1 gpc4346 (
      {stage0_37[428]},
      {stage1_37[219]}
   );
   gpc1_1 gpc4347 (
      {stage0_37[429]},
      {stage1_37[220]}
   );
   gpc1_1 gpc4348 (
      {stage0_37[430]},
      {stage1_37[221]}
   );
   gpc1_1 gpc4349 (
      {stage0_37[431]},
      {stage1_37[222]}
   );
   gpc1_1 gpc4350 (
      {stage0_37[432]},
      {stage1_37[223]}
   );
   gpc1_1 gpc4351 (
      {stage0_37[433]},
      {stage1_37[224]}
   );
   gpc1_1 gpc4352 (
      {stage0_37[434]},
      {stage1_37[225]}
   );
   gpc1_1 gpc4353 (
      {stage0_37[435]},
      {stage1_37[226]}
   );
   gpc1_1 gpc4354 (
      {stage0_37[436]},
      {stage1_37[227]}
   );
   gpc1_1 gpc4355 (
      {stage0_37[437]},
      {stage1_37[228]}
   );
   gpc1_1 gpc4356 (
      {stage0_37[438]},
      {stage1_37[229]}
   );
   gpc1_1 gpc4357 (
      {stage0_37[439]},
      {stage1_37[230]}
   );
   gpc1_1 gpc4358 (
      {stage0_37[440]},
      {stage1_37[231]}
   );
   gpc1_1 gpc4359 (
      {stage0_37[441]},
      {stage1_37[232]}
   );
   gpc1_1 gpc4360 (
      {stage0_37[442]},
      {stage1_37[233]}
   );
   gpc1_1 gpc4361 (
      {stage0_37[443]},
      {stage1_37[234]}
   );
   gpc1_1 gpc4362 (
      {stage0_37[444]},
      {stage1_37[235]}
   );
   gpc1_1 gpc4363 (
      {stage0_37[445]},
      {stage1_37[236]}
   );
   gpc1_1 gpc4364 (
      {stage0_37[446]},
      {stage1_37[237]}
   );
   gpc1_1 gpc4365 (
      {stage0_37[447]},
      {stage1_37[238]}
   );
   gpc1_1 gpc4366 (
      {stage0_37[448]},
      {stage1_37[239]}
   );
   gpc1_1 gpc4367 (
      {stage0_37[449]},
      {stage1_37[240]}
   );
   gpc1_1 gpc4368 (
      {stage0_37[450]},
      {stage1_37[241]}
   );
   gpc1_1 gpc4369 (
      {stage0_37[451]},
      {stage1_37[242]}
   );
   gpc1_1 gpc4370 (
      {stage0_37[452]},
      {stage1_37[243]}
   );
   gpc1_1 gpc4371 (
      {stage0_37[453]},
      {stage1_37[244]}
   );
   gpc1_1 gpc4372 (
      {stage0_37[454]},
      {stage1_37[245]}
   );
   gpc1_1 gpc4373 (
      {stage0_37[455]},
      {stage1_37[246]}
   );
   gpc1_1 gpc4374 (
      {stage0_37[456]},
      {stage1_37[247]}
   );
   gpc1_1 gpc4375 (
      {stage0_37[457]},
      {stage1_37[248]}
   );
   gpc1_1 gpc4376 (
      {stage0_37[458]},
      {stage1_37[249]}
   );
   gpc1_1 gpc4377 (
      {stage0_37[459]},
      {stage1_37[250]}
   );
   gpc1_1 gpc4378 (
      {stage0_37[460]},
      {stage1_37[251]}
   );
   gpc1_1 gpc4379 (
      {stage0_37[461]},
      {stage1_37[252]}
   );
   gpc1_1 gpc4380 (
      {stage0_37[462]},
      {stage1_37[253]}
   );
   gpc1_1 gpc4381 (
      {stage0_37[463]},
      {stage1_37[254]}
   );
   gpc1_1 gpc4382 (
      {stage0_37[464]},
      {stage1_37[255]}
   );
   gpc1_1 gpc4383 (
      {stage0_37[465]},
      {stage1_37[256]}
   );
   gpc1_1 gpc4384 (
      {stage0_37[466]},
      {stage1_37[257]}
   );
   gpc1_1 gpc4385 (
      {stage0_37[467]},
      {stage1_37[258]}
   );
   gpc1_1 gpc4386 (
      {stage0_37[468]},
      {stage1_37[259]}
   );
   gpc1_1 gpc4387 (
      {stage0_37[469]},
      {stage1_37[260]}
   );
   gpc1_1 gpc4388 (
      {stage0_37[470]},
      {stage1_37[261]}
   );
   gpc1_1 gpc4389 (
      {stage0_37[471]},
      {stage1_37[262]}
   );
   gpc1_1 gpc4390 (
      {stage0_37[472]},
      {stage1_37[263]}
   );
   gpc1_1 gpc4391 (
      {stage0_37[473]},
      {stage1_37[264]}
   );
   gpc1_1 gpc4392 (
      {stage0_37[474]},
      {stage1_37[265]}
   );
   gpc1_1 gpc4393 (
      {stage0_37[475]},
      {stage1_37[266]}
   );
   gpc1_1 gpc4394 (
      {stage0_37[476]},
      {stage1_37[267]}
   );
   gpc1_1 gpc4395 (
      {stage0_37[477]},
      {stage1_37[268]}
   );
   gpc1_1 gpc4396 (
      {stage0_37[478]},
      {stage1_37[269]}
   );
   gpc1_1 gpc4397 (
      {stage0_37[479]},
      {stage1_37[270]}
   );
   gpc1_1 gpc4398 (
      {stage0_37[480]},
      {stage1_37[271]}
   );
   gpc1_1 gpc4399 (
      {stage0_37[481]},
      {stage1_37[272]}
   );
   gpc1_1 gpc4400 (
      {stage0_37[482]},
      {stage1_37[273]}
   );
   gpc1_1 gpc4401 (
      {stage0_37[483]},
      {stage1_37[274]}
   );
   gpc1_1 gpc4402 (
      {stage0_37[484]},
      {stage1_37[275]}
   );
   gpc1_1 gpc4403 (
      {stage0_37[485]},
      {stage1_37[276]}
   );
   gpc1_1 gpc4404 (
      {stage0_37[486]},
      {stage1_37[277]}
   );
   gpc1_1 gpc4405 (
      {stage0_37[487]},
      {stage1_37[278]}
   );
   gpc1_1 gpc4406 (
      {stage0_37[488]},
      {stage1_37[279]}
   );
   gpc1_1 gpc4407 (
      {stage0_37[489]},
      {stage1_37[280]}
   );
   gpc1_1 gpc4408 (
      {stage0_37[490]},
      {stage1_37[281]}
   );
   gpc1_1 gpc4409 (
      {stage0_37[491]},
      {stage1_37[282]}
   );
   gpc1_1 gpc4410 (
      {stage0_37[492]},
      {stage1_37[283]}
   );
   gpc1_1 gpc4411 (
      {stage0_37[493]},
      {stage1_37[284]}
   );
   gpc1_1 gpc4412 (
      {stage0_37[494]},
      {stage1_37[285]}
   );
   gpc1_1 gpc4413 (
      {stage0_37[495]},
      {stage1_37[286]}
   );
   gpc1_1 gpc4414 (
      {stage0_37[496]},
      {stage1_37[287]}
   );
   gpc1_1 gpc4415 (
      {stage0_37[497]},
      {stage1_37[288]}
   );
   gpc1_1 gpc4416 (
      {stage0_37[498]},
      {stage1_37[289]}
   );
   gpc1_1 gpc4417 (
      {stage0_37[499]},
      {stage1_37[290]}
   );
   gpc1_1 gpc4418 (
      {stage0_37[500]},
      {stage1_37[291]}
   );
   gpc1_1 gpc4419 (
      {stage0_37[501]},
      {stage1_37[292]}
   );
   gpc1_1 gpc4420 (
      {stage0_37[502]},
      {stage1_37[293]}
   );
   gpc1_1 gpc4421 (
      {stage0_37[503]},
      {stage1_37[294]}
   );
   gpc1_1 gpc4422 (
      {stage0_37[504]},
      {stage1_37[295]}
   );
   gpc1_1 gpc4423 (
      {stage0_37[505]},
      {stage1_37[296]}
   );
   gpc1_1 gpc4424 (
      {stage0_37[506]},
      {stage1_37[297]}
   );
   gpc1_1 gpc4425 (
      {stage0_37[507]},
      {stage1_37[298]}
   );
   gpc1_1 gpc4426 (
      {stage0_37[508]},
      {stage1_37[299]}
   );
   gpc1_1 gpc4427 (
      {stage0_37[509]},
      {stage1_37[300]}
   );
   gpc1_1 gpc4428 (
      {stage0_37[510]},
      {stage1_37[301]}
   );
   gpc1_1 gpc4429 (
      {stage0_37[511]},
      {stage1_37[302]}
   );
   gpc1_1 gpc4430 (
      {stage0_38[382]},
      {stage1_38[147]}
   );
   gpc1_1 gpc4431 (
      {stage0_38[383]},
      {stage1_38[148]}
   );
   gpc1_1 gpc4432 (
      {stage0_38[384]},
      {stage1_38[149]}
   );
   gpc1_1 gpc4433 (
      {stage0_38[385]},
      {stage1_38[150]}
   );
   gpc1_1 gpc4434 (
      {stage0_38[386]},
      {stage1_38[151]}
   );
   gpc1_1 gpc4435 (
      {stage0_38[387]},
      {stage1_38[152]}
   );
   gpc1_1 gpc4436 (
      {stage0_38[388]},
      {stage1_38[153]}
   );
   gpc1_1 gpc4437 (
      {stage0_38[389]},
      {stage1_38[154]}
   );
   gpc1_1 gpc4438 (
      {stage0_38[390]},
      {stage1_38[155]}
   );
   gpc1_1 gpc4439 (
      {stage0_38[391]},
      {stage1_38[156]}
   );
   gpc1_1 gpc4440 (
      {stage0_38[392]},
      {stage1_38[157]}
   );
   gpc1_1 gpc4441 (
      {stage0_38[393]},
      {stage1_38[158]}
   );
   gpc1_1 gpc4442 (
      {stage0_38[394]},
      {stage1_38[159]}
   );
   gpc1_1 gpc4443 (
      {stage0_38[395]},
      {stage1_38[160]}
   );
   gpc1_1 gpc4444 (
      {stage0_38[396]},
      {stage1_38[161]}
   );
   gpc1_1 gpc4445 (
      {stage0_38[397]},
      {stage1_38[162]}
   );
   gpc1_1 gpc4446 (
      {stage0_38[398]},
      {stage1_38[163]}
   );
   gpc1_1 gpc4447 (
      {stage0_38[399]},
      {stage1_38[164]}
   );
   gpc1_1 gpc4448 (
      {stage0_38[400]},
      {stage1_38[165]}
   );
   gpc1_1 gpc4449 (
      {stage0_38[401]},
      {stage1_38[166]}
   );
   gpc1_1 gpc4450 (
      {stage0_38[402]},
      {stage1_38[167]}
   );
   gpc1_1 gpc4451 (
      {stage0_38[403]},
      {stage1_38[168]}
   );
   gpc1_1 gpc4452 (
      {stage0_38[404]},
      {stage1_38[169]}
   );
   gpc1_1 gpc4453 (
      {stage0_38[405]},
      {stage1_38[170]}
   );
   gpc1_1 gpc4454 (
      {stage0_38[406]},
      {stage1_38[171]}
   );
   gpc1_1 gpc4455 (
      {stage0_38[407]},
      {stage1_38[172]}
   );
   gpc1_1 gpc4456 (
      {stage0_38[408]},
      {stage1_38[173]}
   );
   gpc1_1 gpc4457 (
      {stage0_38[409]},
      {stage1_38[174]}
   );
   gpc1_1 gpc4458 (
      {stage0_38[410]},
      {stage1_38[175]}
   );
   gpc1_1 gpc4459 (
      {stage0_38[411]},
      {stage1_38[176]}
   );
   gpc1_1 gpc4460 (
      {stage0_38[412]},
      {stage1_38[177]}
   );
   gpc1_1 gpc4461 (
      {stage0_38[413]},
      {stage1_38[178]}
   );
   gpc1_1 gpc4462 (
      {stage0_38[414]},
      {stage1_38[179]}
   );
   gpc1_1 gpc4463 (
      {stage0_38[415]},
      {stage1_38[180]}
   );
   gpc1_1 gpc4464 (
      {stage0_38[416]},
      {stage1_38[181]}
   );
   gpc1_1 gpc4465 (
      {stage0_38[417]},
      {stage1_38[182]}
   );
   gpc1_1 gpc4466 (
      {stage0_38[418]},
      {stage1_38[183]}
   );
   gpc1_1 gpc4467 (
      {stage0_38[419]},
      {stage1_38[184]}
   );
   gpc1_1 gpc4468 (
      {stage0_38[420]},
      {stage1_38[185]}
   );
   gpc1_1 gpc4469 (
      {stage0_38[421]},
      {stage1_38[186]}
   );
   gpc1_1 gpc4470 (
      {stage0_38[422]},
      {stage1_38[187]}
   );
   gpc1_1 gpc4471 (
      {stage0_38[423]},
      {stage1_38[188]}
   );
   gpc1_1 gpc4472 (
      {stage0_38[424]},
      {stage1_38[189]}
   );
   gpc1_1 gpc4473 (
      {stage0_38[425]},
      {stage1_38[190]}
   );
   gpc1_1 gpc4474 (
      {stage0_38[426]},
      {stage1_38[191]}
   );
   gpc1_1 gpc4475 (
      {stage0_38[427]},
      {stage1_38[192]}
   );
   gpc1_1 gpc4476 (
      {stage0_38[428]},
      {stage1_38[193]}
   );
   gpc1_1 gpc4477 (
      {stage0_38[429]},
      {stage1_38[194]}
   );
   gpc1_1 gpc4478 (
      {stage0_38[430]},
      {stage1_38[195]}
   );
   gpc1_1 gpc4479 (
      {stage0_38[431]},
      {stage1_38[196]}
   );
   gpc1_1 gpc4480 (
      {stage0_38[432]},
      {stage1_38[197]}
   );
   gpc1_1 gpc4481 (
      {stage0_38[433]},
      {stage1_38[198]}
   );
   gpc1_1 gpc4482 (
      {stage0_38[434]},
      {stage1_38[199]}
   );
   gpc1_1 gpc4483 (
      {stage0_38[435]},
      {stage1_38[200]}
   );
   gpc1_1 gpc4484 (
      {stage0_38[436]},
      {stage1_38[201]}
   );
   gpc1_1 gpc4485 (
      {stage0_38[437]},
      {stage1_38[202]}
   );
   gpc1_1 gpc4486 (
      {stage0_38[438]},
      {stage1_38[203]}
   );
   gpc1_1 gpc4487 (
      {stage0_38[439]},
      {stage1_38[204]}
   );
   gpc1_1 gpc4488 (
      {stage0_38[440]},
      {stage1_38[205]}
   );
   gpc1_1 gpc4489 (
      {stage0_38[441]},
      {stage1_38[206]}
   );
   gpc1_1 gpc4490 (
      {stage0_38[442]},
      {stage1_38[207]}
   );
   gpc1_1 gpc4491 (
      {stage0_38[443]},
      {stage1_38[208]}
   );
   gpc1_1 gpc4492 (
      {stage0_38[444]},
      {stage1_38[209]}
   );
   gpc1_1 gpc4493 (
      {stage0_38[445]},
      {stage1_38[210]}
   );
   gpc1_1 gpc4494 (
      {stage0_38[446]},
      {stage1_38[211]}
   );
   gpc1_1 gpc4495 (
      {stage0_38[447]},
      {stage1_38[212]}
   );
   gpc1_1 gpc4496 (
      {stage0_38[448]},
      {stage1_38[213]}
   );
   gpc1_1 gpc4497 (
      {stage0_38[449]},
      {stage1_38[214]}
   );
   gpc1_1 gpc4498 (
      {stage0_38[450]},
      {stage1_38[215]}
   );
   gpc1_1 gpc4499 (
      {stage0_38[451]},
      {stage1_38[216]}
   );
   gpc1_1 gpc4500 (
      {stage0_38[452]},
      {stage1_38[217]}
   );
   gpc1_1 gpc4501 (
      {stage0_38[453]},
      {stage1_38[218]}
   );
   gpc1_1 gpc4502 (
      {stage0_38[454]},
      {stage1_38[219]}
   );
   gpc1_1 gpc4503 (
      {stage0_38[455]},
      {stage1_38[220]}
   );
   gpc1_1 gpc4504 (
      {stage0_38[456]},
      {stage1_38[221]}
   );
   gpc1_1 gpc4505 (
      {stage0_38[457]},
      {stage1_38[222]}
   );
   gpc1_1 gpc4506 (
      {stage0_38[458]},
      {stage1_38[223]}
   );
   gpc1_1 gpc4507 (
      {stage0_38[459]},
      {stage1_38[224]}
   );
   gpc1_1 gpc4508 (
      {stage0_38[460]},
      {stage1_38[225]}
   );
   gpc1_1 gpc4509 (
      {stage0_38[461]},
      {stage1_38[226]}
   );
   gpc1_1 gpc4510 (
      {stage0_38[462]},
      {stage1_38[227]}
   );
   gpc1_1 gpc4511 (
      {stage0_38[463]},
      {stage1_38[228]}
   );
   gpc1_1 gpc4512 (
      {stage0_38[464]},
      {stage1_38[229]}
   );
   gpc1_1 gpc4513 (
      {stage0_38[465]},
      {stage1_38[230]}
   );
   gpc1_1 gpc4514 (
      {stage0_38[466]},
      {stage1_38[231]}
   );
   gpc1_1 gpc4515 (
      {stage0_38[467]},
      {stage1_38[232]}
   );
   gpc1_1 gpc4516 (
      {stage0_38[468]},
      {stage1_38[233]}
   );
   gpc1_1 gpc4517 (
      {stage0_38[469]},
      {stage1_38[234]}
   );
   gpc1_1 gpc4518 (
      {stage0_38[470]},
      {stage1_38[235]}
   );
   gpc1_1 gpc4519 (
      {stage0_38[471]},
      {stage1_38[236]}
   );
   gpc1_1 gpc4520 (
      {stage0_38[472]},
      {stage1_38[237]}
   );
   gpc1_1 gpc4521 (
      {stage0_38[473]},
      {stage1_38[238]}
   );
   gpc1_1 gpc4522 (
      {stage0_38[474]},
      {stage1_38[239]}
   );
   gpc1_1 gpc4523 (
      {stage0_38[475]},
      {stage1_38[240]}
   );
   gpc1_1 gpc4524 (
      {stage0_38[476]},
      {stage1_38[241]}
   );
   gpc1_1 gpc4525 (
      {stage0_38[477]},
      {stage1_38[242]}
   );
   gpc1_1 gpc4526 (
      {stage0_38[478]},
      {stage1_38[243]}
   );
   gpc1_1 gpc4527 (
      {stage0_38[479]},
      {stage1_38[244]}
   );
   gpc1_1 gpc4528 (
      {stage0_38[480]},
      {stage1_38[245]}
   );
   gpc1_1 gpc4529 (
      {stage0_38[481]},
      {stage1_38[246]}
   );
   gpc1_1 gpc4530 (
      {stage0_38[482]},
      {stage1_38[247]}
   );
   gpc1_1 gpc4531 (
      {stage0_38[483]},
      {stage1_38[248]}
   );
   gpc1_1 gpc4532 (
      {stage0_38[484]},
      {stage1_38[249]}
   );
   gpc1_1 gpc4533 (
      {stage0_38[485]},
      {stage1_38[250]}
   );
   gpc1_1 gpc4534 (
      {stage0_38[486]},
      {stage1_38[251]}
   );
   gpc1_1 gpc4535 (
      {stage0_38[487]},
      {stage1_38[252]}
   );
   gpc1_1 gpc4536 (
      {stage0_38[488]},
      {stage1_38[253]}
   );
   gpc1_1 gpc4537 (
      {stage0_38[489]},
      {stage1_38[254]}
   );
   gpc1_1 gpc4538 (
      {stage0_38[490]},
      {stage1_38[255]}
   );
   gpc1_1 gpc4539 (
      {stage0_38[491]},
      {stage1_38[256]}
   );
   gpc1_1 gpc4540 (
      {stage0_38[492]},
      {stage1_38[257]}
   );
   gpc1_1 gpc4541 (
      {stage0_38[493]},
      {stage1_38[258]}
   );
   gpc1_1 gpc4542 (
      {stage0_38[494]},
      {stage1_38[259]}
   );
   gpc1_1 gpc4543 (
      {stage0_38[495]},
      {stage1_38[260]}
   );
   gpc1_1 gpc4544 (
      {stage0_38[496]},
      {stage1_38[261]}
   );
   gpc1_1 gpc4545 (
      {stage0_38[497]},
      {stage1_38[262]}
   );
   gpc1_1 gpc4546 (
      {stage0_38[498]},
      {stage1_38[263]}
   );
   gpc1_1 gpc4547 (
      {stage0_38[499]},
      {stage1_38[264]}
   );
   gpc1_1 gpc4548 (
      {stage0_38[500]},
      {stage1_38[265]}
   );
   gpc1_1 gpc4549 (
      {stage0_38[501]},
      {stage1_38[266]}
   );
   gpc1_1 gpc4550 (
      {stage0_38[502]},
      {stage1_38[267]}
   );
   gpc1_1 gpc4551 (
      {stage0_38[503]},
      {stage1_38[268]}
   );
   gpc1_1 gpc4552 (
      {stage0_38[504]},
      {stage1_38[269]}
   );
   gpc1_1 gpc4553 (
      {stage0_38[505]},
      {stage1_38[270]}
   );
   gpc1_1 gpc4554 (
      {stage0_38[506]},
      {stage1_38[271]}
   );
   gpc1_1 gpc4555 (
      {stage0_38[507]},
      {stage1_38[272]}
   );
   gpc1_1 gpc4556 (
      {stage0_38[508]},
      {stage1_38[273]}
   );
   gpc1_1 gpc4557 (
      {stage0_38[509]},
      {stage1_38[274]}
   );
   gpc1_1 gpc4558 (
      {stage0_38[510]},
      {stage1_38[275]}
   );
   gpc1_1 gpc4559 (
      {stage0_38[511]},
      {stage1_38[276]}
   );
   gpc1_1 gpc4560 (
      {stage0_39[491]},
      {stage1_39[176]}
   );
   gpc1_1 gpc4561 (
      {stage0_39[492]},
      {stage1_39[177]}
   );
   gpc1_1 gpc4562 (
      {stage0_39[493]},
      {stage1_39[178]}
   );
   gpc1_1 gpc4563 (
      {stage0_39[494]},
      {stage1_39[179]}
   );
   gpc1_1 gpc4564 (
      {stage0_39[495]},
      {stage1_39[180]}
   );
   gpc1_1 gpc4565 (
      {stage0_39[496]},
      {stage1_39[181]}
   );
   gpc1_1 gpc4566 (
      {stage0_39[497]},
      {stage1_39[182]}
   );
   gpc1_1 gpc4567 (
      {stage0_39[498]},
      {stage1_39[183]}
   );
   gpc1_1 gpc4568 (
      {stage0_39[499]},
      {stage1_39[184]}
   );
   gpc1_1 gpc4569 (
      {stage0_39[500]},
      {stage1_39[185]}
   );
   gpc1_1 gpc4570 (
      {stage0_39[501]},
      {stage1_39[186]}
   );
   gpc1_1 gpc4571 (
      {stage0_39[502]},
      {stage1_39[187]}
   );
   gpc1_1 gpc4572 (
      {stage0_39[503]},
      {stage1_39[188]}
   );
   gpc1_1 gpc4573 (
      {stage0_39[504]},
      {stage1_39[189]}
   );
   gpc1_1 gpc4574 (
      {stage0_39[505]},
      {stage1_39[190]}
   );
   gpc1_1 gpc4575 (
      {stage0_39[506]},
      {stage1_39[191]}
   );
   gpc1_1 gpc4576 (
      {stage0_39[507]},
      {stage1_39[192]}
   );
   gpc1_1 gpc4577 (
      {stage0_39[508]},
      {stage1_39[193]}
   );
   gpc1_1 gpc4578 (
      {stage0_39[509]},
      {stage1_39[194]}
   );
   gpc1_1 gpc4579 (
      {stage0_39[510]},
      {stage1_39[195]}
   );
   gpc1_1 gpc4580 (
      {stage0_39[511]},
      {stage1_39[196]}
   );
   gpc1_1 gpc4581 (
      {stage0_40[489]},
      {stage1_40[207]}
   );
   gpc1_1 gpc4582 (
      {stage0_40[490]},
      {stage1_40[208]}
   );
   gpc1_1 gpc4583 (
      {stage0_40[491]},
      {stage1_40[209]}
   );
   gpc1_1 gpc4584 (
      {stage0_40[492]},
      {stage1_40[210]}
   );
   gpc1_1 gpc4585 (
      {stage0_40[493]},
      {stage1_40[211]}
   );
   gpc1_1 gpc4586 (
      {stage0_40[494]},
      {stage1_40[212]}
   );
   gpc1_1 gpc4587 (
      {stage0_40[495]},
      {stage1_40[213]}
   );
   gpc1_1 gpc4588 (
      {stage0_40[496]},
      {stage1_40[214]}
   );
   gpc1_1 gpc4589 (
      {stage0_40[497]},
      {stage1_40[215]}
   );
   gpc1_1 gpc4590 (
      {stage0_40[498]},
      {stage1_40[216]}
   );
   gpc1_1 gpc4591 (
      {stage0_40[499]},
      {stage1_40[217]}
   );
   gpc1_1 gpc4592 (
      {stage0_40[500]},
      {stage1_40[218]}
   );
   gpc1_1 gpc4593 (
      {stage0_40[501]},
      {stage1_40[219]}
   );
   gpc1_1 gpc4594 (
      {stage0_40[502]},
      {stage1_40[220]}
   );
   gpc1_1 gpc4595 (
      {stage0_40[503]},
      {stage1_40[221]}
   );
   gpc1_1 gpc4596 (
      {stage0_40[504]},
      {stage1_40[222]}
   );
   gpc1_1 gpc4597 (
      {stage0_40[505]},
      {stage1_40[223]}
   );
   gpc1_1 gpc4598 (
      {stage0_40[506]},
      {stage1_40[224]}
   );
   gpc1_1 gpc4599 (
      {stage0_40[507]},
      {stage1_40[225]}
   );
   gpc1_1 gpc4600 (
      {stage0_40[508]},
      {stage1_40[226]}
   );
   gpc1_1 gpc4601 (
      {stage0_40[509]},
      {stage1_40[227]}
   );
   gpc1_1 gpc4602 (
      {stage0_40[510]},
      {stage1_40[228]}
   );
   gpc1_1 gpc4603 (
      {stage0_40[511]},
      {stage1_40[229]}
   );
   gpc1_1 gpc4604 (
      {stage0_41[420]},
      {stage1_41[185]}
   );
   gpc1_1 gpc4605 (
      {stage0_41[421]},
      {stage1_41[186]}
   );
   gpc1_1 gpc4606 (
      {stage0_41[422]},
      {stage1_41[187]}
   );
   gpc1_1 gpc4607 (
      {stage0_41[423]},
      {stage1_41[188]}
   );
   gpc1_1 gpc4608 (
      {stage0_41[424]},
      {stage1_41[189]}
   );
   gpc1_1 gpc4609 (
      {stage0_41[425]},
      {stage1_41[190]}
   );
   gpc1_1 gpc4610 (
      {stage0_41[426]},
      {stage1_41[191]}
   );
   gpc1_1 gpc4611 (
      {stage0_41[427]},
      {stage1_41[192]}
   );
   gpc1_1 gpc4612 (
      {stage0_41[428]},
      {stage1_41[193]}
   );
   gpc1_1 gpc4613 (
      {stage0_41[429]},
      {stage1_41[194]}
   );
   gpc1_1 gpc4614 (
      {stage0_41[430]},
      {stage1_41[195]}
   );
   gpc1_1 gpc4615 (
      {stage0_41[431]},
      {stage1_41[196]}
   );
   gpc1_1 gpc4616 (
      {stage0_41[432]},
      {stage1_41[197]}
   );
   gpc1_1 gpc4617 (
      {stage0_41[433]},
      {stage1_41[198]}
   );
   gpc1_1 gpc4618 (
      {stage0_41[434]},
      {stage1_41[199]}
   );
   gpc1_1 gpc4619 (
      {stage0_41[435]},
      {stage1_41[200]}
   );
   gpc1_1 gpc4620 (
      {stage0_41[436]},
      {stage1_41[201]}
   );
   gpc1_1 gpc4621 (
      {stage0_41[437]},
      {stage1_41[202]}
   );
   gpc1_1 gpc4622 (
      {stage0_41[438]},
      {stage1_41[203]}
   );
   gpc1_1 gpc4623 (
      {stage0_41[439]},
      {stage1_41[204]}
   );
   gpc1_1 gpc4624 (
      {stage0_41[440]},
      {stage1_41[205]}
   );
   gpc1_1 gpc4625 (
      {stage0_41[441]},
      {stage1_41[206]}
   );
   gpc1_1 gpc4626 (
      {stage0_41[442]},
      {stage1_41[207]}
   );
   gpc1_1 gpc4627 (
      {stage0_41[443]},
      {stage1_41[208]}
   );
   gpc1_1 gpc4628 (
      {stage0_41[444]},
      {stage1_41[209]}
   );
   gpc1_1 gpc4629 (
      {stage0_41[445]},
      {stage1_41[210]}
   );
   gpc1_1 gpc4630 (
      {stage0_41[446]},
      {stage1_41[211]}
   );
   gpc1_1 gpc4631 (
      {stage0_41[447]},
      {stage1_41[212]}
   );
   gpc1_1 gpc4632 (
      {stage0_41[448]},
      {stage1_41[213]}
   );
   gpc1_1 gpc4633 (
      {stage0_41[449]},
      {stage1_41[214]}
   );
   gpc1_1 gpc4634 (
      {stage0_41[450]},
      {stage1_41[215]}
   );
   gpc1_1 gpc4635 (
      {stage0_41[451]},
      {stage1_41[216]}
   );
   gpc1_1 gpc4636 (
      {stage0_41[452]},
      {stage1_41[217]}
   );
   gpc1_1 gpc4637 (
      {stage0_41[453]},
      {stage1_41[218]}
   );
   gpc1_1 gpc4638 (
      {stage0_41[454]},
      {stage1_41[219]}
   );
   gpc1_1 gpc4639 (
      {stage0_41[455]},
      {stage1_41[220]}
   );
   gpc1_1 gpc4640 (
      {stage0_41[456]},
      {stage1_41[221]}
   );
   gpc1_1 gpc4641 (
      {stage0_41[457]},
      {stage1_41[222]}
   );
   gpc1_1 gpc4642 (
      {stage0_41[458]},
      {stage1_41[223]}
   );
   gpc1_1 gpc4643 (
      {stage0_41[459]},
      {stage1_41[224]}
   );
   gpc1_1 gpc4644 (
      {stage0_41[460]},
      {stage1_41[225]}
   );
   gpc1_1 gpc4645 (
      {stage0_41[461]},
      {stage1_41[226]}
   );
   gpc1_1 gpc4646 (
      {stage0_41[462]},
      {stage1_41[227]}
   );
   gpc1_1 gpc4647 (
      {stage0_41[463]},
      {stage1_41[228]}
   );
   gpc1_1 gpc4648 (
      {stage0_41[464]},
      {stage1_41[229]}
   );
   gpc1_1 gpc4649 (
      {stage0_41[465]},
      {stage1_41[230]}
   );
   gpc1_1 gpc4650 (
      {stage0_41[466]},
      {stage1_41[231]}
   );
   gpc1_1 gpc4651 (
      {stage0_41[467]},
      {stage1_41[232]}
   );
   gpc1_1 gpc4652 (
      {stage0_41[468]},
      {stage1_41[233]}
   );
   gpc1_1 gpc4653 (
      {stage0_41[469]},
      {stage1_41[234]}
   );
   gpc1_1 gpc4654 (
      {stage0_41[470]},
      {stage1_41[235]}
   );
   gpc1_1 gpc4655 (
      {stage0_41[471]},
      {stage1_41[236]}
   );
   gpc1_1 gpc4656 (
      {stage0_41[472]},
      {stage1_41[237]}
   );
   gpc1_1 gpc4657 (
      {stage0_41[473]},
      {stage1_41[238]}
   );
   gpc1_1 gpc4658 (
      {stage0_41[474]},
      {stage1_41[239]}
   );
   gpc1_1 gpc4659 (
      {stage0_41[475]},
      {stage1_41[240]}
   );
   gpc1_1 gpc4660 (
      {stage0_41[476]},
      {stage1_41[241]}
   );
   gpc1_1 gpc4661 (
      {stage0_41[477]},
      {stage1_41[242]}
   );
   gpc1_1 gpc4662 (
      {stage0_41[478]},
      {stage1_41[243]}
   );
   gpc1_1 gpc4663 (
      {stage0_41[479]},
      {stage1_41[244]}
   );
   gpc1_1 gpc4664 (
      {stage0_41[480]},
      {stage1_41[245]}
   );
   gpc1_1 gpc4665 (
      {stage0_41[481]},
      {stage1_41[246]}
   );
   gpc1_1 gpc4666 (
      {stage0_41[482]},
      {stage1_41[247]}
   );
   gpc1_1 gpc4667 (
      {stage0_41[483]},
      {stage1_41[248]}
   );
   gpc1_1 gpc4668 (
      {stage0_41[484]},
      {stage1_41[249]}
   );
   gpc1_1 gpc4669 (
      {stage0_41[485]},
      {stage1_41[250]}
   );
   gpc1_1 gpc4670 (
      {stage0_41[486]},
      {stage1_41[251]}
   );
   gpc1_1 gpc4671 (
      {stage0_41[487]},
      {stage1_41[252]}
   );
   gpc1_1 gpc4672 (
      {stage0_41[488]},
      {stage1_41[253]}
   );
   gpc1_1 gpc4673 (
      {stage0_41[489]},
      {stage1_41[254]}
   );
   gpc1_1 gpc4674 (
      {stage0_41[490]},
      {stage1_41[255]}
   );
   gpc1_1 gpc4675 (
      {stage0_41[491]},
      {stage1_41[256]}
   );
   gpc1_1 gpc4676 (
      {stage0_41[492]},
      {stage1_41[257]}
   );
   gpc1_1 gpc4677 (
      {stage0_41[493]},
      {stage1_41[258]}
   );
   gpc1_1 gpc4678 (
      {stage0_41[494]},
      {stage1_41[259]}
   );
   gpc1_1 gpc4679 (
      {stage0_41[495]},
      {stage1_41[260]}
   );
   gpc1_1 gpc4680 (
      {stage0_41[496]},
      {stage1_41[261]}
   );
   gpc1_1 gpc4681 (
      {stage0_41[497]},
      {stage1_41[262]}
   );
   gpc1_1 gpc4682 (
      {stage0_41[498]},
      {stage1_41[263]}
   );
   gpc1_1 gpc4683 (
      {stage0_41[499]},
      {stage1_41[264]}
   );
   gpc1_1 gpc4684 (
      {stage0_41[500]},
      {stage1_41[265]}
   );
   gpc1_1 gpc4685 (
      {stage0_41[501]},
      {stage1_41[266]}
   );
   gpc1_1 gpc4686 (
      {stage0_41[502]},
      {stage1_41[267]}
   );
   gpc1_1 gpc4687 (
      {stage0_41[503]},
      {stage1_41[268]}
   );
   gpc1_1 gpc4688 (
      {stage0_41[504]},
      {stage1_41[269]}
   );
   gpc1_1 gpc4689 (
      {stage0_41[505]},
      {stage1_41[270]}
   );
   gpc1_1 gpc4690 (
      {stage0_41[506]},
      {stage1_41[271]}
   );
   gpc1_1 gpc4691 (
      {stage0_41[507]},
      {stage1_41[272]}
   );
   gpc1_1 gpc4692 (
      {stage0_41[508]},
      {stage1_41[273]}
   );
   gpc1_1 gpc4693 (
      {stage0_41[509]},
      {stage1_41[274]}
   );
   gpc1_1 gpc4694 (
      {stage0_41[510]},
      {stage1_41[275]}
   );
   gpc1_1 gpc4695 (
      {stage0_41[511]},
      {stage1_41[276]}
   );
   gpc1_1 gpc4696 (
      {stage0_42[451]},
      {stage1_42[168]}
   );
   gpc1_1 gpc4697 (
      {stage0_42[452]},
      {stage1_42[169]}
   );
   gpc1_1 gpc4698 (
      {stage0_42[453]},
      {stage1_42[170]}
   );
   gpc1_1 gpc4699 (
      {stage0_42[454]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4700 (
      {stage0_42[455]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4701 (
      {stage0_42[456]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4702 (
      {stage0_42[457]},
      {stage1_42[174]}
   );
   gpc1_1 gpc4703 (
      {stage0_42[458]},
      {stage1_42[175]}
   );
   gpc1_1 gpc4704 (
      {stage0_42[459]},
      {stage1_42[176]}
   );
   gpc1_1 gpc4705 (
      {stage0_42[460]},
      {stage1_42[177]}
   );
   gpc1_1 gpc4706 (
      {stage0_42[461]},
      {stage1_42[178]}
   );
   gpc1_1 gpc4707 (
      {stage0_42[462]},
      {stage1_42[179]}
   );
   gpc1_1 gpc4708 (
      {stage0_42[463]},
      {stage1_42[180]}
   );
   gpc1_1 gpc4709 (
      {stage0_42[464]},
      {stage1_42[181]}
   );
   gpc1_1 gpc4710 (
      {stage0_42[465]},
      {stage1_42[182]}
   );
   gpc1_1 gpc4711 (
      {stage0_42[466]},
      {stage1_42[183]}
   );
   gpc1_1 gpc4712 (
      {stage0_42[467]},
      {stage1_42[184]}
   );
   gpc1_1 gpc4713 (
      {stage0_42[468]},
      {stage1_42[185]}
   );
   gpc1_1 gpc4714 (
      {stage0_42[469]},
      {stage1_42[186]}
   );
   gpc1_1 gpc4715 (
      {stage0_42[470]},
      {stage1_42[187]}
   );
   gpc1_1 gpc4716 (
      {stage0_42[471]},
      {stage1_42[188]}
   );
   gpc1_1 gpc4717 (
      {stage0_42[472]},
      {stage1_42[189]}
   );
   gpc1_1 gpc4718 (
      {stage0_42[473]},
      {stage1_42[190]}
   );
   gpc1_1 gpc4719 (
      {stage0_42[474]},
      {stage1_42[191]}
   );
   gpc1_1 gpc4720 (
      {stage0_42[475]},
      {stage1_42[192]}
   );
   gpc1_1 gpc4721 (
      {stage0_42[476]},
      {stage1_42[193]}
   );
   gpc1_1 gpc4722 (
      {stage0_42[477]},
      {stage1_42[194]}
   );
   gpc1_1 gpc4723 (
      {stage0_42[478]},
      {stage1_42[195]}
   );
   gpc1_1 gpc4724 (
      {stage0_42[479]},
      {stage1_42[196]}
   );
   gpc1_1 gpc4725 (
      {stage0_42[480]},
      {stage1_42[197]}
   );
   gpc1_1 gpc4726 (
      {stage0_42[481]},
      {stage1_42[198]}
   );
   gpc1_1 gpc4727 (
      {stage0_42[482]},
      {stage1_42[199]}
   );
   gpc1_1 gpc4728 (
      {stage0_42[483]},
      {stage1_42[200]}
   );
   gpc1_1 gpc4729 (
      {stage0_42[484]},
      {stage1_42[201]}
   );
   gpc1_1 gpc4730 (
      {stage0_42[485]},
      {stage1_42[202]}
   );
   gpc1_1 gpc4731 (
      {stage0_42[486]},
      {stage1_42[203]}
   );
   gpc1_1 gpc4732 (
      {stage0_42[487]},
      {stage1_42[204]}
   );
   gpc1_1 gpc4733 (
      {stage0_42[488]},
      {stage1_42[205]}
   );
   gpc1_1 gpc4734 (
      {stage0_42[489]},
      {stage1_42[206]}
   );
   gpc1_1 gpc4735 (
      {stage0_42[490]},
      {stage1_42[207]}
   );
   gpc1_1 gpc4736 (
      {stage0_42[491]},
      {stage1_42[208]}
   );
   gpc1_1 gpc4737 (
      {stage0_42[492]},
      {stage1_42[209]}
   );
   gpc1_1 gpc4738 (
      {stage0_42[493]},
      {stage1_42[210]}
   );
   gpc1_1 gpc4739 (
      {stage0_42[494]},
      {stage1_42[211]}
   );
   gpc1_1 gpc4740 (
      {stage0_42[495]},
      {stage1_42[212]}
   );
   gpc1_1 gpc4741 (
      {stage0_42[496]},
      {stage1_42[213]}
   );
   gpc1_1 gpc4742 (
      {stage0_42[497]},
      {stage1_42[214]}
   );
   gpc1_1 gpc4743 (
      {stage0_42[498]},
      {stage1_42[215]}
   );
   gpc1_1 gpc4744 (
      {stage0_42[499]},
      {stage1_42[216]}
   );
   gpc1_1 gpc4745 (
      {stage0_42[500]},
      {stage1_42[217]}
   );
   gpc1_1 gpc4746 (
      {stage0_42[501]},
      {stage1_42[218]}
   );
   gpc1_1 gpc4747 (
      {stage0_42[502]},
      {stage1_42[219]}
   );
   gpc1_1 gpc4748 (
      {stage0_42[503]},
      {stage1_42[220]}
   );
   gpc1_1 gpc4749 (
      {stage0_42[504]},
      {stage1_42[221]}
   );
   gpc1_1 gpc4750 (
      {stage0_42[505]},
      {stage1_42[222]}
   );
   gpc1_1 gpc4751 (
      {stage0_42[506]},
      {stage1_42[223]}
   );
   gpc1_1 gpc4752 (
      {stage0_42[507]},
      {stage1_42[224]}
   );
   gpc1_1 gpc4753 (
      {stage0_42[508]},
      {stage1_42[225]}
   );
   gpc1_1 gpc4754 (
      {stage0_42[509]},
      {stage1_42[226]}
   );
   gpc1_1 gpc4755 (
      {stage0_42[510]},
      {stage1_42[227]}
   );
   gpc1_1 gpc4756 (
      {stage0_42[511]},
      {stage1_42[228]}
   );
   gpc1_1 gpc4757 (
      {stage0_43[475]},
      {stage1_43[207]}
   );
   gpc1_1 gpc4758 (
      {stage0_43[476]},
      {stage1_43[208]}
   );
   gpc1_1 gpc4759 (
      {stage0_43[477]},
      {stage1_43[209]}
   );
   gpc1_1 gpc4760 (
      {stage0_43[478]},
      {stage1_43[210]}
   );
   gpc1_1 gpc4761 (
      {stage0_43[479]},
      {stage1_43[211]}
   );
   gpc1_1 gpc4762 (
      {stage0_43[480]},
      {stage1_43[212]}
   );
   gpc1_1 gpc4763 (
      {stage0_43[481]},
      {stage1_43[213]}
   );
   gpc1_1 gpc4764 (
      {stage0_43[482]},
      {stage1_43[214]}
   );
   gpc1_1 gpc4765 (
      {stage0_43[483]},
      {stage1_43[215]}
   );
   gpc1_1 gpc4766 (
      {stage0_43[484]},
      {stage1_43[216]}
   );
   gpc1_1 gpc4767 (
      {stage0_43[485]},
      {stage1_43[217]}
   );
   gpc1_1 gpc4768 (
      {stage0_43[486]},
      {stage1_43[218]}
   );
   gpc1_1 gpc4769 (
      {stage0_43[487]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4770 (
      {stage0_43[488]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4771 (
      {stage0_43[489]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4772 (
      {stage0_43[490]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4773 (
      {stage0_43[491]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4774 (
      {stage0_43[492]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4775 (
      {stage0_43[493]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4776 (
      {stage0_43[494]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4777 (
      {stage0_43[495]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4778 (
      {stage0_43[496]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4779 (
      {stage0_43[497]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4780 (
      {stage0_43[498]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4781 (
      {stage0_43[499]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4782 (
      {stage0_43[500]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4783 (
      {stage0_43[501]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4784 (
      {stage0_43[502]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4785 (
      {stage0_43[503]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4786 (
      {stage0_43[504]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4787 (
      {stage0_43[505]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4788 (
      {stage0_43[506]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4789 (
      {stage0_43[507]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4790 (
      {stage0_43[508]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4791 (
      {stage0_43[509]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4792 (
      {stage0_43[510]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4793 (
      {stage0_43[511]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4794 (
      {stage0_44[448]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4795 (
      {stage0_44[449]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4796 (
      {stage0_44[450]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4797 (
      {stage0_44[451]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4798 (
      {stage0_44[452]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4799 (
      {stage0_44[453]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4800 (
      {stage0_44[454]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4801 (
      {stage0_44[455]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4802 (
      {stage0_44[456]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4803 (
      {stage0_44[457]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4804 (
      {stage0_44[458]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4805 (
      {stage0_44[459]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4806 (
      {stage0_44[460]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4807 (
      {stage0_44[461]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4808 (
      {stage0_44[462]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4809 (
      {stage0_44[463]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4810 (
      {stage0_44[464]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4811 (
      {stage0_44[465]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4812 (
      {stage0_44[466]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4813 (
      {stage0_44[467]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4814 (
      {stage0_44[468]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4815 (
      {stage0_44[469]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4816 (
      {stage0_44[470]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4817 (
      {stage0_44[471]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4818 (
      {stage0_44[472]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4819 (
      {stage0_44[473]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4820 (
      {stage0_44[474]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4821 (
      {stage0_44[475]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4822 (
      {stage0_44[476]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4823 (
      {stage0_44[477]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4824 (
      {stage0_44[478]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4825 (
      {stage0_44[479]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4826 (
      {stage0_44[480]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4827 (
      {stage0_44[481]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4828 (
      {stage0_44[482]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4829 (
      {stage0_44[483]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4830 (
      {stage0_44[484]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4831 (
      {stage0_44[485]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4832 (
      {stage0_44[486]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4833 (
      {stage0_44[487]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4834 (
      {stage0_44[488]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4835 (
      {stage0_44[489]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4836 (
      {stage0_44[490]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4837 (
      {stage0_44[491]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4838 (
      {stage0_44[492]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4839 (
      {stage0_44[493]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4840 (
      {stage0_44[494]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4841 (
      {stage0_44[495]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4842 (
      {stage0_44[496]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4843 (
      {stage0_44[497]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4844 (
      {stage0_44[498]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4845 (
      {stage0_44[499]},
      {stage1_44[256]}
   );
   gpc1_1 gpc4846 (
      {stage0_44[500]},
      {stage1_44[257]}
   );
   gpc1_1 gpc4847 (
      {stage0_44[501]},
      {stage1_44[258]}
   );
   gpc1_1 gpc4848 (
      {stage0_44[502]},
      {stage1_44[259]}
   );
   gpc1_1 gpc4849 (
      {stage0_44[503]},
      {stage1_44[260]}
   );
   gpc1_1 gpc4850 (
      {stage0_44[504]},
      {stage1_44[261]}
   );
   gpc1_1 gpc4851 (
      {stage0_44[505]},
      {stage1_44[262]}
   );
   gpc1_1 gpc4852 (
      {stage0_44[506]},
      {stage1_44[263]}
   );
   gpc1_1 gpc4853 (
      {stage0_44[507]},
      {stage1_44[264]}
   );
   gpc1_1 gpc4854 (
      {stage0_44[508]},
      {stage1_44[265]}
   );
   gpc1_1 gpc4855 (
      {stage0_44[509]},
      {stage1_44[266]}
   );
   gpc1_1 gpc4856 (
      {stage0_44[510]},
      {stage1_44[267]}
   );
   gpc1_1 gpc4857 (
      {stage0_44[511]},
      {stage1_44[268]}
   );
   gpc1_1 gpc4858 (
      {stage0_45[498]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4859 (
      {stage0_45[499]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4860 (
      {stage0_45[500]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4861 (
      {stage0_45[501]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4862 (
      {stage0_45[502]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4863 (
      {stage0_45[503]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4864 (
      {stage0_45[504]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4865 (
      {stage0_45[505]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4866 (
      {stage0_45[506]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4867 (
      {stage0_45[507]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4868 (
      {stage0_45[508]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4869 (
      {stage0_45[509]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4870 (
      {stage0_45[510]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4871 (
      {stage0_45[511]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4872 (
      {stage0_46[388]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4873 (
      {stage0_46[389]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4874 (
      {stage0_46[390]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4875 (
      {stage0_46[391]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4876 (
      {stage0_46[392]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4877 (
      {stage0_46[393]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4878 (
      {stage0_46[394]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4879 (
      {stage0_46[395]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4880 (
      {stage0_46[396]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4881 (
      {stage0_46[397]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4882 (
      {stage0_46[398]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4883 (
      {stage0_46[399]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4884 (
      {stage0_46[400]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4885 (
      {stage0_46[401]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4886 (
      {stage0_46[402]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4887 (
      {stage0_46[403]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4888 (
      {stage0_46[404]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4889 (
      {stage0_46[405]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4890 (
      {stage0_46[406]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4891 (
      {stage0_46[407]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4892 (
      {stage0_46[408]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4893 (
      {stage0_46[409]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4894 (
      {stage0_46[410]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4895 (
      {stage0_46[411]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4896 (
      {stage0_46[412]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4897 (
      {stage0_46[413]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4898 (
      {stage0_46[414]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4899 (
      {stage0_46[415]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4900 (
      {stage0_46[416]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4901 (
      {stage0_46[417]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4902 (
      {stage0_46[418]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4903 (
      {stage0_46[419]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4904 (
      {stage0_46[420]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4905 (
      {stage0_46[421]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4906 (
      {stage0_46[422]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4907 (
      {stage0_46[423]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4908 (
      {stage0_46[424]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4909 (
      {stage0_46[425]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4910 (
      {stage0_46[426]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4911 (
      {stage0_46[427]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4912 (
      {stage0_46[428]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4913 (
      {stage0_46[429]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4914 (
      {stage0_46[430]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4915 (
      {stage0_46[431]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4916 (
      {stage0_46[432]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4917 (
      {stage0_46[433]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4918 (
      {stage0_46[434]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4919 (
      {stage0_46[435]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4920 (
      {stage0_46[436]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4921 (
      {stage0_46[437]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4922 (
      {stage0_46[438]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4923 (
      {stage0_46[439]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4924 (
      {stage0_46[440]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4925 (
      {stage0_46[441]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4926 (
      {stage0_46[442]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4927 (
      {stage0_46[443]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4928 (
      {stage0_46[444]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4929 (
      {stage0_46[445]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4930 (
      {stage0_46[446]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4931 (
      {stage0_46[447]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4932 (
      {stage0_46[448]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4933 (
      {stage0_46[449]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4934 (
      {stage0_46[450]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4935 (
      {stage0_46[451]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4936 (
      {stage0_46[452]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4937 (
      {stage0_46[453]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4938 (
      {stage0_46[454]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4939 (
      {stage0_46[455]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4940 (
      {stage0_46[456]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4941 (
      {stage0_46[457]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4942 (
      {stage0_46[458]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4943 (
      {stage0_46[459]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4944 (
      {stage0_46[460]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4945 (
      {stage0_46[461]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4946 (
      {stage0_46[462]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4947 (
      {stage0_46[463]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4948 (
      {stage0_46[464]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4949 (
      {stage0_46[465]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4950 (
      {stage0_46[466]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4951 (
      {stage0_46[467]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4952 (
      {stage0_46[468]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4953 (
      {stage0_46[469]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4954 (
      {stage0_46[470]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4955 (
      {stage0_46[471]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4956 (
      {stage0_46[472]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4957 (
      {stage0_46[473]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4958 (
      {stage0_46[474]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4959 (
      {stage0_46[475]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4960 (
      {stage0_46[476]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4961 (
      {stage0_46[477]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4962 (
      {stage0_46[478]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4963 (
      {stage0_46[479]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4964 (
      {stage0_46[480]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4965 (
      {stage0_46[481]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4966 (
      {stage0_46[482]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4967 (
      {stage0_46[483]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4968 (
      {stage0_46[484]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4969 (
      {stage0_46[485]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4970 (
      {stage0_46[486]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4971 (
      {stage0_46[487]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4972 (
      {stage0_46[488]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4973 (
      {stage0_46[489]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4974 (
      {stage0_46[490]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4975 (
      {stage0_46[491]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4976 (
      {stage0_46[492]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4977 (
      {stage0_46[493]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4978 (
      {stage0_46[494]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4979 (
      {stage0_46[495]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4980 (
      {stage0_46[496]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4981 (
      {stage0_46[497]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4982 (
      {stage0_46[498]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4983 (
      {stage0_46[499]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4984 (
      {stage0_46[500]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4985 (
      {stage0_46[501]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4986 (
      {stage0_46[502]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4987 (
      {stage0_46[503]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4988 (
      {stage0_46[504]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4989 (
      {stage0_46[505]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4990 (
      {stage0_46[506]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4991 (
      {stage0_46[507]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4992 (
      {stage0_46[508]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4993 (
      {stage0_46[509]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4994 (
      {stage0_46[510]},
      {stage1_46[298]}
   );
   gpc1_1 gpc4995 (
      {stage0_46[511]},
      {stage1_46[299]}
   );
   gpc1_1 gpc4996 (
      {stage0_47[437]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4997 (
      {stage0_47[438]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4998 (
      {stage0_47[439]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4999 (
      {stage0_47[440]},
      {stage1_47[206]}
   );
   gpc1_1 gpc5000 (
      {stage0_47[441]},
      {stage1_47[207]}
   );
   gpc1_1 gpc5001 (
      {stage0_47[442]},
      {stage1_47[208]}
   );
   gpc1_1 gpc5002 (
      {stage0_47[443]},
      {stage1_47[209]}
   );
   gpc1_1 gpc5003 (
      {stage0_47[444]},
      {stage1_47[210]}
   );
   gpc1_1 gpc5004 (
      {stage0_47[445]},
      {stage1_47[211]}
   );
   gpc1_1 gpc5005 (
      {stage0_47[446]},
      {stage1_47[212]}
   );
   gpc1_1 gpc5006 (
      {stage0_47[447]},
      {stage1_47[213]}
   );
   gpc1_1 gpc5007 (
      {stage0_47[448]},
      {stage1_47[214]}
   );
   gpc1_1 gpc5008 (
      {stage0_47[449]},
      {stage1_47[215]}
   );
   gpc1_1 gpc5009 (
      {stage0_47[450]},
      {stage1_47[216]}
   );
   gpc1_1 gpc5010 (
      {stage0_47[451]},
      {stage1_47[217]}
   );
   gpc1_1 gpc5011 (
      {stage0_47[452]},
      {stage1_47[218]}
   );
   gpc1_1 gpc5012 (
      {stage0_47[453]},
      {stage1_47[219]}
   );
   gpc1_1 gpc5013 (
      {stage0_47[454]},
      {stage1_47[220]}
   );
   gpc1_1 gpc5014 (
      {stage0_47[455]},
      {stage1_47[221]}
   );
   gpc1_1 gpc5015 (
      {stage0_47[456]},
      {stage1_47[222]}
   );
   gpc1_1 gpc5016 (
      {stage0_47[457]},
      {stage1_47[223]}
   );
   gpc1_1 gpc5017 (
      {stage0_47[458]},
      {stage1_47[224]}
   );
   gpc1_1 gpc5018 (
      {stage0_47[459]},
      {stage1_47[225]}
   );
   gpc1_1 gpc5019 (
      {stage0_47[460]},
      {stage1_47[226]}
   );
   gpc1_1 gpc5020 (
      {stage0_47[461]},
      {stage1_47[227]}
   );
   gpc1_1 gpc5021 (
      {stage0_47[462]},
      {stage1_47[228]}
   );
   gpc1_1 gpc5022 (
      {stage0_47[463]},
      {stage1_47[229]}
   );
   gpc1_1 gpc5023 (
      {stage0_47[464]},
      {stage1_47[230]}
   );
   gpc1_1 gpc5024 (
      {stage0_47[465]},
      {stage1_47[231]}
   );
   gpc1_1 gpc5025 (
      {stage0_47[466]},
      {stage1_47[232]}
   );
   gpc1_1 gpc5026 (
      {stage0_47[467]},
      {stage1_47[233]}
   );
   gpc1_1 gpc5027 (
      {stage0_47[468]},
      {stage1_47[234]}
   );
   gpc1_1 gpc5028 (
      {stage0_47[469]},
      {stage1_47[235]}
   );
   gpc1_1 gpc5029 (
      {stage0_47[470]},
      {stage1_47[236]}
   );
   gpc1_1 gpc5030 (
      {stage0_47[471]},
      {stage1_47[237]}
   );
   gpc1_1 gpc5031 (
      {stage0_47[472]},
      {stage1_47[238]}
   );
   gpc1_1 gpc5032 (
      {stage0_47[473]},
      {stage1_47[239]}
   );
   gpc1_1 gpc5033 (
      {stage0_47[474]},
      {stage1_47[240]}
   );
   gpc1_1 gpc5034 (
      {stage0_47[475]},
      {stage1_47[241]}
   );
   gpc1_1 gpc5035 (
      {stage0_47[476]},
      {stage1_47[242]}
   );
   gpc1_1 gpc5036 (
      {stage0_47[477]},
      {stage1_47[243]}
   );
   gpc1_1 gpc5037 (
      {stage0_47[478]},
      {stage1_47[244]}
   );
   gpc1_1 gpc5038 (
      {stage0_47[479]},
      {stage1_47[245]}
   );
   gpc1_1 gpc5039 (
      {stage0_47[480]},
      {stage1_47[246]}
   );
   gpc1_1 gpc5040 (
      {stage0_47[481]},
      {stage1_47[247]}
   );
   gpc1_1 gpc5041 (
      {stage0_47[482]},
      {stage1_47[248]}
   );
   gpc1_1 gpc5042 (
      {stage0_47[483]},
      {stage1_47[249]}
   );
   gpc1_1 gpc5043 (
      {stage0_47[484]},
      {stage1_47[250]}
   );
   gpc1_1 gpc5044 (
      {stage0_47[485]},
      {stage1_47[251]}
   );
   gpc1_1 gpc5045 (
      {stage0_47[486]},
      {stage1_47[252]}
   );
   gpc1_1 gpc5046 (
      {stage0_47[487]},
      {stage1_47[253]}
   );
   gpc1_1 gpc5047 (
      {stage0_47[488]},
      {stage1_47[254]}
   );
   gpc1_1 gpc5048 (
      {stage0_47[489]},
      {stage1_47[255]}
   );
   gpc1_1 gpc5049 (
      {stage0_47[490]},
      {stage1_47[256]}
   );
   gpc1_1 gpc5050 (
      {stage0_47[491]},
      {stage1_47[257]}
   );
   gpc1_1 gpc5051 (
      {stage0_47[492]},
      {stage1_47[258]}
   );
   gpc1_1 gpc5052 (
      {stage0_47[493]},
      {stage1_47[259]}
   );
   gpc1_1 gpc5053 (
      {stage0_47[494]},
      {stage1_47[260]}
   );
   gpc1_1 gpc5054 (
      {stage0_47[495]},
      {stage1_47[261]}
   );
   gpc1_1 gpc5055 (
      {stage0_47[496]},
      {stage1_47[262]}
   );
   gpc1_1 gpc5056 (
      {stage0_47[497]},
      {stage1_47[263]}
   );
   gpc1_1 gpc5057 (
      {stage0_47[498]},
      {stage1_47[264]}
   );
   gpc1_1 gpc5058 (
      {stage0_47[499]},
      {stage1_47[265]}
   );
   gpc1_1 gpc5059 (
      {stage0_47[500]},
      {stage1_47[266]}
   );
   gpc1_1 gpc5060 (
      {stage0_47[501]},
      {stage1_47[267]}
   );
   gpc1_1 gpc5061 (
      {stage0_47[502]},
      {stage1_47[268]}
   );
   gpc1_1 gpc5062 (
      {stage0_47[503]},
      {stage1_47[269]}
   );
   gpc1_1 gpc5063 (
      {stage0_47[504]},
      {stage1_47[270]}
   );
   gpc1_1 gpc5064 (
      {stage0_47[505]},
      {stage1_47[271]}
   );
   gpc1_1 gpc5065 (
      {stage0_47[506]},
      {stage1_47[272]}
   );
   gpc1_1 gpc5066 (
      {stage0_47[507]},
      {stage1_47[273]}
   );
   gpc1_1 gpc5067 (
      {stage0_47[508]},
      {stage1_47[274]}
   );
   gpc1_1 gpc5068 (
      {stage0_47[509]},
      {stage1_47[275]}
   );
   gpc1_1 gpc5069 (
      {stage0_47[510]},
      {stage1_47[276]}
   );
   gpc1_1 gpc5070 (
      {stage0_47[511]},
      {stage1_47[277]}
   );
   gpc1_1 gpc5071 (
      {stage0_48[495]},
      {stage1_48[194]}
   );
   gpc1_1 gpc5072 (
      {stage0_48[496]},
      {stage1_48[195]}
   );
   gpc1_1 gpc5073 (
      {stage0_48[497]},
      {stage1_48[196]}
   );
   gpc1_1 gpc5074 (
      {stage0_48[498]},
      {stage1_48[197]}
   );
   gpc1_1 gpc5075 (
      {stage0_48[499]},
      {stage1_48[198]}
   );
   gpc1_1 gpc5076 (
      {stage0_48[500]},
      {stage1_48[199]}
   );
   gpc1_1 gpc5077 (
      {stage0_48[501]},
      {stage1_48[200]}
   );
   gpc1_1 gpc5078 (
      {stage0_48[502]},
      {stage1_48[201]}
   );
   gpc1_1 gpc5079 (
      {stage0_48[503]},
      {stage1_48[202]}
   );
   gpc1_1 gpc5080 (
      {stage0_48[504]},
      {stage1_48[203]}
   );
   gpc1_1 gpc5081 (
      {stage0_48[505]},
      {stage1_48[204]}
   );
   gpc1_1 gpc5082 (
      {stage0_48[506]},
      {stage1_48[205]}
   );
   gpc1_1 gpc5083 (
      {stage0_48[507]},
      {stage1_48[206]}
   );
   gpc1_1 gpc5084 (
      {stage0_48[508]},
      {stage1_48[207]}
   );
   gpc1_1 gpc5085 (
      {stage0_48[509]},
      {stage1_48[208]}
   );
   gpc1_1 gpc5086 (
      {stage0_48[510]},
      {stage1_48[209]}
   );
   gpc1_1 gpc5087 (
      {stage0_48[511]},
      {stage1_48[210]}
   );
   gpc1_1 gpc5088 (
      {stage0_49[444]},
      {stage1_49[174]}
   );
   gpc1_1 gpc5089 (
      {stage0_49[445]},
      {stage1_49[175]}
   );
   gpc1_1 gpc5090 (
      {stage0_49[446]},
      {stage1_49[176]}
   );
   gpc1_1 gpc5091 (
      {stage0_49[447]},
      {stage1_49[177]}
   );
   gpc1_1 gpc5092 (
      {stage0_49[448]},
      {stage1_49[178]}
   );
   gpc1_1 gpc5093 (
      {stage0_49[449]},
      {stage1_49[179]}
   );
   gpc1_1 gpc5094 (
      {stage0_49[450]},
      {stage1_49[180]}
   );
   gpc1_1 gpc5095 (
      {stage0_49[451]},
      {stage1_49[181]}
   );
   gpc1_1 gpc5096 (
      {stage0_49[452]},
      {stage1_49[182]}
   );
   gpc1_1 gpc5097 (
      {stage0_49[453]},
      {stage1_49[183]}
   );
   gpc1_1 gpc5098 (
      {stage0_49[454]},
      {stage1_49[184]}
   );
   gpc1_1 gpc5099 (
      {stage0_49[455]},
      {stage1_49[185]}
   );
   gpc1_1 gpc5100 (
      {stage0_49[456]},
      {stage1_49[186]}
   );
   gpc1_1 gpc5101 (
      {stage0_49[457]},
      {stage1_49[187]}
   );
   gpc1_1 gpc5102 (
      {stage0_49[458]},
      {stage1_49[188]}
   );
   gpc1_1 gpc5103 (
      {stage0_49[459]},
      {stage1_49[189]}
   );
   gpc1_1 gpc5104 (
      {stage0_49[460]},
      {stage1_49[190]}
   );
   gpc1_1 gpc5105 (
      {stage0_49[461]},
      {stage1_49[191]}
   );
   gpc1_1 gpc5106 (
      {stage0_49[462]},
      {stage1_49[192]}
   );
   gpc1_1 gpc5107 (
      {stage0_49[463]},
      {stage1_49[193]}
   );
   gpc1_1 gpc5108 (
      {stage0_49[464]},
      {stage1_49[194]}
   );
   gpc1_1 gpc5109 (
      {stage0_49[465]},
      {stage1_49[195]}
   );
   gpc1_1 gpc5110 (
      {stage0_49[466]},
      {stage1_49[196]}
   );
   gpc1_1 gpc5111 (
      {stage0_49[467]},
      {stage1_49[197]}
   );
   gpc1_1 gpc5112 (
      {stage0_49[468]},
      {stage1_49[198]}
   );
   gpc1_1 gpc5113 (
      {stage0_49[469]},
      {stage1_49[199]}
   );
   gpc1_1 gpc5114 (
      {stage0_49[470]},
      {stage1_49[200]}
   );
   gpc1_1 gpc5115 (
      {stage0_49[471]},
      {stage1_49[201]}
   );
   gpc1_1 gpc5116 (
      {stage0_49[472]},
      {stage1_49[202]}
   );
   gpc1_1 gpc5117 (
      {stage0_49[473]},
      {stage1_49[203]}
   );
   gpc1_1 gpc5118 (
      {stage0_49[474]},
      {stage1_49[204]}
   );
   gpc1_1 gpc5119 (
      {stage0_49[475]},
      {stage1_49[205]}
   );
   gpc1_1 gpc5120 (
      {stage0_49[476]},
      {stage1_49[206]}
   );
   gpc1_1 gpc5121 (
      {stage0_49[477]},
      {stage1_49[207]}
   );
   gpc1_1 gpc5122 (
      {stage0_49[478]},
      {stage1_49[208]}
   );
   gpc1_1 gpc5123 (
      {stage0_49[479]},
      {stage1_49[209]}
   );
   gpc1_1 gpc5124 (
      {stage0_49[480]},
      {stage1_49[210]}
   );
   gpc1_1 gpc5125 (
      {stage0_49[481]},
      {stage1_49[211]}
   );
   gpc1_1 gpc5126 (
      {stage0_49[482]},
      {stage1_49[212]}
   );
   gpc1_1 gpc5127 (
      {stage0_49[483]},
      {stage1_49[213]}
   );
   gpc1_1 gpc5128 (
      {stage0_49[484]},
      {stage1_49[214]}
   );
   gpc1_1 gpc5129 (
      {stage0_49[485]},
      {stage1_49[215]}
   );
   gpc1_1 gpc5130 (
      {stage0_49[486]},
      {stage1_49[216]}
   );
   gpc1_1 gpc5131 (
      {stage0_49[487]},
      {stage1_49[217]}
   );
   gpc1_1 gpc5132 (
      {stage0_49[488]},
      {stage1_49[218]}
   );
   gpc1_1 gpc5133 (
      {stage0_49[489]},
      {stage1_49[219]}
   );
   gpc1_1 gpc5134 (
      {stage0_49[490]},
      {stage1_49[220]}
   );
   gpc1_1 gpc5135 (
      {stage0_49[491]},
      {stage1_49[221]}
   );
   gpc1_1 gpc5136 (
      {stage0_49[492]},
      {stage1_49[222]}
   );
   gpc1_1 gpc5137 (
      {stage0_49[493]},
      {stage1_49[223]}
   );
   gpc1_1 gpc5138 (
      {stage0_49[494]},
      {stage1_49[224]}
   );
   gpc1_1 gpc5139 (
      {stage0_49[495]},
      {stage1_49[225]}
   );
   gpc1_1 gpc5140 (
      {stage0_49[496]},
      {stage1_49[226]}
   );
   gpc1_1 gpc5141 (
      {stage0_49[497]},
      {stage1_49[227]}
   );
   gpc1_1 gpc5142 (
      {stage0_49[498]},
      {stage1_49[228]}
   );
   gpc1_1 gpc5143 (
      {stage0_49[499]},
      {stage1_49[229]}
   );
   gpc1_1 gpc5144 (
      {stage0_49[500]},
      {stage1_49[230]}
   );
   gpc1_1 gpc5145 (
      {stage0_49[501]},
      {stage1_49[231]}
   );
   gpc1_1 gpc5146 (
      {stage0_49[502]},
      {stage1_49[232]}
   );
   gpc1_1 gpc5147 (
      {stage0_49[503]},
      {stage1_49[233]}
   );
   gpc1_1 gpc5148 (
      {stage0_49[504]},
      {stage1_49[234]}
   );
   gpc1_1 gpc5149 (
      {stage0_49[505]},
      {stage1_49[235]}
   );
   gpc1_1 gpc5150 (
      {stage0_49[506]},
      {stage1_49[236]}
   );
   gpc1_1 gpc5151 (
      {stage0_49[507]},
      {stage1_49[237]}
   );
   gpc1_1 gpc5152 (
      {stage0_49[508]},
      {stage1_49[238]}
   );
   gpc1_1 gpc5153 (
      {stage0_49[509]},
      {stage1_49[239]}
   );
   gpc1_1 gpc5154 (
      {stage0_49[510]},
      {stage1_49[240]}
   );
   gpc1_1 gpc5155 (
      {stage0_49[511]},
      {stage1_49[241]}
   );
   gpc1_1 gpc5156 (
      {stage0_50[474]},
      {stage1_50[179]}
   );
   gpc1_1 gpc5157 (
      {stage0_50[475]},
      {stage1_50[180]}
   );
   gpc1_1 gpc5158 (
      {stage0_50[476]},
      {stage1_50[181]}
   );
   gpc1_1 gpc5159 (
      {stage0_50[477]},
      {stage1_50[182]}
   );
   gpc1_1 gpc5160 (
      {stage0_50[478]},
      {stage1_50[183]}
   );
   gpc1_1 gpc5161 (
      {stage0_50[479]},
      {stage1_50[184]}
   );
   gpc1_1 gpc5162 (
      {stage0_50[480]},
      {stage1_50[185]}
   );
   gpc1_1 gpc5163 (
      {stage0_50[481]},
      {stage1_50[186]}
   );
   gpc1_1 gpc5164 (
      {stage0_50[482]},
      {stage1_50[187]}
   );
   gpc1_1 gpc5165 (
      {stage0_50[483]},
      {stage1_50[188]}
   );
   gpc1_1 gpc5166 (
      {stage0_50[484]},
      {stage1_50[189]}
   );
   gpc1_1 gpc5167 (
      {stage0_50[485]},
      {stage1_50[190]}
   );
   gpc1_1 gpc5168 (
      {stage0_50[486]},
      {stage1_50[191]}
   );
   gpc1_1 gpc5169 (
      {stage0_50[487]},
      {stage1_50[192]}
   );
   gpc1_1 gpc5170 (
      {stage0_50[488]},
      {stage1_50[193]}
   );
   gpc1_1 gpc5171 (
      {stage0_50[489]},
      {stage1_50[194]}
   );
   gpc1_1 gpc5172 (
      {stage0_50[490]},
      {stage1_50[195]}
   );
   gpc1_1 gpc5173 (
      {stage0_50[491]},
      {stage1_50[196]}
   );
   gpc1_1 gpc5174 (
      {stage0_50[492]},
      {stage1_50[197]}
   );
   gpc1_1 gpc5175 (
      {stage0_50[493]},
      {stage1_50[198]}
   );
   gpc1_1 gpc5176 (
      {stage0_50[494]},
      {stage1_50[199]}
   );
   gpc1_1 gpc5177 (
      {stage0_50[495]},
      {stage1_50[200]}
   );
   gpc1_1 gpc5178 (
      {stage0_50[496]},
      {stage1_50[201]}
   );
   gpc1_1 gpc5179 (
      {stage0_50[497]},
      {stage1_50[202]}
   );
   gpc1_1 gpc5180 (
      {stage0_50[498]},
      {stage1_50[203]}
   );
   gpc1_1 gpc5181 (
      {stage0_50[499]},
      {stage1_50[204]}
   );
   gpc1_1 gpc5182 (
      {stage0_50[500]},
      {stage1_50[205]}
   );
   gpc1_1 gpc5183 (
      {stage0_50[501]},
      {stage1_50[206]}
   );
   gpc1_1 gpc5184 (
      {stage0_50[502]},
      {stage1_50[207]}
   );
   gpc1_1 gpc5185 (
      {stage0_50[503]},
      {stage1_50[208]}
   );
   gpc1_1 gpc5186 (
      {stage0_50[504]},
      {stage1_50[209]}
   );
   gpc1_1 gpc5187 (
      {stage0_50[505]},
      {stage1_50[210]}
   );
   gpc1_1 gpc5188 (
      {stage0_50[506]},
      {stage1_50[211]}
   );
   gpc1_1 gpc5189 (
      {stage0_50[507]},
      {stage1_50[212]}
   );
   gpc1_1 gpc5190 (
      {stage0_50[508]},
      {stage1_50[213]}
   );
   gpc1_1 gpc5191 (
      {stage0_50[509]},
      {stage1_50[214]}
   );
   gpc1_1 gpc5192 (
      {stage0_50[510]},
      {stage1_50[215]}
   );
   gpc1_1 gpc5193 (
      {stage0_50[511]},
      {stage1_50[216]}
   );
   gpc1_1 gpc5194 (
      {stage0_51[501]},
      {stage1_51[216]}
   );
   gpc1_1 gpc5195 (
      {stage0_51[502]},
      {stage1_51[217]}
   );
   gpc1_1 gpc5196 (
      {stage0_51[503]},
      {stage1_51[218]}
   );
   gpc1_1 gpc5197 (
      {stage0_51[504]},
      {stage1_51[219]}
   );
   gpc1_1 gpc5198 (
      {stage0_51[505]},
      {stage1_51[220]}
   );
   gpc1_1 gpc5199 (
      {stage0_51[506]},
      {stage1_51[221]}
   );
   gpc1_1 gpc5200 (
      {stage0_51[507]},
      {stage1_51[222]}
   );
   gpc1_1 gpc5201 (
      {stage0_51[508]},
      {stage1_51[223]}
   );
   gpc1_1 gpc5202 (
      {stage0_51[509]},
      {stage1_51[224]}
   );
   gpc1_1 gpc5203 (
      {stage0_51[510]},
      {stage1_51[225]}
   );
   gpc1_1 gpc5204 (
      {stage0_51[511]},
      {stage1_51[226]}
   );
   gpc1_1 gpc5205 (
      {stage0_52[410]},
      {stage1_52[202]}
   );
   gpc1_1 gpc5206 (
      {stage0_52[411]},
      {stage1_52[203]}
   );
   gpc1_1 gpc5207 (
      {stage0_52[412]},
      {stage1_52[204]}
   );
   gpc1_1 gpc5208 (
      {stage0_52[413]},
      {stage1_52[205]}
   );
   gpc1_1 gpc5209 (
      {stage0_52[414]},
      {stage1_52[206]}
   );
   gpc1_1 gpc5210 (
      {stage0_52[415]},
      {stage1_52[207]}
   );
   gpc1_1 gpc5211 (
      {stage0_52[416]},
      {stage1_52[208]}
   );
   gpc1_1 gpc5212 (
      {stage0_52[417]},
      {stage1_52[209]}
   );
   gpc1_1 gpc5213 (
      {stage0_52[418]},
      {stage1_52[210]}
   );
   gpc1_1 gpc5214 (
      {stage0_52[419]},
      {stage1_52[211]}
   );
   gpc1_1 gpc5215 (
      {stage0_52[420]},
      {stage1_52[212]}
   );
   gpc1_1 gpc5216 (
      {stage0_52[421]},
      {stage1_52[213]}
   );
   gpc1_1 gpc5217 (
      {stage0_52[422]},
      {stage1_52[214]}
   );
   gpc1_1 gpc5218 (
      {stage0_52[423]},
      {stage1_52[215]}
   );
   gpc1_1 gpc5219 (
      {stage0_52[424]},
      {stage1_52[216]}
   );
   gpc1_1 gpc5220 (
      {stage0_52[425]},
      {stage1_52[217]}
   );
   gpc1_1 gpc5221 (
      {stage0_52[426]},
      {stage1_52[218]}
   );
   gpc1_1 gpc5222 (
      {stage0_52[427]},
      {stage1_52[219]}
   );
   gpc1_1 gpc5223 (
      {stage0_52[428]},
      {stage1_52[220]}
   );
   gpc1_1 gpc5224 (
      {stage0_52[429]},
      {stage1_52[221]}
   );
   gpc1_1 gpc5225 (
      {stage0_52[430]},
      {stage1_52[222]}
   );
   gpc1_1 gpc5226 (
      {stage0_52[431]},
      {stage1_52[223]}
   );
   gpc1_1 gpc5227 (
      {stage0_52[432]},
      {stage1_52[224]}
   );
   gpc1_1 gpc5228 (
      {stage0_52[433]},
      {stage1_52[225]}
   );
   gpc1_1 gpc5229 (
      {stage0_52[434]},
      {stage1_52[226]}
   );
   gpc1_1 gpc5230 (
      {stage0_52[435]},
      {stage1_52[227]}
   );
   gpc1_1 gpc5231 (
      {stage0_52[436]},
      {stage1_52[228]}
   );
   gpc1_1 gpc5232 (
      {stage0_52[437]},
      {stage1_52[229]}
   );
   gpc1_1 gpc5233 (
      {stage0_52[438]},
      {stage1_52[230]}
   );
   gpc1_1 gpc5234 (
      {stage0_52[439]},
      {stage1_52[231]}
   );
   gpc1_1 gpc5235 (
      {stage0_52[440]},
      {stage1_52[232]}
   );
   gpc1_1 gpc5236 (
      {stage0_52[441]},
      {stage1_52[233]}
   );
   gpc1_1 gpc5237 (
      {stage0_52[442]},
      {stage1_52[234]}
   );
   gpc1_1 gpc5238 (
      {stage0_52[443]},
      {stage1_52[235]}
   );
   gpc1_1 gpc5239 (
      {stage0_52[444]},
      {stage1_52[236]}
   );
   gpc1_1 gpc5240 (
      {stage0_52[445]},
      {stage1_52[237]}
   );
   gpc1_1 gpc5241 (
      {stage0_52[446]},
      {stage1_52[238]}
   );
   gpc1_1 gpc5242 (
      {stage0_52[447]},
      {stage1_52[239]}
   );
   gpc1_1 gpc5243 (
      {stage0_52[448]},
      {stage1_52[240]}
   );
   gpc1_1 gpc5244 (
      {stage0_52[449]},
      {stage1_52[241]}
   );
   gpc1_1 gpc5245 (
      {stage0_52[450]},
      {stage1_52[242]}
   );
   gpc1_1 gpc5246 (
      {stage0_52[451]},
      {stage1_52[243]}
   );
   gpc1_1 gpc5247 (
      {stage0_52[452]},
      {stage1_52[244]}
   );
   gpc1_1 gpc5248 (
      {stage0_52[453]},
      {stage1_52[245]}
   );
   gpc1_1 gpc5249 (
      {stage0_52[454]},
      {stage1_52[246]}
   );
   gpc1_1 gpc5250 (
      {stage0_52[455]},
      {stage1_52[247]}
   );
   gpc1_1 gpc5251 (
      {stage0_52[456]},
      {stage1_52[248]}
   );
   gpc1_1 gpc5252 (
      {stage0_52[457]},
      {stage1_52[249]}
   );
   gpc1_1 gpc5253 (
      {stage0_52[458]},
      {stage1_52[250]}
   );
   gpc1_1 gpc5254 (
      {stage0_52[459]},
      {stage1_52[251]}
   );
   gpc1_1 gpc5255 (
      {stage0_52[460]},
      {stage1_52[252]}
   );
   gpc1_1 gpc5256 (
      {stage0_52[461]},
      {stage1_52[253]}
   );
   gpc1_1 gpc5257 (
      {stage0_52[462]},
      {stage1_52[254]}
   );
   gpc1_1 gpc5258 (
      {stage0_52[463]},
      {stage1_52[255]}
   );
   gpc1_1 gpc5259 (
      {stage0_52[464]},
      {stage1_52[256]}
   );
   gpc1_1 gpc5260 (
      {stage0_52[465]},
      {stage1_52[257]}
   );
   gpc1_1 gpc5261 (
      {stage0_52[466]},
      {stage1_52[258]}
   );
   gpc1_1 gpc5262 (
      {stage0_52[467]},
      {stage1_52[259]}
   );
   gpc1_1 gpc5263 (
      {stage0_52[468]},
      {stage1_52[260]}
   );
   gpc1_1 gpc5264 (
      {stage0_52[469]},
      {stage1_52[261]}
   );
   gpc1_1 gpc5265 (
      {stage0_52[470]},
      {stage1_52[262]}
   );
   gpc1_1 gpc5266 (
      {stage0_52[471]},
      {stage1_52[263]}
   );
   gpc1_1 gpc5267 (
      {stage0_52[472]},
      {stage1_52[264]}
   );
   gpc1_1 gpc5268 (
      {stage0_52[473]},
      {stage1_52[265]}
   );
   gpc1_1 gpc5269 (
      {stage0_52[474]},
      {stage1_52[266]}
   );
   gpc1_1 gpc5270 (
      {stage0_52[475]},
      {stage1_52[267]}
   );
   gpc1_1 gpc5271 (
      {stage0_52[476]},
      {stage1_52[268]}
   );
   gpc1_1 gpc5272 (
      {stage0_52[477]},
      {stage1_52[269]}
   );
   gpc1_1 gpc5273 (
      {stage0_52[478]},
      {stage1_52[270]}
   );
   gpc1_1 gpc5274 (
      {stage0_52[479]},
      {stage1_52[271]}
   );
   gpc1_1 gpc5275 (
      {stage0_52[480]},
      {stage1_52[272]}
   );
   gpc1_1 gpc5276 (
      {stage0_52[481]},
      {stage1_52[273]}
   );
   gpc1_1 gpc5277 (
      {stage0_52[482]},
      {stage1_52[274]}
   );
   gpc1_1 gpc5278 (
      {stage0_52[483]},
      {stage1_52[275]}
   );
   gpc1_1 gpc5279 (
      {stage0_52[484]},
      {stage1_52[276]}
   );
   gpc1_1 gpc5280 (
      {stage0_52[485]},
      {stage1_52[277]}
   );
   gpc1_1 gpc5281 (
      {stage0_52[486]},
      {stage1_52[278]}
   );
   gpc1_1 gpc5282 (
      {stage0_52[487]},
      {stage1_52[279]}
   );
   gpc1_1 gpc5283 (
      {stage0_52[488]},
      {stage1_52[280]}
   );
   gpc1_1 gpc5284 (
      {stage0_52[489]},
      {stage1_52[281]}
   );
   gpc1_1 gpc5285 (
      {stage0_52[490]},
      {stage1_52[282]}
   );
   gpc1_1 gpc5286 (
      {stage0_52[491]},
      {stage1_52[283]}
   );
   gpc1_1 gpc5287 (
      {stage0_52[492]},
      {stage1_52[284]}
   );
   gpc1_1 gpc5288 (
      {stage0_52[493]},
      {stage1_52[285]}
   );
   gpc1_1 gpc5289 (
      {stage0_52[494]},
      {stage1_52[286]}
   );
   gpc1_1 gpc5290 (
      {stage0_52[495]},
      {stage1_52[287]}
   );
   gpc1_1 gpc5291 (
      {stage0_52[496]},
      {stage1_52[288]}
   );
   gpc1_1 gpc5292 (
      {stage0_52[497]},
      {stage1_52[289]}
   );
   gpc1_1 gpc5293 (
      {stage0_52[498]},
      {stage1_52[290]}
   );
   gpc1_1 gpc5294 (
      {stage0_52[499]},
      {stage1_52[291]}
   );
   gpc1_1 gpc5295 (
      {stage0_52[500]},
      {stage1_52[292]}
   );
   gpc1_1 gpc5296 (
      {stage0_52[501]},
      {stage1_52[293]}
   );
   gpc1_1 gpc5297 (
      {stage0_52[502]},
      {stage1_52[294]}
   );
   gpc1_1 gpc5298 (
      {stage0_52[503]},
      {stage1_52[295]}
   );
   gpc1_1 gpc5299 (
      {stage0_52[504]},
      {stage1_52[296]}
   );
   gpc1_1 gpc5300 (
      {stage0_52[505]},
      {stage1_52[297]}
   );
   gpc1_1 gpc5301 (
      {stage0_52[506]},
      {stage1_52[298]}
   );
   gpc1_1 gpc5302 (
      {stage0_52[507]},
      {stage1_52[299]}
   );
   gpc1_1 gpc5303 (
      {stage0_52[508]},
      {stage1_52[300]}
   );
   gpc1_1 gpc5304 (
      {stage0_52[509]},
      {stage1_52[301]}
   );
   gpc1_1 gpc5305 (
      {stage0_52[510]},
      {stage1_52[302]}
   );
   gpc1_1 gpc5306 (
      {stage0_52[511]},
      {stage1_52[303]}
   );
   gpc1_1 gpc5307 (
      {stage0_53[497]},
      {stage1_53[172]}
   );
   gpc1_1 gpc5308 (
      {stage0_53[498]},
      {stage1_53[173]}
   );
   gpc1_1 gpc5309 (
      {stage0_53[499]},
      {stage1_53[174]}
   );
   gpc1_1 gpc5310 (
      {stage0_53[500]},
      {stage1_53[175]}
   );
   gpc1_1 gpc5311 (
      {stage0_53[501]},
      {stage1_53[176]}
   );
   gpc1_1 gpc5312 (
      {stage0_53[502]},
      {stage1_53[177]}
   );
   gpc1_1 gpc5313 (
      {stage0_53[503]},
      {stage1_53[178]}
   );
   gpc1_1 gpc5314 (
      {stage0_53[504]},
      {stage1_53[179]}
   );
   gpc1_1 gpc5315 (
      {stage0_53[505]},
      {stage1_53[180]}
   );
   gpc1_1 gpc5316 (
      {stage0_53[506]},
      {stage1_53[181]}
   );
   gpc1_1 gpc5317 (
      {stage0_53[507]},
      {stage1_53[182]}
   );
   gpc1_1 gpc5318 (
      {stage0_53[508]},
      {stage1_53[183]}
   );
   gpc1_1 gpc5319 (
      {stage0_53[509]},
      {stage1_53[184]}
   );
   gpc1_1 gpc5320 (
      {stage0_53[510]},
      {stage1_53[185]}
   );
   gpc1_1 gpc5321 (
      {stage0_53[511]},
      {stage1_53[186]}
   );
   gpc1_1 gpc5322 (
      {stage0_54[441]},
      {stage1_54[192]}
   );
   gpc1_1 gpc5323 (
      {stage0_54[442]},
      {stage1_54[193]}
   );
   gpc1_1 gpc5324 (
      {stage0_54[443]},
      {stage1_54[194]}
   );
   gpc1_1 gpc5325 (
      {stage0_54[444]},
      {stage1_54[195]}
   );
   gpc1_1 gpc5326 (
      {stage0_54[445]},
      {stage1_54[196]}
   );
   gpc1_1 gpc5327 (
      {stage0_54[446]},
      {stage1_54[197]}
   );
   gpc1_1 gpc5328 (
      {stage0_54[447]},
      {stage1_54[198]}
   );
   gpc1_1 gpc5329 (
      {stage0_54[448]},
      {stage1_54[199]}
   );
   gpc1_1 gpc5330 (
      {stage0_54[449]},
      {stage1_54[200]}
   );
   gpc1_1 gpc5331 (
      {stage0_54[450]},
      {stage1_54[201]}
   );
   gpc1_1 gpc5332 (
      {stage0_54[451]},
      {stage1_54[202]}
   );
   gpc1_1 gpc5333 (
      {stage0_54[452]},
      {stage1_54[203]}
   );
   gpc1_1 gpc5334 (
      {stage0_54[453]},
      {stage1_54[204]}
   );
   gpc1_1 gpc5335 (
      {stage0_54[454]},
      {stage1_54[205]}
   );
   gpc1_1 gpc5336 (
      {stage0_54[455]},
      {stage1_54[206]}
   );
   gpc1_1 gpc5337 (
      {stage0_54[456]},
      {stage1_54[207]}
   );
   gpc1_1 gpc5338 (
      {stage0_54[457]},
      {stage1_54[208]}
   );
   gpc1_1 gpc5339 (
      {stage0_54[458]},
      {stage1_54[209]}
   );
   gpc1_1 gpc5340 (
      {stage0_54[459]},
      {stage1_54[210]}
   );
   gpc1_1 gpc5341 (
      {stage0_54[460]},
      {stage1_54[211]}
   );
   gpc1_1 gpc5342 (
      {stage0_54[461]},
      {stage1_54[212]}
   );
   gpc1_1 gpc5343 (
      {stage0_54[462]},
      {stage1_54[213]}
   );
   gpc1_1 gpc5344 (
      {stage0_54[463]},
      {stage1_54[214]}
   );
   gpc1_1 gpc5345 (
      {stage0_54[464]},
      {stage1_54[215]}
   );
   gpc1_1 gpc5346 (
      {stage0_54[465]},
      {stage1_54[216]}
   );
   gpc1_1 gpc5347 (
      {stage0_54[466]},
      {stage1_54[217]}
   );
   gpc1_1 gpc5348 (
      {stage0_54[467]},
      {stage1_54[218]}
   );
   gpc1_1 gpc5349 (
      {stage0_54[468]},
      {stage1_54[219]}
   );
   gpc1_1 gpc5350 (
      {stage0_54[469]},
      {stage1_54[220]}
   );
   gpc1_1 gpc5351 (
      {stage0_54[470]},
      {stage1_54[221]}
   );
   gpc1_1 gpc5352 (
      {stage0_54[471]},
      {stage1_54[222]}
   );
   gpc1_1 gpc5353 (
      {stage0_54[472]},
      {stage1_54[223]}
   );
   gpc1_1 gpc5354 (
      {stage0_54[473]},
      {stage1_54[224]}
   );
   gpc1_1 gpc5355 (
      {stage0_54[474]},
      {stage1_54[225]}
   );
   gpc1_1 gpc5356 (
      {stage0_54[475]},
      {stage1_54[226]}
   );
   gpc1_1 gpc5357 (
      {stage0_54[476]},
      {stage1_54[227]}
   );
   gpc1_1 gpc5358 (
      {stage0_54[477]},
      {stage1_54[228]}
   );
   gpc1_1 gpc5359 (
      {stage0_54[478]},
      {stage1_54[229]}
   );
   gpc1_1 gpc5360 (
      {stage0_54[479]},
      {stage1_54[230]}
   );
   gpc1_1 gpc5361 (
      {stage0_54[480]},
      {stage1_54[231]}
   );
   gpc1_1 gpc5362 (
      {stage0_54[481]},
      {stage1_54[232]}
   );
   gpc1_1 gpc5363 (
      {stage0_54[482]},
      {stage1_54[233]}
   );
   gpc1_1 gpc5364 (
      {stage0_54[483]},
      {stage1_54[234]}
   );
   gpc1_1 gpc5365 (
      {stage0_54[484]},
      {stage1_54[235]}
   );
   gpc1_1 gpc5366 (
      {stage0_54[485]},
      {stage1_54[236]}
   );
   gpc1_1 gpc5367 (
      {stage0_54[486]},
      {stage1_54[237]}
   );
   gpc1_1 gpc5368 (
      {stage0_54[487]},
      {stage1_54[238]}
   );
   gpc1_1 gpc5369 (
      {stage0_54[488]},
      {stage1_54[239]}
   );
   gpc1_1 gpc5370 (
      {stage0_54[489]},
      {stage1_54[240]}
   );
   gpc1_1 gpc5371 (
      {stage0_54[490]},
      {stage1_54[241]}
   );
   gpc1_1 gpc5372 (
      {stage0_54[491]},
      {stage1_54[242]}
   );
   gpc1_1 gpc5373 (
      {stage0_54[492]},
      {stage1_54[243]}
   );
   gpc1_1 gpc5374 (
      {stage0_54[493]},
      {stage1_54[244]}
   );
   gpc1_1 gpc5375 (
      {stage0_54[494]},
      {stage1_54[245]}
   );
   gpc1_1 gpc5376 (
      {stage0_54[495]},
      {stage1_54[246]}
   );
   gpc1_1 gpc5377 (
      {stage0_54[496]},
      {stage1_54[247]}
   );
   gpc1_1 gpc5378 (
      {stage0_54[497]},
      {stage1_54[248]}
   );
   gpc1_1 gpc5379 (
      {stage0_54[498]},
      {stage1_54[249]}
   );
   gpc1_1 gpc5380 (
      {stage0_54[499]},
      {stage1_54[250]}
   );
   gpc1_1 gpc5381 (
      {stage0_54[500]},
      {stage1_54[251]}
   );
   gpc1_1 gpc5382 (
      {stage0_54[501]},
      {stage1_54[252]}
   );
   gpc1_1 gpc5383 (
      {stage0_54[502]},
      {stage1_54[253]}
   );
   gpc1_1 gpc5384 (
      {stage0_54[503]},
      {stage1_54[254]}
   );
   gpc1_1 gpc5385 (
      {stage0_54[504]},
      {stage1_54[255]}
   );
   gpc1_1 gpc5386 (
      {stage0_54[505]},
      {stage1_54[256]}
   );
   gpc1_1 gpc5387 (
      {stage0_54[506]},
      {stage1_54[257]}
   );
   gpc1_1 gpc5388 (
      {stage0_54[507]},
      {stage1_54[258]}
   );
   gpc1_1 gpc5389 (
      {stage0_54[508]},
      {stage1_54[259]}
   );
   gpc1_1 gpc5390 (
      {stage0_54[509]},
      {stage1_54[260]}
   );
   gpc1_1 gpc5391 (
      {stage0_54[510]},
      {stage1_54[261]}
   );
   gpc1_1 gpc5392 (
      {stage0_54[511]},
      {stage1_54[262]}
   );
   gpc1_1 gpc5393 (
      {stage0_55[508]},
      {stage1_55[222]}
   );
   gpc1_1 gpc5394 (
      {stage0_55[509]},
      {stage1_55[223]}
   );
   gpc1_1 gpc5395 (
      {stage0_55[510]},
      {stage1_55[224]}
   );
   gpc1_1 gpc5396 (
      {stage0_55[511]},
      {stage1_55[225]}
   );
   gpc1_1 gpc5397 (
      {stage0_56[444]},
      {stage1_56[189]}
   );
   gpc1_1 gpc5398 (
      {stage0_56[445]},
      {stage1_56[190]}
   );
   gpc1_1 gpc5399 (
      {stage0_56[446]},
      {stage1_56[191]}
   );
   gpc1_1 gpc5400 (
      {stage0_56[447]},
      {stage1_56[192]}
   );
   gpc1_1 gpc5401 (
      {stage0_56[448]},
      {stage1_56[193]}
   );
   gpc1_1 gpc5402 (
      {stage0_56[449]},
      {stage1_56[194]}
   );
   gpc1_1 gpc5403 (
      {stage0_56[450]},
      {stage1_56[195]}
   );
   gpc1_1 gpc5404 (
      {stage0_56[451]},
      {stage1_56[196]}
   );
   gpc1_1 gpc5405 (
      {stage0_56[452]},
      {stage1_56[197]}
   );
   gpc1_1 gpc5406 (
      {stage0_56[453]},
      {stage1_56[198]}
   );
   gpc1_1 gpc5407 (
      {stage0_56[454]},
      {stage1_56[199]}
   );
   gpc1_1 gpc5408 (
      {stage0_56[455]},
      {stage1_56[200]}
   );
   gpc1_1 gpc5409 (
      {stage0_56[456]},
      {stage1_56[201]}
   );
   gpc1_1 gpc5410 (
      {stage0_56[457]},
      {stage1_56[202]}
   );
   gpc1_1 gpc5411 (
      {stage0_56[458]},
      {stage1_56[203]}
   );
   gpc1_1 gpc5412 (
      {stage0_56[459]},
      {stage1_56[204]}
   );
   gpc1_1 gpc5413 (
      {stage0_56[460]},
      {stage1_56[205]}
   );
   gpc1_1 gpc5414 (
      {stage0_56[461]},
      {stage1_56[206]}
   );
   gpc1_1 gpc5415 (
      {stage0_56[462]},
      {stage1_56[207]}
   );
   gpc1_1 gpc5416 (
      {stage0_56[463]},
      {stage1_56[208]}
   );
   gpc1_1 gpc5417 (
      {stage0_56[464]},
      {stage1_56[209]}
   );
   gpc1_1 gpc5418 (
      {stage0_56[465]},
      {stage1_56[210]}
   );
   gpc1_1 gpc5419 (
      {stage0_56[466]},
      {stage1_56[211]}
   );
   gpc1_1 gpc5420 (
      {stage0_56[467]},
      {stage1_56[212]}
   );
   gpc1_1 gpc5421 (
      {stage0_56[468]},
      {stage1_56[213]}
   );
   gpc1_1 gpc5422 (
      {stage0_56[469]},
      {stage1_56[214]}
   );
   gpc1_1 gpc5423 (
      {stage0_56[470]},
      {stage1_56[215]}
   );
   gpc1_1 gpc5424 (
      {stage0_56[471]},
      {stage1_56[216]}
   );
   gpc1_1 gpc5425 (
      {stage0_56[472]},
      {stage1_56[217]}
   );
   gpc1_1 gpc5426 (
      {stage0_56[473]},
      {stage1_56[218]}
   );
   gpc1_1 gpc5427 (
      {stage0_56[474]},
      {stage1_56[219]}
   );
   gpc1_1 gpc5428 (
      {stage0_56[475]},
      {stage1_56[220]}
   );
   gpc1_1 gpc5429 (
      {stage0_56[476]},
      {stage1_56[221]}
   );
   gpc1_1 gpc5430 (
      {stage0_56[477]},
      {stage1_56[222]}
   );
   gpc1_1 gpc5431 (
      {stage0_56[478]},
      {stage1_56[223]}
   );
   gpc1_1 gpc5432 (
      {stage0_56[479]},
      {stage1_56[224]}
   );
   gpc1_1 gpc5433 (
      {stage0_56[480]},
      {stage1_56[225]}
   );
   gpc1_1 gpc5434 (
      {stage0_56[481]},
      {stage1_56[226]}
   );
   gpc1_1 gpc5435 (
      {stage0_56[482]},
      {stage1_56[227]}
   );
   gpc1_1 gpc5436 (
      {stage0_56[483]},
      {stage1_56[228]}
   );
   gpc1_1 gpc5437 (
      {stage0_56[484]},
      {stage1_56[229]}
   );
   gpc1_1 gpc5438 (
      {stage0_56[485]},
      {stage1_56[230]}
   );
   gpc1_1 gpc5439 (
      {stage0_56[486]},
      {stage1_56[231]}
   );
   gpc1_1 gpc5440 (
      {stage0_56[487]},
      {stage1_56[232]}
   );
   gpc1_1 gpc5441 (
      {stage0_56[488]},
      {stage1_56[233]}
   );
   gpc1_1 gpc5442 (
      {stage0_56[489]},
      {stage1_56[234]}
   );
   gpc1_1 gpc5443 (
      {stage0_56[490]},
      {stage1_56[235]}
   );
   gpc1_1 gpc5444 (
      {stage0_56[491]},
      {stage1_56[236]}
   );
   gpc1_1 gpc5445 (
      {stage0_56[492]},
      {stage1_56[237]}
   );
   gpc1_1 gpc5446 (
      {stage0_56[493]},
      {stage1_56[238]}
   );
   gpc1_1 gpc5447 (
      {stage0_56[494]},
      {stage1_56[239]}
   );
   gpc1_1 gpc5448 (
      {stage0_56[495]},
      {stage1_56[240]}
   );
   gpc1_1 gpc5449 (
      {stage0_56[496]},
      {stage1_56[241]}
   );
   gpc1_1 gpc5450 (
      {stage0_56[497]},
      {stage1_56[242]}
   );
   gpc1_1 gpc5451 (
      {stage0_56[498]},
      {stage1_56[243]}
   );
   gpc1_1 gpc5452 (
      {stage0_56[499]},
      {stage1_56[244]}
   );
   gpc1_1 gpc5453 (
      {stage0_56[500]},
      {stage1_56[245]}
   );
   gpc1_1 gpc5454 (
      {stage0_56[501]},
      {stage1_56[246]}
   );
   gpc1_1 gpc5455 (
      {stage0_56[502]},
      {stage1_56[247]}
   );
   gpc1_1 gpc5456 (
      {stage0_56[503]},
      {stage1_56[248]}
   );
   gpc1_1 gpc5457 (
      {stage0_56[504]},
      {stage1_56[249]}
   );
   gpc1_1 gpc5458 (
      {stage0_56[505]},
      {stage1_56[250]}
   );
   gpc1_1 gpc5459 (
      {stage0_56[506]},
      {stage1_56[251]}
   );
   gpc1_1 gpc5460 (
      {stage0_56[507]},
      {stage1_56[252]}
   );
   gpc1_1 gpc5461 (
      {stage0_56[508]},
      {stage1_56[253]}
   );
   gpc1_1 gpc5462 (
      {stage0_56[509]},
      {stage1_56[254]}
   );
   gpc1_1 gpc5463 (
      {stage0_56[510]},
      {stage1_56[255]}
   );
   gpc1_1 gpc5464 (
      {stage0_56[511]},
      {stage1_56[256]}
   );
   gpc1_1 gpc5465 (
      {stage0_57[510]},
      {stage1_57[178]}
   );
   gpc1_1 gpc5466 (
      {stage0_57[511]},
      {stage1_57[179]}
   );
   gpc1_1 gpc5467 (
      {stage0_58[493]},
      {stage1_58[224]}
   );
   gpc1_1 gpc5468 (
      {stage0_58[494]},
      {stage1_58[225]}
   );
   gpc1_1 gpc5469 (
      {stage0_58[495]},
      {stage1_58[226]}
   );
   gpc1_1 gpc5470 (
      {stage0_58[496]},
      {stage1_58[227]}
   );
   gpc1_1 gpc5471 (
      {stage0_58[497]},
      {stage1_58[228]}
   );
   gpc1_1 gpc5472 (
      {stage0_58[498]},
      {stage1_58[229]}
   );
   gpc1_1 gpc5473 (
      {stage0_58[499]},
      {stage1_58[230]}
   );
   gpc1_1 gpc5474 (
      {stage0_58[500]},
      {stage1_58[231]}
   );
   gpc1_1 gpc5475 (
      {stage0_58[501]},
      {stage1_58[232]}
   );
   gpc1_1 gpc5476 (
      {stage0_58[502]},
      {stage1_58[233]}
   );
   gpc1_1 gpc5477 (
      {stage0_58[503]},
      {stage1_58[234]}
   );
   gpc1_1 gpc5478 (
      {stage0_58[504]},
      {stage1_58[235]}
   );
   gpc1_1 gpc5479 (
      {stage0_58[505]},
      {stage1_58[236]}
   );
   gpc1_1 gpc5480 (
      {stage0_58[506]},
      {stage1_58[237]}
   );
   gpc1_1 gpc5481 (
      {stage0_58[507]},
      {stage1_58[238]}
   );
   gpc1_1 gpc5482 (
      {stage0_58[508]},
      {stage1_58[239]}
   );
   gpc1_1 gpc5483 (
      {stage0_58[509]},
      {stage1_58[240]}
   );
   gpc1_1 gpc5484 (
      {stage0_58[510]},
      {stage1_58[241]}
   );
   gpc1_1 gpc5485 (
      {stage0_58[511]},
      {stage1_58[242]}
   );
   gpc1_1 gpc5486 (
      {stage0_59[412]},
      {stage1_59[194]}
   );
   gpc1_1 gpc5487 (
      {stage0_59[413]},
      {stage1_59[195]}
   );
   gpc1_1 gpc5488 (
      {stage0_59[414]},
      {stage1_59[196]}
   );
   gpc1_1 gpc5489 (
      {stage0_59[415]},
      {stage1_59[197]}
   );
   gpc1_1 gpc5490 (
      {stage0_59[416]},
      {stage1_59[198]}
   );
   gpc1_1 gpc5491 (
      {stage0_59[417]},
      {stage1_59[199]}
   );
   gpc1_1 gpc5492 (
      {stage0_59[418]},
      {stage1_59[200]}
   );
   gpc1_1 gpc5493 (
      {stage0_59[419]},
      {stage1_59[201]}
   );
   gpc1_1 gpc5494 (
      {stage0_59[420]},
      {stage1_59[202]}
   );
   gpc1_1 gpc5495 (
      {stage0_59[421]},
      {stage1_59[203]}
   );
   gpc1_1 gpc5496 (
      {stage0_59[422]},
      {stage1_59[204]}
   );
   gpc1_1 gpc5497 (
      {stage0_59[423]},
      {stage1_59[205]}
   );
   gpc1_1 gpc5498 (
      {stage0_59[424]},
      {stage1_59[206]}
   );
   gpc1_1 gpc5499 (
      {stage0_59[425]},
      {stage1_59[207]}
   );
   gpc1_1 gpc5500 (
      {stage0_59[426]},
      {stage1_59[208]}
   );
   gpc1_1 gpc5501 (
      {stage0_59[427]},
      {stage1_59[209]}
   );
   gpc1_1 gpc5502 (
      {stage0_59[428]},
      {stage1_59[210]}
   );
   gpc1_1 gpc5503 (
      {stage0_59[429]},
      {stage1_59[211]}
   );
   gpc1_1 gpc5504 (
      {stage0_59[430]},
      {stage1_59[212]}
   );
   gpc1_1 gpc5505 (
      {stage0_59[431]},
      {stage1_59[213]}
   );
   gpc1_1 gpc5506 (
      {stage0_59[432]},
      {stage1_59[214]}
   );
   gpc1_1 gpc5507 (
      {stage0_59[433]},
      {stage1_59[215]}
   );
   gpc1_1 gpc5508 (
      {stage0_59[434]},
      {stage1_59[216]}
   );
   gpc1_1 gpc5509 (
      {stage0_59[435]},
      {stage1_59[217]}
   );
   gpc1_1 gpc5510 (
      {stage0_59[436]},
      {stage1_59[218]}
   );
   gpc1_1 gpc5511 (
      {stage0_59[437]},
      {stage1_59[219]}
   );
   gpc1_1 gpc5512 (
      {stage0_59[438]},
      {stage1_59[220]}
   );
   gpc1_1 gpc5513 (
      {stage0_59[439]},
      {stage1_59[221]}
   );
   gpc1_1 gpc5514 (
      {stage0_59[440]},
      {stage1_59[222]}
   );
   gpc1_1 gpc5515 (
      {stage0_59[441]},
      {stage1_59[223]}
   );
   gpc1_1 gpc5516 (
      {stage0_59[442]},
      {stage1_59[224]}
   );
   gpc1_1 gpc5517 (
      {stage0_59[443]},
      {stage1_59[225]}
   );
   gpc1_1 gpc5518 (
      {stage0_59[444]},
      {stage1_59[226]}
   );
   gpc1_1 gpc5519 (
      {stage0_59[445]},
      {stage1_59[227]}
   );
   gpc1_1 gpc5520 (
      {stage0_59[446]},
      {stage1_59[228]}
   );
   gpc1_1 gpc5521 (
      {stage0_59[447]},
      {stage1_59[229]}
   );
   gpc1_1 gpc5522 (
      {stage0_59[448]},
      {stage1_59[230]}
   );
   gpc1_1 gpc5523 (
      {stage0_59[449]},
      {stage1_59[231]}
   );
   gpc1_1 gpc5524 (
      {stage0_59[450]},
      {stage1_59[232]}
   );
   gpc1_1 gpc5525 (
      {stage0_59[451]},
      {stage1_59[233]}
   );
   gpc1_1 gpc5526 (
      {stage0_59[452]},
      {stage1_59[234]}
   );
   gpc1_1 gpc5527 (
      {stage0_59[453]},
      {stage1_59[235]}
   );
   gpc1_1 gpc5528 (
      {stage0_59[454]},
      {stage1_59[236]}
   );
   gpc1_1 gpc5529 (
      {stage0_59[455]},
      {stage1_59[237]}
   );
   gpc1_1 gpc5530 (
      {stage0_59[456]},
      {stage1_59[238]}
   );
   gpc1_1 gpc5531 (
      {stage0_59[457]},
      {stage1_59[239]}
   );
   gpc1_1 gpc5532 (
      {stage0_59[458]},
      {stage1_59[240]}
   );
   gpc1_1 gpc5533 (
      {stage0_59[459]},
      {stage1_59[241]}
   );
   gpc1_1 gpc5534 (
      {stage0_59[460]},
      {stage1_59[242]}
   );
   gpc1_1 gpc5535 (
      {stage0_59[461]},
      {stage1_59[243]}
   );
   gpc1_1 gpc5536 (
      {stage0_59[462]},
      {stage1_59[244]}
   );
   gpc1_1 gpc5537 (
      {stage0_59[463]},
      {stage1_59[245]}
   );
   gpc1_1 gpc5538 (
      {stage0_59[464]},
      {stage1_59[246]}
   );
   gpc1_1 gpc5539 (
      {stage0_59[465]},
      {stage1_59[247]}
   );
   gpc1_1 gpc5540 (
      {stage0_59[466]},
      {stage1_59[248]}
   );
   gpc1_1 gpc5541 (
      {stage0_59[467]},
      {stage1_59[249]}
   );
   gpc1_1 gpc5542 (
      {stage0_59[468]},
      {stage1_59[250]}
   );
   gpc1_1 gpc5543 (
      {stage0_59[469]},
      {stage1_59[251]}
   );
   gpc1_1 gpc5544 (
      {stage0_59[470]},
      {stage1_59[252]}
   );
   gpc1_1 gpc5545 (
      {stage0_59[471]},
      {stage1_59[253]}
   );
   gpc1_1 gpc5546 (
      {stage0_59[472]},
      {stage1_59[254]}
   );
   gpc1_1 gpc5547 (
      {stage0_59[473]},
      {stage1_59[255]}
   );
   gpc1_1 gpc5548 (
      {stage0_59[474]},
      {stage1_59[256]}
   );
   gpc1_1 gpc5549 (
      {stage0_59[475]},
      {stage1_59[257]}
   );
   gpc1_1 gpc5550 (
      {stage0_59[476]},
      {stage1_59[258]}
   );
   gpc1_1 gpc5551 (
      {stage0_59[477]},
      {stage1_59[259]}
   );
   gpc1_1 gpc5552 (
      {stage0_59[478]},
      {stage1_59[260]}
   );
   gpc1_1 gpc5553 (
      {stage0_59[479]},
      {stage1_59[261]}
   );
   gpc1_1 gpc5554 (
      {stage0_59[480]},
      {stage1_59[262]}
   );
   gpc1_1 gpc5555 (
      {stage0_59[481]},
      {stage1_59[263]}
   );
   gpc1_1 gpc5556 (
      {stage0_59[482]},
      {stage1_59[264]}
   );
   gpc1_1 gpc5557 (
      {stage0_59[483]},
      {stage1_59[265]}
   );
   gpc1_1 gpc5558 (
      {stage0_59[484]},
      {stage1_59[266]}
   );
   gpc1_1 gpc5559 (
      {stage0_59[485]},
      {stage1_59[267]}
   );
   gpc1_1 gpc5560 (
      {stage0_59[486]},
      {stage1_59[268]}
   );
   gpc1_1 gpc5561 (
      {stage0_59[487]},
      {stage1_59[269]}
   );
   gpc1_1 gpc5562 (
      {stage0_59[488]},
      {stage1_59[270]}
   );
   gpc1_1 gpc5563 (
      {stage0_59[489]},
      {stage1_59[271]}
   );
   gpc1_1 gpc5564 (
      {stage0_59[490]},
      {stage1_59[272]}
   );
   gpc1_1 gpc5565 (
      {stage0_59[491]},
      {stage1_59[273]}
   );
   gpc1_1 gpc5566 (
      {stage0_59[492]},
      {stage1_59[274]}
   );
   gpc1_1 gpc5567 (
      {stage0_59[493]},
      {stage1_59[275]}
   );
   gpc1_1 gpc5568 (
      {stage0_59[494]},
      {stage1_59[276]}
   );
   gpc1_1 gpc5569 (
      {stage0_59[495]},
      {stage1_59[277]}
   );
   gpc1_1 gpc5570 (
      {stage0_59[496]},
      {stage1_59[278]}
   );
   gpc1_1 gpc5571 (
      {stage0_59[497]},
      {stage1_59[279]}
   );
   gpc1_1 gpc5572 (
      {stage0_59[498]},
      {stage1_59[280]}
   );
   gpc1_1 gpc5573 (
      {stage0_59[499]},
      {stage1_59[281]}
   );
   gpc1_1 gpc5574 (
      {stage0_59[500]},
      {stage1_59[282]}
   );
   gpc1_1 gpc5575 (
      {stage0_59[501]},
      {stage1_59[283]}
   );
   gpc1_1 gpc5576 (
      {stage0_59[502]},
      {stage1_59[284]}
   );
   gpc1_1 gpc5577 (
      {stage0_59[503]},
      {stage1_59[285]}
   );
   gpc1_1 gpc5578 (
      {stage0_59[504]},
      {stage1_59[286]}
   );
   gpc1_1 gpc5579 (
      {stage0_59[505]},
      {stage1_59[287]}
   );
   gpc1_1 gpc5580 (
      {stage0_59[506]},
      {stage1_59[288]}
   );
   gpc1_1 gpc5581 (
      {stage0_59[507]},
      {stage1_59[289]}
   );
   gpc1_1 gpc5582 (
      {stage0_59[508]},
      {stage1_59[290]}
   );
   gpc1_1 gpc5583 (
      {stage0_59[509]},
      {stage1_59[291]}
   );
   gpc1_1 gpc5584 (
      {stage0_59[510]},
      {stage1_59[292]}
   );
   gpc1_1 gpc5585 (
      {stage0_59[511]},
      {stage1_59[293]}
   );
   gpc1_1 gpc5586 (
      {stage0_60[502]},
      {stage1_60[190]}
   );
   gpc1_1 gpc5587 (
      {stage0_60[503]},
      {stage1_60[191]}
   );
   gpc1_1 gpc5588 (
      {stage0_60[504]},
      {stage1_60[192]}
   );
   gpc1_1 gpc5589 (
      {stage0_60[505]},
      {stage1_60[193]}
   );
   gpc1_1 gpc5590 (
      {stage0_60[506]},
      {stage1_60[194]}
   );
   gpc1_1 gpc5591 (
      {stage0_60[507]},
      {stage1_60[195]}
   );
   gpc1_1 gpc5592 (
      {stage0_60[508]},
      {stage1_60[196]}
   );
   gpc1_1 gpc5593 (
      {stage0_60[509]},
      {stage1_60[197]}
   );
   gpc1_1 gpc5594 (
      {stage0_60[510]},
      {stage1_60[198]}
   );
   gpc1_1 gpc5595 (
      {stage0_60[511]},
      {stage1_60[199]}
   );
   gpc1_1 gpc5596 (
      {stage0_62[330]},
      {stage1_62[191]}
   );
   gpc1_1 gpc5597 (
      {stage0_62[331]},
      {stage1_62[192]}
   );
   gpc1_1 gpc5598 (
      {stage0_62[332]},
      {stage1_62[193]}
   );
   gpc1_1 gpc5599 (
      {stage0_62[333]},
      {stage1_62[194]}
   );
   gpc1_1 gpc5600 (
      {stage0_62[334]},
      {stage1_62[195]}
   );
   gpc1_1 gpc5601 (
      {stage0_62[335]},
      {stage1_62[196]}
   );
   gpc1_1 gpc5602 (
      {stage0_62[336]},
      {stage1_62[197]}
   );
   gpc1_1 gpc5603 (
      {stage0_62[337]},
      {stage1_62[198]}
   );
   gpc1_1 gpc5604 (
      {stage0_62[338]},
      {stage1_62[199]}
   );
   gpc1_1 gpc5605 (
      {stage0_62[339]},
      {stage1_62[200]}
   );
   gpc1_1 gpc5606 (
      {stage0_62[340]},
      {stage1_62[201]}
   );
   gpc1_1 gpc5607 (
      {stage0_62[341]},
      {stage1_62[202]}
   );
   gpc1_1 gpc5608 (
      {stage0_62[342]},
      {stage1_62[203]}
   );
   gpc1_1 gpc5609 (
      {stage0_62[343]},
      {stage1_62[204]}
   );
   gpc1_1 gpc5610 (
      {stage0_62[344]},
      {stage1_62[205]}
   );
   gpc1_1 gpc5611 (
      {stage0_62[345]},
      {stage1_62[206]}
   );
   gpc1_1 gpc5612 (
      {stage0_62[346]},
      {stage1_62[207]}
   );
   gpc1_1 gpc5613 (
      {stage0_62[347]},
      {stage1_62[208]}
   );
   gpc1_1 gpc5614 (
      {stage0_62[348]},
      {stage1_62[209]}
   );
   gpc1_1 gpc5615 (
      {stage0_62[349]},
      {stage1_62[210]}
   );
   gpc1_1 gpc5616 (
      {stage0_62[350]},
      {stage1_62[211]}
   );
   gpc1_1 gpc5617 (
      {stage0_62[351]},
      {stage1_62[212]}
   );
   gpc1_1 gpc5618 (
      {stage0_62[352]},
      {stage1_62[213]}
   );
   gpc1_1 gpc5619 (
      {stage0_62[353]},
      {stage1_62[214]}
   );
   gpc1_1 gpc5620 (
      {stage0_62[354]},
      {stage1_62[215]}
   );
   gpc1_1 gpc5621 (
      {stage0_62[355]},
      {stage1_62[216]}
   );
   gpc1_1 gpc5622 (
      {stage0_62[356]},
      {stage1_62[217]}
   );
   gpc1_1 gpc5623 (
      {stage0_62[357]},
      {stage1_62[218]}
   );
   gpc1_1 gpc5624 (
      {stage0_62[358]},
      {stage1_62[219]}
   );
   gpc1_1 gpc5625 (
      {stage0_62[359]},
      {stage1_62[220]}
   );
   gpc1_1 gpc5626 (
      {stage0_62[360]},
      {stage1_62[221]}
   );
   gpc1_1 gpc5627 (
      {stage0_62[361]},
      {stage1_62[222]}
   );
   gpc1_1 gpc5628 (
      {stage0_62[362]},
      {stage1_62[223]}
   );
   gpc1_1 gpc5629 (
      {stage0_62[363]},
      {stage1_62[224]}
   );
   gpc1_1 gpc5630 (
      {stage0_62[364]},
      {stage1_62[225]}
   );
   gpc1_1 gpc5631 (
      {stage0_62[365]},
      {stage1_62[226]}
   );
   gpc1_1 gpc5632 (
      {stage0_62[366]},
      {stage1_62[227]}
   );
   gpc1_1 gpc5633 (
      {stage0_62[367]},
      {stage1_62[228]}
   );
   gpc1_1 gpc5634 (
      {stage0_62[368]},
      {stage1_62[229]}
   );
   gpc1_1 gpc5635 (
      {stage0_62[369]},
      {stage1_62[230]}
   );
   gpc1_1 gpc5636 (
      {stage0_62[370]},
      {stage1_62[231]}
   );
   gpc1_1 gpc5637 (
      {stage0_62[371]},
      {stage1_62[232]}
   );
   gpc1_1 gpc5638 (
      {stage0_62[372]},
      {stage1_62[233]}
   );
   gpc1_1 gpc5639 (
      {stage0_62[373]},
      {stage1_62[234]}
   );
   gpc1_1 gpc5640 (
      {stage0_62[374]},
      {stage1_62[235]}
   );
   gpc1_1 gpc5641 (
      {stage0_62[375]},
      {stage1_62[236]}
   );
   gpc1_1 gpc5642 (
      {stage0_62[376]},
      {stage1_62[237]}
   );
   gpc1_1 gpc5643 (
      {stage0_62[377]},
      {stage1_62[238]}
   );
   gpc1_1 gpc5644 (
      {stage0_62[378]},
      {stage1_62[239]}
   );
   gpc1_1 gpc5645 (
      {stage0_62[379]},
      {stage1_62[240]}
   );
   gpc1_1 gpc5646 (
      {stage0_62[380]},
      {stage1_62[241]}
   );
   gpc1_1 gpc5647 (
      {stage0_62[381]},
      {stage1_62[242]}
   );
   gpc1_1 gpc5648 (
      {stage0_62[382]},
      {stage1_62[243]}
   );
   gpc1_1 gpc5649 (
      {stage0_62[383]},
      {stage1_62[244]}
   );
   gpc1_1 gpc5650 (
      {stage0_62[384]},
      {stage1_62[245]}
   );
   gpc1_1 gpc5651 (
      {stage0_62[385]},
      {stage1_62[246]}
   );
   gpc1_1 gpc5652 (
      {stage0_62[386]},
      {stage1_62[247]}
   );
   gpc1_1 gpc5653 (
      {stage0_62[387]},
      {stage1_62[248]}
   );
   gpc1_1 gpc5654 (
      {stage0_62[388]},
      {stage1_62[249]}
   );
   gpc1_1 gpc5655 (
      {stage0_62[389]},
      {stage1_62[250]}
   );
   gpc1_1 gpc5656 (
      {stage0_62[390]},
      {stage1_62[251]}
   );
   gpc1_1 gpc5657 (
      {stage0_62[391]},
      {stage1_62[252]}
   );
   gpc1_1 gpc5658 (
      {stage0_62[392]},
      {stage1_62[253]}
   );
   gpc1_1 gpc5659 (
      {stage0_62[393]},
      {stage1_62[254]}
   );
   gpc1_1 gpc5660 (
      {stage0_62[394]},
      {stage1_62[255]}
   );
   gpc1_1 gpc5661 (
      {stage0_62[395]},
      {stage1_62[256]}
   );
   gpc1_1 gpc5662 (
      {stage0_62[396]},
      {stage1_62[257]}
   );
   gpc1_1 gpc5663 (
      {stage0_62[397]},
      {stage1_62[258]}
   );
   gpc1_1 gpc5664 (
      {stage0_62[398]},
      {stage1_62[259]}
   );
   gpc1_1 gpc5665 (
      {stage0_62[399]},
      {stage1_62[260]}
   );
   gpc1_1 gpc5666 (
      {stage0_62[400]},
      {stage1_62[261]}
   );
   gpc1_1 gpc5667 (
      {stage0_62[401]},
      {stage1_62[262]}
   );
   gpc1_1 gpc5668 (
      {stage0_62[402]},
      {stage1_62[263]}
   );
   gpc1_1 gpc5669 (
      {stage0_62[403]},
      {stage1_62[264]}
   );
   gpc1_1 gpc5670 (
      {stage0_62[404]},
      {stage1_62[265]}
   );
   gpc1_1 gpc5671 (
      {stage0_62[405]},
      {stage1_62[266]}
   );
   gpc1_1 gpc5672 (
      {stage0_62[406]},
      {stage1_62[267]}
   );
   gpc1_1 gpc5673 (
      {stage0_62[407]},
      {stage1_62[268]}
   );
   gpc1_1 gpc5674 (
      {stage0_62[408]},
      {stage1_62[269]}
   );
   gpc1_1 gpc5675 (
      {stage0_62[409]},
      {stage1_62[270]}
   );
   gpc1_1 gpc5676 (
      {stage0_62[410]},
      {stage1_62[271]}
   );
   gpc1_1 gpc5677 (
      {stage0_62[411]},
      {stage1_62[272]}
   );
   gpc1_1 gpc5678 (
      {stage0_62[412]},
      {stage1_62[273]}
   );
   gpc1_1 gpc5679 (
      {stage0_62[413]},
      {stage1_62[274]}
   );
   gpc1_1 gpc5680 (
      {stage0_62[414]},
      {stage1_62[275]}
   );
   gpc1_1 gpc5681 (
      {stage0_62[415]},
      {stage1_62[276]}
   );
   gpc1_1 gpc5682 (
      {stage0_62[416]},
      {stage1_62[277]}
   );
   gpc1_1 gpc5683 (
      {stage0_62[417]},
      {stage1_62[278]}
   );
   gpc1_1 gpc5684 (
      {stage0_62[418]},
      {stage1_62[279]}
   );
   gpc1_1 gpc5685 (
      {stage0_62[419]},
      {stage1_62[280]}
   );
   gpc1_1 gpc5686 (
      {stage0_62[420]},
      {stage1_62[281]}
   );
   gpc1_1 gpc5687 (
      {stage0_62[421]},
      {stage1_62[282]}
   );
   gpc1_1 gpc5688 (
      {stage0_62[422]},
      {stage1_62[283]}
   );
   gpc1_1 gpc5689 (
      {stage0_62[423]},
      {stage1_62[284]}
   );
   gpc1_1 gpc5690 (
      {stage0_62[424]},
      {stage1_62[285]}
   );
   gpc1_1 gpc5691 (
      {stage0_62[425]},
      {stage1_62[286]}
   );
   gpc1_1 gpc5692 (
      {stage0_62[426]},
      {stage1_62[287]}
   );
   gpc1_1 gpc5693 (
      {stage0_62[427]},
      {stage1_62[288]}
   );
   gpc1_1 gpc5694 (
      {stage0_62[428]},
      {stage1_62[289]}
   );
   gpc1_1 gpc5695 (
      {stage0_62[429]},
      {stage1_62[290]}
   );
   gpc1_1 gpc5696 (
      {stage0_62[430]},
      {stage1_62[291]}
   );
   gpc1_1 gpc5697 (
      {stage0_62[431]},
      {stage1_62[292]}
   );
   gpc1_1 gpc5698 (
      {stage0_62[432]},
      {stage1_62[293]}
   );
   gpc1_1 gpc5699 (
      {stage0_62[433]},
      {stage1_62[294]}
   );
   gpc1_1 gpc5700 (
      {stage0_62[434]},
      {stage1_62[295]}
   );
   gpc1_1 gpc5701 (
      {stage0_62[435]},
      {stage1_62[296]}
   );
   gpc1_1 gpc5702 (
      {stage0_62[436]},
      {stage1_62[297]}
   );
   gpc1_1 gpc5703 (
      {stage0_62[437]},
      {stage1_62[298]}
   );
   gpc1_1 gpc5704 (
      {stage0_62[438]},
      {stage1_62[299]}
   );
   gpc1_1 gpc5705 (
      {stage0_62[439]},
      {stage1_62[300]}
   );
   gpc1_1 gpc5706 (
      {stage0_62[440]},
      {stage1_62[301]}
   );
   gpc1_1 gpc5707 (
      {stage0_62[441]},
      {stage1_62[302]}
   );
   gpc1_1 gpc5708 (
      {stage0_62[442]},
      {stage1_62[303]}
   );
   gpc1_1 gpc5709 (
      {stage0_62[443]},
      {stage1_62[304]}
   );
   gpc1_1 gpc5710 (
      {stage0_62[444]},
      {stage1_62[305]}
   );
   gpc1_1 gpc5711 (
      {stage0_62[445]},
      {stage1_62[306]}
   );
   gpc1_1 gpc5712 (
      {stage0_62[446]},
      {stage1_62[307]}
   );
   gpc1_1 gpc5713 (
      {stage0_62[447]},
      {stage1_62[308]}
   );
   gpc1_1 gpc5714 (
      {stage0_62[448]},
      {stage1_62[309]}
   );
   gpc1_1 gpc5715 (
      {stage0_62[449]},
      {stage1_62[310]}
   );
   gpc1_1 gpc5716 (
      {stage0_62[450]},
      {stage1_62[311]}
   );
   gpc1_1 gpc5717 (
      {stage0_62[451]},
      {stage1_62[312]}
   );
   gpc1_1 gpc5718 (
      {stage0_62[452]},
      {stage1_62[313]}
   );
   gpc1_1 gpc5719 (
      {stage0_62[453]},
      {stage1_62[314]}
   );
   gpc1_1 gpc5720 (
      {stage0_62[454]},
      {stage1_62[315]}
   );
   gpc1_1 gpc5721 (
      {stage0_62[455]},
      {stage1_62[316]}
   );
   gpc1_1 gpc5722 (
      {stage0_62[456]},
      {stage1_62[317]}
   );
   gpc1_1 gpc5723 (
      {stage0_62[457]},
      {stage1_62[318]}
   );
   gpc1_1 gpc5724 (
      {stage0_62[458]},
      {stage1_62[319]}
   );
   gpc1_1 gpc5725 (
      {stage0_62[459]},
      {stage1_62[320]}
   );
   gpc1_1 gpc5726 (
      {stage0_62[460]},
      {stage1_62[321]}
   );
   gpc1_1 gpc5727 (
      {stage0_62[461]},
      {stage1_62[322]}
   );
   gpc1_1 gpc5728 (
      {stage0_62[462]},
      {stage1_62[323]}
   );
   gpc1_1 gpc5729 (
      {stage0_62[463]},
      {stage1_62[324]}
   );
   gpc1_1 gpc5730 (
      {stage0_62[464]},
      {stage1_62[325]}
   );
   gpc1_1 gpc5731 (
      {stage0_62[465]},
      {stage1_62[326]}
   );
   gpc1_1 gpc5732 (
      {stage0_62[466]},
      {stage1_62[327]}
   );
   gpc1_1 gpc5733 (
      {stage0_62[467]},
      {stage1_62[328]}
   );
   gpc1_1 gpc5734 (
      {stage0_62[468]},
      {stage1_62[329]}
   );
   gpc1_1 gpc5735 (
      {stage0_62[469]},
      {stage1_62[330]}
   );
   gpc1_1 gpc5736 (
      {stage0_62[470]},
      {stage1_62[331]}
   );
   gpc1_1 gpc5737 (
      {stage0_62[471]},
      {stage1_62[332]}
   );
   gpc1_1 gpc5738 (
      {stage0_62[472]},
      {stage1_62[333]}
   );
   gpc1_1 gpc5739 (
      {stage0_62[473]},
      {stage1_62[334]}
   );
   gpc1_1 gpc5740 (
      {stage0_62[474]},
      {stage1_62[335]}
   );
   gpc1_1 gpc5741 (
      {stage0_62[475]},
      {stage1_62[336]}
   );
   gpc1_1 gpc5742 (
      {stage0_62[476]},
      {stage1_62[337]}
   );
   gpc1_1 gpc5743 (
      {stage0_62[477]},
      {stage1_62[338]}
   );
   gpc1_1 gpc5744 (
      {stage0_62[478]},
      {stage1_62[339]}
   );
   gpc1_1 gpc5745 (
      {stage0_62[479]},
      {stage1_62[340]}
   );
   gpc1_1 gpc5746 (
      {stage0_62[480]},
      {stage1_62[341]}
   );
   gpc1_1 gpc5747 (
      {stage0_62[481]},
      {stage1_62[342]}
   );
   gpc1_1 gpc5748 (
      {stage0_62[482]},
      {stage1_62[343]}
   );
   gpc1_1 gpc5749 (
      {stage0_62[483]},
      {stage1_62[344]}
   );
   gpc1_1 gpc5750 (
      {stage0_62[484]},
      {stage1_62[345]}
   );
   gpc1_1 gpc5751 (
      {stage0_62[485]},
      {stage1_62[346]}
   );
   gpc1_1 gpc5752 (
      {stage0_62[486]},
      {stage1_62[347]}
   );
   gpc1_1 gpc5753 (
      {stage0_62[487]},
      {stage1_62[348]}
   );
   gpc1_1 gpc5754 (
      {stage0_62[488]},
      {stage1_62[349]}
   );
   gpc1_1 gpc5755 (
      {stage0_62[489]},
      {stage1_62[350]}
   );
   gpc1_1 gpc5756 (
      {stage0_62[490]},
      {stage1_62[351]}
   );
   gpc1_1 gpc5757 (
      {stage0_62[491]},
      {stage1_62[352]}
   );
   gpc1_1 gpc5758 (
      {stage0_62[492]},
      {stage1_62[353]}
   );
   gpc1_1 gpc5759 (
      {stage0_62[493]},
      {stage1_62[354]}
   );
   gpc1_1 gpc5760 (
      {stage0_62[494]},
      {stage1_62[355]}
   );
   gpc1_1 gpc5761 (
      {stage0_62[495]},
      {stage1_62[356]}
   );
   gpc1_1 gpc5762 (
      {stage0_62[496]},
      {stage1_62[357]}
   );
   gpc1_1 gpc5763 (
      {stage0_62[497]},
      {stage1_62[358]}
   );
   gpc1_1 gpc5764 (
      {stage0_62[498]},
      {stage1_62[359]}
   );
   gpc1_1 gpc5765 (
      {stage0_62[499]},
      {stage1_62[360]}
   );
   gpc1_1 gpc5766 (
      {stage0_62[500]},
      {stage1_62[361]}
   );
   gpc1_1 gpc5767 (
      {stage0_62[501]},
      {stage1_62[362]}
   );
   gpc1_1 gpc5768 (
      {stage0_62[502]},
      {stage1_62[363]}
   );
   gpc1_1 gpc5769 (
      {stage0_62[503]},
      {stage1_62[364]}
   );
   gpc1_1 gpc5770 (
      {stage0_62[504]},
      {stage1_62[365]}
   );
   gpc1_1 gpc5771 (
      {stage0_62[505]},
      {stage1_62[366]}
   );
   gpc1_1 gpc5772 (
      {stage0_62[506]},
      {stage1_62[367]}
   );
   gpc1_1 gpc5773 (
      {stage0_62[507]},
      {stage1_62[368]}
   );
   gpc1_1 gpc5774 (
      {stage0_62[508]},
      {stage1_62[369]}
   );
   gpc1_1 gpc5775 (
      {stage0_62[509]},
      {stage1_62[370]}
   );
   gpc1_1 gpc5776 (
      {stage0_62[510]},
      {stage1_62[371]}
   );
   gpc1_1 gpc5777 (
      {stage0_62[511]},
      {stage1_62[372]}
   );
   gpc1_1 gpc5778 (
      {stage0_63[342]},
      {stage1_63[125]}
   );
   gpc1_1 gpc5779 (
      {stage0_63[343]},
      {stage1_63[126]}
   );
   gpc1_1 gpc5780 (
      {stage0_63[344]},
      {stage1_63[127]}
   );
   gpc1_1 gpc5781 (
      {stage0_63[345]},
      {stage1_63[128]}
   );
   gpc1_1 gpc5782 (
      {stage0_63[346]},
      {stage1_63[129]}
   );
   gpc1_1 gpc5783 (
      {stage0_63[347]},
      {stage1_63[130]}
   );
   gpc1_1 gpc5784 (
      {stage0_63[348]},
      {stage1_63[131]}
   );
   gpc1_1 gpc5785 (
      {stage0_63[349]},
      {stage1_63[132]}
   );
   gpc1_1 gpc5786 (
      {stage0_63[350]},
      {stage1_63[133]}
   );
   gpc1_1 gpc5787 (
      {stage0_63[351]},
      {stage1_63[134]}
   );
   gpc1_1 gpc5788 (
      {stage0_63[352]},
      {stage1_63[135]}
   );
   gpc1_1 gpc5789 (
      {stage0_63[353]},
      {stage1_63[136]}
   );
   gpc1_1 gpc5790 (
      {stage0_63[354]},
      {stage1_63[137]}
   );
   gpc1_1 gpc5791 (
      {stage0_63[355]},
      {stage1_63[138]}
   );
   gpc1_1 gpc5792 (
      {stage0_63[356]},
      {stage1_63[139]}
   );
   gpc1_1 gpc5793 (
      {stage0_63[357]},
      {stage1_63[140]}
   );
   gpc1_1 gpc5794 (
      {stage0_63[358]},
      {stage1_63[141]}
   );
   gpc1_1 gpc5795 (
      {stage0_63[359]},
      {stage1_63[142]}
   );
   gpc1_1 gpc5796 (
      {stage0_63[360]},
      {stage1_63[143]}
   );
   gpc1_1 gpc5797 (
      {stage0_63[361]},
      {stage1_63[144]}
   );
   gpc1_1 gpc5798 (
      {stage0_63[362]},
      {stage1_63[145]}
   );
   gpc1_1 gpc5799 (
      {stage0_63[363]},
      {stage1_63[146]}
   );
   gpc1_1 gpc5800 (
      {stage0_63[364]},
      {stage1_63[147]}
   );
   gpc1_1 gpc5801 (
      {stage0_63[365]},
      {stage1_63[148]}
   );
   gpc1_1 gpc5802 (
      {stage0_63[366]},
      {stage1_63[149]}
   );
   gpc1_1 gpc5803 (
      {stage0_63[367]},
      {stage1_63[150]}
   );
   gpc1_1 gpc5804 (
      {stage0_63[368]},
      {stage1_63[151]}
   );
   gpc1_1 gpc5805 (
      {stage0_63[369]},
      {stage1_63[152]}
   );
   gpc1_1 gpc5806 (
      {stage0_63[370]},
      {stage1_63[153]}
   );
   gpc1_1 gpc5807 (
      {stage0_63[371]},
      {stage1_63[154]}
   );
   gpc1_1 gpc5808 (
      {stage0_63[372]},
      {stage1_63[155]}
   );
   gpc1_1 gpc5809 (
      {stage0_63[373]},
      {stage1_63[156]}
   );
   gpc1_1 gpc5810 (
      {stage0_63[374]},
      {stage1_63[157]}
   );
   gpc1_1 gpc5811 (
      {stage0_63[375]},
      {stage1_63[158]}
   );
   gpc1_1 gpc5812 (
      {stage0_63[376]},
      {stage1_63[159]}
   );
   gpc1_1 gpc5813 (
      {stage0_63[377]},
      {stage1_63[160]}
   );
   gpc1_1 gpc5814 (
      {stage0_63[378]},
      {stage1_63[161]}
   );
   gpc1_1 gpc5815 (
      {stage0_63[379]},
      {stage1_63[162]}
   );
   gpc1_1 gpc5816 (
      {stage0_63[380]},
      {stage1_63[163]}
   );
   gpc1_1 gpc5817 (
      {stage0_63[381]},
      {stage1_63[164]}
   );
   gpc1_1 gpc5818 (
      {stage0_63[382]},
      {stage1_63[165]}
   );
   gpc1_1 gpc5819 (
      {stage0_63[383]},
      {stage1_63[166]}
   );
   gpc1_1 gpc5820 (
      {stage0_63[384]},
      {stage1_63[167]}
   );
   gpc1_1 gpc5821 (
      {stage0_63[385]},
      {stage1_63[168]}
   );
   gpc1_1 gpc5822 (
      {stage0_63[386]},
      {stage1_63[169]}
   );
   gpc1_1 gpc5823 (
      {stage0_63[387]},
      {stage1_63[170]}
   );
   gpc1_1 gpc5824 (
      {stage0_63[388]},
      {stage1_63[171]}
   );
   gpc1_1 gpc5825 (
      {stage0_63[389]},
      {stage1_63[172]}
   );
   gpc1_1 gpc5826 (
      {stage0_63[390]},
      {stage1_63[173]}
   );
   gpc1_1 gpc5827 (
      {stage0_63[391]},
      {stage1_63[174]}
   );
   gpc1_1 gpc5828 (
      {stage0_63[392]},
      {stage1_63[175]}
   );
   gpc1_1 gpc5829 (
      {stage0_63[393]},
      {stage1_63[176]}
   );
   gpc1_1 gpc5830 (
      {stage0_63[394]},
      {stage1_63[177]}
   );
   gpc1_1 gpc5831 (
      {stage0_63[395]},
      {stage1_63[178]}
   );
   gpc1_1 gpc5832 (
      {stage0_63[396]},
      {stage1_63[179]}
   );
   gpc1_1 gpc5833 (
      {stage0_63[397]},
      {stage1_63[180]}
   );
   gpc1_1 gpc5834 (
      {stage0_63[398]},
      {stage1_63[181]}
   );
   gpc1_1 gpc5835 (
      {stage0_63[399]},
      {stage1_63[182]}
   );
   gpc1_1 gpc5836 (
      {stage0_63[400]},
      {stage1_63[183]}
   );
   gpc1_1 gpc5837 (
      {stage0_63[401]},
      {stage1_63[184]}
   );
   gpc1_1 gpc5838 (
      {stage0_63[402]},
      {stage1_63[185]}
   );
   gpc1_1 gpc5839 (
      {stage0_63[403]},
      {stage1_63[186]}
   );
   gpc1_1 gpc5840 (
      {stage0_63[404]},
      {stage1_63[187]}
   );
   gpc1_1 gpc5841 (
      {stage0_63[405]},
      {stage1_63[188]}
   );
   gpc1_1 gpc5842 (
      {stage0_63[406]},
      {stage1_63[189]}
   );
   gpc1_1 gpc5843 (
      {stage0_63[407]},
      {stage1_63[190]}
   );
   gpc1_1 gpc5844 (
      {stage0_63[408]},
      {stage1_63[191]}
   );
   gpc1_1 gpc5845 (
      {stage0_63[409]},
      {stage1_63[192]}
   );
   gpc1_1 gpc5846 (
      {stage0_63[410]},
      {stage1_63[193]}
   );
   gpc1_1 gpc5847 (
      {stage0_63[411]},
      {stage1_63[194]}
   );
   gpc1_1 gpc5848 (
      {stage0_63[412]},
      {stage1_63[195]}
   );
   gpc1_1 gpc5849 (
      {stage0_63[413]},
      {stage1_63[196]}
   );
   gpc1_1 gpc5850 (
      {stage0_63[414]},
      {stage1_63[197]}
   );
   gpc1_1 gpc5851 (
      {stage0_63[415]},
      {stage1_63[198]}
   );
   gpc1_1 gpc5852 (
      {stage0_63[416]},
      {stage1_63[199]}
   );
   gpc1_1 gpc5853 (
      {stage0_63[417]},
      {stage1_63[200]}
   );
   gpc1_1 gpc5854 (
      {stage0_63[418]},
      {stage1_63[201]}
   );
   gpc1_1 gpc5855 (
      {stage0_63[419]},
      {stage1_63[202]}
   );
   gpc1_1 gpc5856 (
      {stage0_63[420]},
      {stage1_63[203]}
   );
   gpc1_1 gpc5857 (
      {stage0_63[421]},
      {stage1_63[204]}
   );
   gpc1_1 gpc5858 (
      {stage0_63[422]},
      {stage1_63[205]}
   );
   gpc1_1 gpc5859 (
      {stage0_63[423]},
      {stage1_63[206]}
   );
   gpc1_1 gpc5860 (
      {stage0_63[424]},
      {stage1_63[207]}
   );
   gpc1_1 gpc5861 (
      {stage0_63[425]},
      {stage1_63[208]}
   );
   gpc1_1 gpc5862 (
      {stage0_63[426]},
      {stage1_63[209]}
   );
   gpc1_1 gpc5863 (
      {stage0_63[427]},
      {stage1_63[210]}
   );
   gpc1_1 gpc5864 (
      {stage0_63[428]},
      {stage1_63[211]}
   );
   gpc1_1 gpc5865 (
      {stage0_63[429]},
      {stage1_63[212]}
   );
   gpc1_1 gpc5866 (
      {stage0_63[430]},
      {stage1_63[213]}
   );
   gpc1_1 gpc5867 (
      {stage0_63[431]},
      {stage1_63[214]}
   );
   gpc1_1 gpc5868 (
      {stage0_63[432]},
      {stage1_63[215]}
   );
   gpc1_1 gpc5869 (
      {stage0_63[433]},
      {stage1_63[216]}
   );
   gpc1_1 gpc5870 (
      {stage0_63[434]},
      {stage1_63[217]}
   );
   gpc1_1 gpc5871 (
      {stage0_63[435]},
      {stage1_63[218]}
   );
   gpc1_1 gpc5872 (
      {stage0_63[436]},
      {stage1_63[219]}
   );
   gpc1_1 gpc5873 (
      {stage0_63[437]},
      {stage1_63[220]}
   );
   gpc1_1 gpc5874 (
      {stage0_63[438]},
      {stage1_63[221]}
   );
   gpc1_1 gpc5875 (
      {stage0_63[439]},
      {stage1_63[222]}
   );
   gpc1_1 gpc5876 (
      {stage0_63[440]},
      {stage1_63[223]}
   );
   gpc1_1 gpc5877 (
      {stage0_63[441]},
      {stage1_63[224]}
   );
   gpc1_1 gpc5878 (
      {stage0_63[442]},
      {stage1_63[225]}
   );
   gpc1_1 gpc5879 (
      {stage0_63[443]},
      {stage1_63[226]}
   );
   gpc1_1 gpc5880 (
      {stage0_63[444]},
      {stage1_63[227]}
   );
   gpc1_1 gpc5881 (
      {stage0_63[445]},
      {stage1_63[228]}
   );
   gpc1_1 gpc5882 (
      {stage0_63[446]},
      {stage1_63[229]}
   );
   gpc1_1 gpc5883 (
      {stage0_63[447]},
      {stage1_63[230]}
   );
   gpc1_1 gpc5884 (
      {stage0_63[448]},
      {stage1_63[231]}
   );
   gpc1_1 gpc5885 (
      {stage0_63[449]},
      {stage1_63[232]}
   );
   gpc1_1 gpc5886 (
      {stage0_63[450]},
      {stage1_63[233]}
   );
   gpc1_1 gpc5887 (
      {stage0_63[451]},
      {stage1_63[234]}
   );
   gpc1_1 gpc5888 (
      {stage0_63[452]},
      {stage1_63[235]}
   );
   gpc1_1 gpc5889 (
      {stage0_63[453]},
      {stage1_63[236]}
   );
   gpc1_1 gpc5890 (
      {stage0_63[454]},
      {stage1_63[237]}
   );
   gpc1_1 gpc5891 (
      {stage0_63[455]},
      {stage1_63[238]}
   );
   gpc1_1 gpc5892 (
      {stage0_63[456]},
      {stage1_63[239]}
   );
   gpc1_1 gpc5893 (
      {stage0_63[457]},
      {stage1_63[240]}
   );
   gpc1_1 gpc5894 (
      {stage0_63[458]},
      {stage1_63[241]}
   );
   gpc1_1 gpc5895 (
      {stage0_63[459]},
      {stage1_63[242]}
   );
   gpc1_1 gpc5896 (
      {stage0_63[460]},
      {stage1_63[243]}
   );
   gpc1_1 gpc5897 (
      {stage0_63[461]},
      {stage1_63[244]}
   );
   gpc1_1 gpc5898 (
      {stage0_63[462]},
      {stage1_63[245]}
   );
   gpc1_1 gpc5899 (
      {stage0_63[463]},
      {stage1_63[246]}
   );
   gpc1_1 gpc5900 (
      {stage0_63[464]},
      {stage1_63[247]}
   );
   gpc1_1 gpc5901 (
      {stage0_63[465]},
      {stage1_63[248]}
   );
   gpc1_1 gpc5902 (
      {stage0_63[466]},
      {stage1_63[249]}
   );
   gpc1_1 gpc5903 (
      {stage0_63[467]},
      {stage1_63[250]}
   );
   gpc1_1 gpc5904 (
      {stage0_63[468]},
      {stage1_63[251]}
   );
   gpc1_1 gpc5905 (
      {stage0_63[469]},
      {stage1_63[252]}
   );
   gpc1_1 gpc5906 (
      {stage0_63[470]},
      {stage1_63[253]}
   );
   gpc1_1 gpc5907 (
      {stage0_63[471]},
      {stage1_63[254]}
   );
   gpc1_1 gpc5908 (
      {stage0_63[472]},
      {stage1_63[255]}
   );
   gpc1_1 gpc5909 (
      {stage0_63[473]},
      {stage1_63[256]}
   );
   gpc1_1 gpc5910 (
      {stage0_63[474]},
      {stage1_63[257]}
   );
   gpc1_1 gpc5911 (
      {stage0_63[475]},
      {stage1_63[258]}
   );
   gpc1_1 gpc5912 (
      {stage0_63[476]},
      {stage1_63[259]}
   );
   gpc1_1 gpc5913 (
      {stage0_63[477]},
      {stage1_63[260]}
   );
   gpc1_1 gpc5914 (
      {stage0_63[478]},
      {stage1_63[261]}
   );
   gpc1_1 gpc5915 (
      {stage0_63[479]},
      {stage1_63[262]}
   );
   gpc1_1 gpc5916 (
      {stage0_63[480]},
      {stage1_63[263]}
   );
   gpc1_1 gpc5917 (
      {stage0_63[481]},
      {stage1_63[264]}
   );
   gpc1_1 gpc5918 (
      {stage0_63[482]},
      {stage1_63[265]}
   );
   gpc1_1 gpc5919 (
      {stage0_63[483]},
      {stage1_63[266]}
   );
   gpc1_1 gpc5920 (
      {stage0_63[484]},
      {stage1_63[267]}
   );
   gpc1_1 gpc5921 (
      {stage0_63[485]},
      {stage1_63[268]}
   );
   gpc1_1 gpc5922 (
      {stage0_63[486]},
      {stage1_63[269]}
   );
   gpc1_1 gpc5923 (
      {stage0_63[487]},
      {stage1_63[270]}
   );
   gpc1_1 gpc5924 (
      {stage0_63[488]},
      {stage1_63[271]}
   );
   gpc1_1 gpc5925 (
      {stage0_63[489]},
      {stage1_63[272]}
   );
   gpc1_1 gpc5926 (
      {stage0_63[490]},
      {stage1_63[273]}
   );
   gpc1_1 gpc5927 (
      {stage0_63[491]},
      {stage1_63[274]}
   );
   gpc1_1 gpc5928 (
      {stage0_63[492]},
      {stage1_63[275]}
   );
   gpc1_1 gpc5929 (
      {stage0_63[493]},
      {stage1_63[276]}
   );
   gpc1_1 gpc5930 (
      {stage0_63[494]},
      {stage1_63[277]}
   );
   gpc1_1 gpc5931 (
      {stage0_63[495]},
      {stage1_63[278]}
   );
   gpc1_1 gpc5932 (
      {stage0_63[496]},
      {stage1_63[279]}
   );
   gpc1_1 gpc5933 (
      {stage0_63[497]},
      {stage1_63[280]}
   );
   gpc1_1 gpc5934 (
      {stage0_63[498]},
      {stage1_63[281]}
   );
   gpc1_1 gpc5935 (
      {stage0_63[499]},
      {stage1_63[282]}
   );
   gpc1_1 gpc5936 (
      {stage0_63[500]},
      {stage1_63[283]}
   );
   gpc1_1 gpc5937 (
      {stage0_63[501]},
      {stage1_63[284]}
   );
   gpc1_1 gpc5938 (
      {stage0_63[502]},
      {stage1_63[285]}
   );
   gpc1_1 gpc5939 (
      {stage0_63[503]},
      {stage1_63[286]}
   );
   gpc1_1 gpc5940 (
      {stage0_63[504]},
      {stage1_63[287]}
   );
   gpc1_1 gpc5941 (
      {stage0_63[505]},
      {stage1_63[288]}
   );
   gpc1_1 gpc5942 (
      {stage0_63[506]},
      {stage1_63[289]}
   );
   gpc1_1 gpc5943 (
      {stage0_63[507]},
      {stage1_63[290]}
   );
   gpc1_1 gpc5944 (
      {stage0_63[508]},
      {stage1_63[291]}
   );
   gpc1_1 gpc5945 (
      {stage0_63[509]},
      {stage1_63[292]}
   );
   gpc1_1 gpc5946 (
      {stage0_63[510]},
      {stage1_63[293]}
   );
   gpc1_1 gpc5947 (
      {stage0_63[511]},
      {stage1_63[294]}
   );
   gpc1163_5 gpc5948 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc5949 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc5950 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc5951 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc5952 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc5953 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc5954 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc5955 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc5956 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc5957 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc5958 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc5959 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc5960 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc5961 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc5962 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc5963 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc5964 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc5965 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc5966 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc5967 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc5968 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc5969 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc5970 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc5971 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc5972 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc615_5 gpc5973 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106]},
      {stage1_1[96]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc615_5 gpc5974 (
      {stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111]},
      {stage1_1[97]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc5975 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[0],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc5976 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[1],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc5977 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[2],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc5978 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[3],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc5979 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[4],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc5980 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[5],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc5981 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[6],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc5982 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage2_5[7],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc5983 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69]},
      {stage2_5[8],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc5984 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage2_5[9],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc5985 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage2_5[10],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc5986 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], 1'b0},
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87]},
      {stage2_5[11],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc5987 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[12],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc5988 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[13],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc5989 (
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[14],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc5990 (
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[15],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc5991 (
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[16],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc606_5 gpc5992 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[17],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc606_5 gpc5993 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[18],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc606_5 gpc5994 (
      {stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[19],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc5995 (
      {stage1_2[130], stage1_2[131], stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[20],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc5996 (
      {stage1_2[136], stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[21],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc606_5 gpc5997 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[22],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc606_5 gpc5998 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152], stage1_2[153]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[23],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc606_5 gpc5999 (
      {stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157], stage1_2[158], stage1_2[159]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[24],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc606_5 gpc6000 (
      {stage1_2[160], stage1_2[161], stage1_2[162], stage1_2[163], stage1_2[164], stage1_2[165]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[25],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc606_5 gpc6001 (
      {stage1_2[166], stage1_2[167], stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[26],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc606_5 gpc6002 (
      {stage1_2[172], stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[27],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc606_5 gpc6003 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182], stage1_2[183]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[28],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc606_5 gpc6004 (
      {stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187], stage1_2[188], stage1_2[189]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[29],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc606_5 gpc6005 (
      {stage1_2[190], stage1_2[191], stage1_2[192], stage1_2[193], stage1_2[194], stage1_2[195]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[30],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc606_5 gpc6006 (
      {stage1_2[196], stage1_2[197], stage1_2[198], stage1_2[199], stage1_2[200], stage1_2[201]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[31],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc606_5 gpc6007 (
      {stage1_2[202], stage1_2[203], stage1_2[204], stage1_2[205], stage1_2[206], stage1_2[207]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[32],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc1415_5 gpc6008 (
      {stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92]},
      {stage1_4[126]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[21],stage2_5[33],stage2_4[60],stage2_3[60]}
   );
   gpc1415_5 gpc6009 (
      {stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage1_4[127]},
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7]},
      {stage1_6[1]},
      {stage2_7[1],stage2_6[22],stage2_5[34],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc6010 (
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102]},
      {stage1_4[128]},
      {stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13]},
      {stage2_7[2],stage2_6[23],stage2_5[35],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc6011 (
      {stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage1_4[129]},
      {stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19]},
      {stage2_7[3],stage2_6[24],stage2_5[36],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc6012 (
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112]},
      {stage1_4[130]},
      {stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25]},
      {stage2_7[4],stage2_6[25],stage2_5[37],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc6013 (
      {stage1_3[113], stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117]},
      {stage1_4[131]},
      {stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31]},
      {stage2_7[5],stage2_6[26],stage2_5[38],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc6014 (
      {stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122]},
      {stage1_4[132]},
      {stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37]},
      {stage2_7[6],stage2_6[27],stage2_5[39],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc6015 (
      {stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage1_4[133]},
      {stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43]},
      {stage2_7[7],stage2_6[28],stage2_5[40],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc6016 (
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132]},
      {stage1_4[134]},
      {stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49]},
      {stage2_7[8],stage2_6[29],stage2_5[41],stage2_4[68],stage2_3[68]}
   );
   gpc623_5 gpc6017 (
      {stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[135], stage1_4[136]},
      {stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55]},
      {stage2_7[9],stage2_6[30],stage2_5[42],stage2_4[69],stage2_3[69]}
   );
   gpc623_5 gpc6018 (
      {stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[137], stage1_4[138]},
      {stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61]},
      {stage2_7[10],stage2_6[31],stage2_5[43],stage2_4[70],stage2_3[70]}
   );
   gpc606_5 gpc6019 (
      {stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[11],stage2_6[32],stage2_5[44],stage2_4[71]}
   );
   gpc606_5 gpc6020 (
      {stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[12],stage2_6[33],stage2_5[45],stage2_4[72]}
   );
   gpc606_5 gpc6021 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[13],stage2_6[34],stage2_5[46],stage2_4[73]}
   );
   gpc606_5 gpc6022 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162]},
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage2_8[3],stage2_7[14],stage2_6[35],stage2_5[47],stage2_4[74]}
   );
   gpc606_5 gpc6023 (
      {stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168]},
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage2_8[4],stage2_7[15],stage2_6[36],stage2_5[48],stage2_4[75]}
   );
   gpc606_5 gpc6024 (
      {stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174]},
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36], stage1_6[37]},
      {stage2_8[5],stage2_7[16],stage2_6[37],stage2_5[49],stage2_4[76]}
   );
   gpc606_5 gpc6025 (
      {stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42], stage1_6[43]},
      {stage2_8[6],stage2_7[17],stage2_6[38],stage2_5[50],stage2_4[77]}
   );
   gpc606_5 gpc6026 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49]},
      {stage2_8[7],stage2_7[18],stage2_6[39],stage2_5[51],stage2_4[78]}
   );
   gpc606_5 gpc6027 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192]},
      {stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage2_8[8],stage2_7[19],stage2_6[40],stage2_5[52],stage2_4[79]}
   );
   gpc606_5 gpc6028 (
      {stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198]},
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage2_8[9],stage2_7[20],stage2_6[41],stage2_5[53],stage2_4[80]}
   );
   gpc606_5 gpc6029 (
      {stage1_4[199], stage1_4[200], stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204]},
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66], stage1_6[67]},
      {stage2_8[10],stage2_7[21],stage2_6[42],stage2_5[54],stage2_4[81]}
   );
   gpc606_5 gpc6030 (
      {stage1_4[205], stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72], stage1_6[73]},
      {stage2_8[11],stage2_7[22],stage2_6[43],stage2_5[55],stage2_4[82]}
   );
   gpc606_5 gpc6031 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79]},
      {stage2_8[12],stage2_7[23],stage2_6[44],stage2_5[56],stage2_4[83]}
   );
   gpc606_5 gpc6032 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221], stage1_4[222]},
      {stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage2_8[13],stage2_7[24],stage2_6[45],stage2_5[57],stage2_4[84]}
   );
   gpc606_5 gpc6033 (
      {stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227], stage1_4[228]},
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage2_8[14],stage2_7[25],stage2_6[46],stage2_5[58],stage2_4[85]}
   );
   gpc606_5 gpc6034 (
      {stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233], stage1_4[234]},
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96], stage1_6[97]},
      {stage2_8[15],stage2_7[26],stage2_6[47],stage2_5[59],stage2_4[86]}
   );
   gpc606_5 gpc6035 (
      {stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239], stage1_4[240]},
      {stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102], stage1_6[103]},
      {stage2_8[16],stage2_7[27],stage2_6[48],stage2_5[60],stage2_4[87]}
   );
   gpc606_5 gpc6036 (
      {stage1_4[241], stage1_4[242], stage1_4[243], stage1_4[244], stage1_4[245], stage1_4[246]},
      {stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108], stage1_6[109]},
      {stage2_8[17],stage2_7[28],stage2_6[49],stage2_5[61],stage2_4[88]}
   );
   gpc606_5 gpc6037 (
      {stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[18],stage2_7[29],stage2_6[50],stage2_5[62]}
   );
   gpc606_5 gpc6038 (
      {stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[19],stage2_7[30],stage2_6[51],stage2_5[63]}
   );
   gpc606_5 gpc6039 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[20],stage2_7[31],stage2_6[52],stage2_5[64]}
   );
   gpc606_5 gpc6040 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[21],stage2_7[32],stage2_6[53],stage2_5[65]}
   );
   gpc606_5 gpc6041 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[22],stage2_7[33],stage2_6[54],stage2_5[66]}
   );
   gpc606_5 gpc6042 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[23],stage2_7[34],stage2_6[55],stage2_5[67]}
   );
   gpc606_5 gpc6043 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[24],stage2_7[35],stage2_6[56],stage2_5[68]}
   );
   gpc606_5 gpc6044 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[25],stage2_7[36],stage2_6[57],stage2_5[69]}
   );
   gpc606_5 gpc6045 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[26],stage2_7[37],stage2_6[58],stage2_5[70]}
   );
   gpc606_5 gpc6046 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[27],stage2_7[38],stage2_6[59],stage2_5[71]}
   );
   gpc606_5 gpc6047 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[28],stage2_7[39],stage2_6[60],stage2_5[72]}
   );
   gpc606_5 gpc6048 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[29],stage2_7[40],stage2_6[61],stage2_5[73]}
   );
   gpc606_5 gpc6049 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[30],stage2_7[41],stage2_6[62],stage2_5[74]}
   );
   gpc606_5 gpc6050 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[31],stage2_7[42],stage2_6[63],stage2_5[75]}
   );
   gpc606_5 gpc6051 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[32],stage2_7[43],stage2_6[64],stage2_5[76]}
   );
   gpc606_5 gpc6052 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[33],stage2_7[44],stage2_6[65],stage2_5[77]}
   );
   gpc606_5 gpc6053 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[34],stage2_7[45],stage2_6[66],stage2_5[78]}
   );
   gpc606_5 gpc6054 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[35],stage2_7[46],stage2_6[67],stage2_5[79]}
   );
   gpc606_5 gpc6055 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[36],stage2_7[47],stage2_6[68],stage2_5[80]}
   );
   gpc606_5 gpc6056 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[114], stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage2_9[19],stage2_8[37],stage2_7[48],stage2_6[69],stage2_5[81]}
   );
   gpc606_5 gpc6057 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage2_9[20],stage2_8[38],stage2_7[49],stage2_6[70],stage2_5[82]}
   );
   gpc615_5 gpc6058 (
      {stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_7[126]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[21],stage2_8[39],stage2_7[50],stage2_6[71]}
   );
   gpc615_5 gpc6059 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_7[127]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[22],stage2_8[40],stage2_7[51],stage2_6[72]}
   );
   gpc615_5 gpc6060 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124]},
      {stage1_7[128]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[23],stage2_8[41],stage2_7[52],stage2_6[73]}
   );
   gpc615_5 gpc6061 (
      {stage1_6[125], stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129]},
      {stage1_7[129]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[24],stage2_8[42],stage2_7[53],stage2_6[74]}
   );
   gpc615_5 gpc6062 (
      {stage1_6[130], stage1_6[131], stage1_6[132], stage1_6[133], stage1_6[134]},
      {stage1_7[130]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[25],stage2_8[43],stage2_7[54],stage2_6[75]}
   );
   gpc615_5 gpc6063 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[26],stage2_8[44],stage2_7[55]}
   );
   gpc615_5 gpc6064 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[27],stage2_8[45],stage2_7[56]}
   );
   gpc615_5 gpc6065 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[28],stage2_8[46],stage2_7[57]}
   );
   gpc615_5 gpc6066 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[29],stage2_8[47],stage2_7[58]}
   );
   gpc615_5 gpc6067 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[30],stage2_8[48],stage2_7[59]}
   );
   gpc615_5 gpc6068 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[31],stage2_8[49],stage2_7[60]}
   );
   gpc615_5 gpc6069 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[36]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[32],stage2_8[50],stage2_7[61]}
   );
   gpc615_5 gpc6070 (
      {stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170]},
      {stage1_8[37]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[33],stage2_8[51],stage2_7[62]}
   );
   gpc615_5 gpc6071 (
      {stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175]},
      {stage1_8[38]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[34],stage2_8[52],stage2_7[63]}
   );
   gpc615_5 gpc6072 (
      {stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_8[39]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[35],stage2_8[53],stage2_7[64]}
   );
   gpc615_5 gpc6073 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185]},
      {stage1_8[40]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[36],stage2_8[54],stage2_7[65]}
   );
   gpc615_5 gpc6074 (
      {stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190]},
      {stage1_8[41]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[37],stage2_8[55],stage2_7[66]}
   );
   gpc615_5 gpc6075 (
      {stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195]},
      {stage1_8[42]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[38],stage2_8[56],stage2_7[67]}
   );
   gpc615_5 gpc6076 (
      {stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200]},
      {stage1_8[43]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[39],stage2_8[57],stage2_7[68]}
   );
   gpc615_5 gpc6077 (
      {stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205]},
      {stage1_8[44]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[40],stage2_8[58],stage2_7[69]}
   );
   gpc615_5 gpc6078 (
      {stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_8[45]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[41],stage2_8[59],stage2_7[70]}
   );
   gpc615_5 gpc6079 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215]},
      {stage1_8[46]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[42],stage2_8[60],stage2_7[71]}
   );
   gpc615_5 gpc6080 (
      {stage1_7[216], stage1_7[217], stage1_7[218], stage1_7[219], stage1_7[220]},
      {stage1_8[47]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[43],stage2_8[61],stage2_7[72]}
   );
   gpc615_5 gpc6081 (
      {stage1_7[221], stage1_7[222], stage1_7[223], stage1_7[224], stage1_7[225]},
      {stage1_8[48]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[44],stage2_8[62],stage2_7[73]}
   );
   gpc615_5 gpc6082 (
      {stage1_7[226], stage1_7[227], stage1_7[228], stage1_7[229], stage1_7[230]},
      {stage1_8[49]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[45],stage2_8[63],stage2_7[74]}
   );
   gpc615_5 gpc6083 (
      {stage1_7[231], stage1_7[232], stage1_7[233], stage1_7[234], stage1_7[235]},
      {stage1_8[50]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[46],stage2_8[64],stage2_7[75]}
   );
   gpc615_5 gpc6084 (
      {stage1_7[236], stage1_7[237], stage1_7[238], stage1_7[239], stage1_7[240]},
      {stage1_8[51]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[26],stage2_9[47],stage2_8[65],stage2_7[76]}
   );
   gpc615_5 gpc6085 (
      {stage1_7[241], stage1_7[242], stage1_7[243], stage1_7[244], stage1_7[245]},
      {stage1_8[52]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[27],stage2_9[48],stage2_8[66],stage2_7[77]}
   );
   gpc615_5 gpc6086 (
      {stage1_7[246], stage1_7[247], stage1_7[248], stage1_7[249], stage1_7[250]},
      {stage1_8[53]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[28],stage2_9[49],stage2_8[67],stage2_7[78]}
   );
   gpc615_5 gpc6087 (
      {stage1_7[251], stage1_7[252], stage1_7[253], stage1_7[254], stage1_7[255]},
      {stage1_8[54]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[29],stage2_9[50],stage2_8[68],stage2_7[79]}
   );
   gpc615_5 gpc6088 (
      {stage1_7[256], stage1_7[257], stage1_7[258], stage1_7[259], stage1_7[260]},
      {stage1_8[55]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[30],stage2_9[51],stage2_8[69],stage2_7[80]}
   );
   gpc615_5 gpc6089 (
      {stage1_7[261], stage1_7[262], stage1_7[263], stage1_7[264], stage1_7[265]},
      {stage1_8[56]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[31],stage2_9[52],stage2_8[70],stage2_7[81]}
   );
   gpc615_5 gpc6090 (
      {stage1_7[266], stage1_7[267], stage1_7[268], stage1_7[269], stage1_7[270]},
      {stage1_8[57]},
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage2_11[27],stage2_10[32],stage2_9[53],stage2_8[71],stage2_7[82]}
   );
   gpc615_5 gpc6091 (
      {stage1_7[271], stage1_7[272], stage1_7[273], stage1_7[274], stage1_7[275]},
      {stage1_8[58]},
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage2_11[28],stage2_10[33],stage2_9[54],stage2_8[72],stage2_7[83]}
   );
   gpc615_5 gpc6092 (
      {stage1_7[276], stage1_7[277], stage1_7[278], stage1_7[279], stage1_7[280]},
      {stage1_8[59]},
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage2_11[29],stage2_10[34],stage2_9[55],stage2_8[73],stage2_7[84]}
   );
   gpc615_5 gpc6093 (
      {stage1_7[281], stage1_7[282], stage1_7[283], stage1_7[284], stage1_7[285]},
      {stage1_8[60]},
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage2_11[30],stage2_10[35],stage2_9[56],stage2_8[74],stage2_7[85]}
   );
   gpc615_5 gpc6094 (
      {stage1_7[286], stage1_7[287], stage1_7[288], stage1_7[289], stage1_7[290]},
      {stage1_8[61]},
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage2_11[31],stage2_10[36],stage2_9[57],stage2_8[75],stage2_7[86]}
   );
   gpc615_5 gpc6095 (
      {stage1_7[291], stage1_7[292], stage1_7[293], stage1_7[294], stage1_7[295]},
      {stage1_8[62]},
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage2_11[32],stage2_10[37],stage2_9[58],stage2_8[76],stage2_7[87]}
   );
   gpc615_5 gpc6096 (
      {stage1_7[296], stage1_7[297], stage1_7[298], stage1_7[299], stage1_7[300]},
      {stage1_8[63]},
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage2_11[33],stage2_10[38],stage2_9[59],stage2_8[77],stage2_7[88]}
   );
   gpc615_5 gpc6097 (
      {stage1_7[301], stage1_7[302], stage1_7[303], stage1_7[304], stage1_7[305]},
      {stage1_8[64]},
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage2_11[34],stage2_10[39],stage2_9[60],stage2_8[78],stage2_7[89]}
   );
   gpc615_5 gpc6098 (
      {stage1_7[306], stage1_7[307], stage1_7[308], stage1_7[309], stage1_7[310]},
      {stage1_8[65]},
      {stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213], stage1_9[214], stage1_9[215]},
      {stage2_11[35],stage2_10[40],stage2_9[61],stage2_8[79],stage2_7[90]}
   );
   gpc615_5 gpc6099 (
      {stage1_7[311], stage1_7[312], stage1_7[313], stage1_7[314], stage1_7[315]},
      {stage1_8[66]},
      {stage1_9[216], stage1_9[217], stage1_9[218], stage1_9[219], stage1_9[220], stage1_9[221]},
      {stage2_11[36],stage2_10[41],stage2_9[62],stage2_8[80],stage2_7[91]}
   );
   gpc615_5 gpc6100 (
      {stage1_7[316], stage1_7[317], stage1_7[318], stage1_7[319], stage1_7[320]},
      {stage1_8[67]},
      {stage1_9[222], stage1_9[223], stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227]},
      {stage2_11[37],stage2_10[42],stage2_9[63],stage2_8[81],stage2_7[92]}
   );
   gpc615_5 gpc6101 (
      {stage1_7[321], stage1_7[322], stage1_7[323], stage1_7[324], stage1_7[325]},
      {stage1_8[68]},
      {stage1_9[228], stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage2_11[38],stage2_10[43],stage2_9[64],stage2_8[82],stage2_7[93]}
   );
   gpc615_5 gpc6102 (
      {stage1_7[326], stage1_7[327], stage1_7[328], stage1_7[329], stage1_7[330]},
      {stage1_8[69]},
      {stage1_9[234], stage1_9[235], stage1_9[236], stage1_9[237], stage1_9[238], stage1_9[239]},
      {stage2_11[39],stage2_10[44],stage2_9[65],stage2_8[83],stage2_7[94]}
   );
   gpc615_5 gpc6103 (
      {stage1_7[331], stage1_7[332], stage1_7[333], stage1_7[334], stage1_7[335]},
      {stage1_8[70]},
      {stage1_9[240], stage1_9[241], stage1_9[242], stage1_9[243], stage1_9[244], stage1_9[245]},
      {stage2_11[40],stage2_10[45],stage2_9[66],stage2_8[84],stage2_7[95]}
   );
   gpc615_5 gpc6104 (
      {stage1_7[336], stage1_7[337], stage1_7[338], stage1_7[339], 1'b0},
      {stage1_8[71]},
      {stage1_9[246], stage1_9[247], stage1_9[248], stage1_9[249], stage1_9[250], stage1_9[251]},
      {stage2_11[41],stage2_10[46],stage2_9[67],stage2_8[85],stage2_7[96]}
   );
   gpc606_5 gpc6105 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[42],stage2_10[47],stage2_9[68],stage2_8[86]}
   );
   gpc606_5 gpc6106 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[43],stage2_10[48],stage2_9[69],stage2_8[87]}
   );
   gpc606_5 gpc6107 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[44],stage2_10[49],stage2_9[70],stage2_8[88]}
   );
   gpc606_5 gpc6108 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[45],stage2_10[50],stage2_9[71],stage2_8[89]}
   );
   gpc606_5 gpc6109 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[46],stage2_10[51],stage2_9[72],stage2_8[90]}
   );
   gpc606_5 gpc6110 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[47],stage2_10[52],stage2_9[73],stage2_8[91]}
   );
   gpc606_5 gpc6111 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[48],stage2_10[53],stage2_9[74],stage2_8[92]}
   );
   gpc606_5 gpc6112 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[49],stage2_10[54],stage2_9[75],stage2_8[93]}
   );
   gpc606_5 gpc6113 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[50],stage2_10[55],stage2_9[76],stage2_8[94]}
   );
   gpc606_5 gpc6114 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[51],stage2_10[56],stage2_9[77],stage2_8[95]}
   );
   gpc606_5 gpc6115 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[52],stage2_10[57],stage2_9[78],stage2_8[96]}
   );
   gpc606_5 gpc6116 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[53],stage2_10[58],stage2_9[79],stage2_8[97]}
   );
   gpc606_5 gpc6117 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[54],stage2_10[59],stage2_9[80],stage2_8[98]}
   );
   gpc606_5 gpc6118 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[55],stage2_10[60],stage2_9[81],stage2_8[99]}
   );
   gpc606_5 gpc6119 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[56],stage2_10[61],stage2_9[82],stage2_8[100]}
   );
   gpc606_5 gpc6120 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[57],stage2_10[62],stage2_9[83],stage2_8[101]}
   );
   gpc606_5 gpc6121 (
      {stage1_9[252], stage1_9[253], stage1_9[254], stage1_9[255], stage1_9[256], stage1_9[257]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[16],stage2_11[58],stage2_10[63],stage2_9[84]}
   );
   gpc606_5 gpc6122 (
      {stage1_9[258], stage1_9[259], stage1_9[260], stage1_9[261], stage1_9[262], stage1_9[263]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[17],stage2_11[59],stage2_10[64],stage2_9[85]}
   );
   gpc606_5 gpc6123 (
      {stage1_9[264], stage1_9[265], stage1_9[266], stage1_9[267], stage1_9[268], stage1_9[269]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[18],stage2_11[60],stage2_10[65],stage2_9[86]}
   );
   gpc606_5 gpc6124 (
      {stage1_9[270], stage1_9[271], stage1_9[272], stage1_9[273], stage1_9[274], stage1_9[275]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[19],stage2_11[61],stage2_10[66],stage2_9[87]}
   );
   gpc606_5 gpc6125 (
      {stage1_9[276], stage1_9[277], stage1_9[278], stage1_9[279], stage1_9[280], stage1_9[281]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[20],stage2_11[62],stage2_10[67],stage2_9[88]}
   );
   gpc606_5 gpc6126 (
      {stage1_9[282], stage1_9[283], stage1_9[284], stage1_9[285], stage1_9[286], stage1_9[287]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[21],stage2_11[63],stage2_10[68],stage2_9[89]}
   );
   gpc606_5 gpc6127 (
      {stage1_9[288], stage1_9[289], stage1_9[290], stage1_9[291], stage1_9[292], stage1_9[293]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[22],stage2_11[64],stage2_10[69],stage2_9[90]}
   );
   gpc606_5 gpc6128 (
      {stage1_9[294], stage1_9[295], stage1_9[296], stage1_9[297], stage1_9[298], stage1_9[299]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[23],stage2_11[65],stage2_10[70],stage2_9[91]}
   );
   gpc606_5 gpc6129 (
      {stage1_9[300], stage1_9[301], stage1_9[302], stage1_9[303], stage1_9[304], stage1_9[305]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[24],stage2_11[66],stage2_10[71],stage2_9[92]}
   );
   gpc606_5 gpc6130 (
      {stage1_9[306], stage1_9[307], stage1_9[308], stage1_9[309], stage1_9[310], stage1_9[311]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[25],stage2_11[67],stage2_10[72],stage2_9[93]}
   );
   gpc606_5 gpc6131 (
      {stage1_9[312], stage1_9[313], stage1_9[314], stage1_9[315], stage1_9[316], stage1_9[317]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[26],stage2_11[68],stage2_10[73],stage2_9[94]}
   );
   gpc606_5 gpc6132 (
      {stage1_9[318], stage1_9[319], stage1_9[320], stage1_9[321], stage1_9[322], stage1_9[323]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[27],stage2_11[69],stage2_10[74],stage2_9[95]}
   );
   gpc606_5 gpc6133 (
      {stage1_9[324], stage1_9[325], stage1_9[326], stage1_9[327], stage1_9[328], stage1_9[329]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[28],stage2_11[70],stage2_10[75],stage2_9[96]}
   );
   gpc606_5 gpc6134 (
      {stage1_9[330], stage1_9[331], stage1_9[332], stage1_9[333], stage1_9[334], stage1_9[335]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[29],stage2_11[71],stage2_10[76],stage2_9[97]}
   );
   gpc606_5 gpc6135 (
      {stage1_9[336], stage1_9[337], stage1_9[338], stage1_9[339], stage1_9[340], stage1_9[341]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[30],stage2_11[72],stage2_10[77],stage2_9[98]}
   );
   gpc606_5 gpc6136 (
      {stage1_9[342], stage1_9[343], stage1_9[344], stage1_9[345], stage1_9[346], stage1_9[347]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[31],stage2_11[73],stage2_10[78],stage2_9[99]}
   );
   gpc606_5 gpc6137 (
      {stage1_9[348], stage1_9[349], stage1_9[350], stage1_9[351], stage1_9[352], stage1_9[353]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[32],stage2_11[74],stage2_10[79],stage2_9[100]}
   );
   gpc606_5 gpc6138 (
      {stage1_9[354], stage1_9[355], stage1_9[356], stage1_9[357], stage1_9[358], stage1_9[359]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[33],stage2_11[75],stage2_10[80],stage2_9[101]}
   );
   gpc615_5 gpc6139 (
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_11[108]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[34],stage2_11[76],stage2_10[81]}
   );
   gpc1163_5 gpc6140 (
      {stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_13[0]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[19],stage2_12[35],stage2_11[77]}
   );
   gpc1163_5 gpc6141 (
      {stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage1_13[1]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[20],stage2_12[36],stage2_11[78]}
   );
   gpc1163_5 gpc6142 (
      {stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage1_13[2]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[21],stage2_12[37],stage2_11[79]}
   );
   gpc1163_5 gpc6143 (
      {stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage1_13[3]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[22],stage2_12[38],stage2_11[80]}
   );
   gpc1163_5 gpc6144 (
      {stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage1_13[4]},
      {stage1_14[4]},
      {stage2_15[4],stage2_14[5],stage2_13[23],stage2_12[39],stage2_11[81]}
   );
   gpc1163_5 gpc6145 (
      {stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[5]},
      {stage1_14[5]},
      {stage2_15[5],stage2_14[6],stage2_13[24],stage2_12[40],stage2_11[82]}
   );
   gpc1163_5 gpc6146 (
      {stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_13[6]},
      {stage1_14[6]},
      {stage2_15[6],stage2_14[7],stage2_13[25],stage2_12[41],stage2_11[83]}
   );
   gpc1163_5 gpc6147 (
      {stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_13[7]},
      {stage1_14[7]},
      {stage2_15[7],stage2_14[8],stage2_13[26],stage2_12[42],stage2_11[84]}
   );
   gpc1163_5 gpc6148 (
      {stage1_11[133], stage1_11[134], stage1_11[135]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[8]},
      {stage1_14[8]},
      {stage2_15[8],stage2_14[9],stage2_13[27],stage2_12[43],stage2_11[85]}
   );
   gpc1163_5 gpc6149 (
      {stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_13[9]},
      {stage1_14[9]},
      {stage2_15[9],stage2_14[10],stage2_13[28],stage2_12[44],stage2_11[86]}
   );
   gpc1163_5 gpc6150 (
      {stage1_11[139], stage1_11[140], stage1_11[141]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage1_13[10]},
      {stage1_14[10]},
      {stage2_15[10],stage2_14[11],stage2_13[29],stage2_12[45],stage2_11[87]}
   );
   gpc1163_5 gpc6151 (
      {stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage1_13[11]},
      {stage1_14[11]},
      {stage2_15[11],stage2_14[12],stage2_13[30],stage2_12[46],stage2_11[88]}
   );
   gpc1163_5 gpc6152 (
      {stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage1_13[12]},
      {stage1_14[12]},
      {stage2_15[12],stage2_14[13],stage2_13[31],stage2_12[47],stage2_11[89]}
   );
   gpc1163_5 gpc6153 (
      {stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[13]},
      {stage1_14[13]},
      {stage2_15[13],stage2_14[14],stage2_13[32],stage2_12[48],stage2_11[90]}
   );
   gpc1163_5 gpc6154 (
      {stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage1_13[14]},
      {stage1_14[14]},
      {stage2_15[14],stage2_14[15],stage2_13[33],stage2_12[49],stage2_11[91]}
   );
   gpc1163_5 gpc6155 (
      {stage1_11[154], stage1_11[155], stage1_11[156]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_13[15]},
      {stage1_14[15]},
      {stage2_15[15],stage2_14[16],stage2_13[34],stage2_12[50],stage2_11[92]}
   );
   gpc1163_5 gpc6156 (
      {stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage1_13[16]},
      {stage1_14[16]},
      {stage2_15[16],stage2_14[17],stage2_13[35],stage2_12[51],stage2_11[93]}
   );
   gpc1163_5 gpc6157 (
      {stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_13[17]},
      {stage1_14[17]},
      {stage2_15[17],stage2_14[18],stage2_13[36],stage2_12[52],stage2_11[94]}
   );
   gpc1163_5 gpc6158 (
      {stage1_11[163], stage1_11[164], stage1_11[165]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[18]},
      {stage1_14[18]},
      {stage2_15[18],stage2_14[19],stage2_13[37],stage2_12[53],stage2_11[95]}
   );
   gpc1163_5 gpc6159 (
      {stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_13[19]},
      {stage1_14[19]},
      {stage2_15[19],stage2_14[20],stage2_13[38],stage2_12[54],stage2_11[96]}
   );
   gpc1163_5 gpc6160 (
      {stage1_11[169], stage1_11[170], stage1_11[171]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_13[20]},
      {stage1_14[20]},
      {stage2_15[20],stage2_14[21],stage2_13[39],stage2_12[55],stage2_11[97]}
   );
   gpc615_5 gpc6161 (
      {stage1_11[172], stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176]},
      {stage1_12[132]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[21],stage2_14[22],stage2_13[40],stage2_12[56],stage2_11[98]}
   );
   gpc615_5 gpc6162 (
      {stage1_11[177], stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181]},
      {stage1_12[133]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[22],stage2_14[23],stage2_13[41],stage2_12[57],stage2_11[99]}
   );
   gpc615_5 gpc6163 (
      {stage1_11[182], stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186]},
      {stage1_12[134]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[23],stage2_14[24],stage2_13[42],stage2_12[58],stage2_11[100]}
   );
   gpc615_5 gpc6164 (
      {stage1_11[187], stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191]},
      {stage1_12[135]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[24],stage2_14[25],stage2_13[43],stage2_12[59],stage2_11[101]}
   );
   gpc615_5 gpc6165 (
      {stage1_11[192], stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196]},
      {stage1_12[136]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[25],stage2_14[26],stage2_13[44],stage2_12[60],stage2_11[102]}
   );
   gpc615_5 gpc6166 (
      {stage1_11[197], stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201]},
      {stage1_12[137]},
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage2_15[26],stage2_14[27],stage2_13[45],stage2_12[61],stage2_11[103]}
   );
   gpc615_5 gpc6167 (
      {stage1_11[202], stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206]},
      {stage1_12[138]},
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage2_15[27],stage2_14[28],stage2_13[46],stage2_12[62],stage2_11[104]}
   );
   gpc615_5 gpc6168 (
      {stage1_11[207], stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211]},
      {stage1_12[139]},
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage2_15[28],stage2_14[29],stage2_13[47],stage2_12[63],stage2_11[105]}
   );
   gpc615_5 gpc6169 (
      {stage1_11[212], stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216]},
      {stage1_12[140]},
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage2_15[29],stage2_14[30],stage2_13[48],stage2_12[64],stage2_11[106]}
   );
   gpc615_5 gpc6170 (
      {stage1_11[217], stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221]},
      {stage1_12[141]},
      {stage1_13[75], stage1_13[76], stage1_13[77], stage1_13[78], stage1_13[79], stage1_13[80]},
      {stage2_15[30],stage2_14[31],stage2_13[49],stage2_12[65],stage2_11[107]}
   );
   gpc615_5 gpc6171 (
      {stage1_11[222], stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226]},
      {stage1_12[142]},
      {stage1_13[81], stage1_13[82], stage1_13[83], stage1_13[84], stage1_13[85], stage1_13[86]},
      {stage2_15[31],stage2_14[32],stage2_13[50],stage2_12[66],stage2_11[108]}
   );
   gpc615_5 gpc6172 (
      {stage1_11[227], stage1_11[228], stage1_11[229], stage1_11[230], stage1_11[231]},
      {stage1_12[143]},
      {stage1_13[87], stage1_13[88], stage1_13[89], stage1_13[90], stage1_13[91], stage1_13[92]},
      {stage2_15[32],stage2_14[33],stage2_13[51],stage2_12[67],stage2_11[109]}
   );
   gpc615_5 gpc6173 (
      {stage1_11[232], stage1_11[233], stage1_11[234], stage1_11[235], stage1_11[236]},
      {stage1_12[144]},
      {stage1_13[93], stage1_13[94], stage1_13[95], stage1_13[96], stage1_13[97], stage1_13[98]},
      {stage2_15[33],stage2_14[34],stage2_13[52],stage2_12[68],stage2_11[110]}
   );
   gpc615_5 gpc6174 (
      {stage1_11[237], stage1_11[238], stage1_11[239], stage1_11[240], stage1_11[241]},
      {stage1_12[145]},
      {stage1_13[99], stage1_13[100], stage1_13[101], stage1_13[102], stage1_13[103], stage1_13[104]},
      {stage2_15[34],stage2_14[35],stage2_13[53],stage2_12[69],stage2_11[111]}
   );
   gpc615_5 gpc6175 (
      {stage1_11[242], stage1_11[243], stage1_11[244], stage1_11[245], stage1_11[246]},
      {stage1_12[146]},
      {stage1_13[105], stage1_13[106], stage1_13[107], stage1_13[108], stage1_13[109], stage1_13[110]},
      {stage2_15[35],stage2_14[36],stage2_13[54],stage2_12[70],stage2_11[112]}
   );
   gpc615_5 gpc6176 (
      {stage1_11[247], stage1_11[248], stage1_11[249], stage1_11[250], stage1_11[251]},
      {stage1_12[147]},
      {stage1_13[111], stage1_13[112], stage1_13[113], stage1_13[114], stage1_13[115], stage1_13[116]},
      {stage2_15[36],stage2_14[37],stage2_13[55],stage2_12[71],stage2_11[113]}
   );
   gpc615_5 gpc6177 (
      {stage1_11[252], stage1_11[253], stage1_11[254], stage1_11[255], stage1_11[256]},
      {stage1_12[148]},
      {stage1_13[117], stage1_13[118], stage1_13[119], stage1_13[120], stage1_13[121], stage1_13[122]},
      {stage2_15[37],stage2_14[38],stage2_13[56],stage2_12[72],stage2_11[114]}
   );
   gpc615_5 gpc6178 (
      {stage1_11[257], stage1_11[258], stage1_11[259], stage1_11[260], stage1_11[261]},
      {stage1_12[149]},
      {stage1_13[123], stage1_13[124], stage1_13[125], stage1_13[126], stage1_13[127], stage1_13[128]},
      {stage2_15[38],stage2_14[39],stage2_13[57],stage2_12[73],stage2_11[115]}
   );
   gpc615_5 gpc6179 (
      {stage1_11[262], stage1_11[263], stage1_11[264], stage1_11[265], stage1_11[266]},
      {stage1_12[150]},
      {stage1_13[129], stage1_13[130], stage1_13[131], stage1_13[132], stage1_13[133], stage1_13[134]},
      {stage2_15[39],stage2_14[40],stage2_13[58],stage2_12[74],stage2_11[116]}
   );
   gpc615_5 gpc6180 (
      {stage1_11[267], stage1_11[268], stage1_11[269], stage1_11[270], stage1_11[271]},
      {stage1_12[151]},
      {stage1_13[135], stage1_13[136], stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140]},
      {stage2_15[40],stage2_14[41],stage2_13[59],stage2_12[75],stage2_11[117]}
   );
   gpc615_5 gpc6181 (
      {stage1_11[272], stage1_11[273], stage1_11[274], stage1_11[275], stage1_11[276]},
      {stage1_12[152]},
      {stage1_13[141], stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage2_15[41],stage2_14[42],stage2_13[60],stage2_12[76],stage2_11[118]}
   );
   gpc615_5 gpc6182 (
      {stage1_11[277], stage1_11[278], stage1_11[279], stage1_11[280], stage1_11[281]},
      {stage1_12[153]},
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151], stage1_13[152]},
      {stage2_15[42],stage2_14[43],stage2_13[61],stage2_12[77],stage2_11[119]}
   );
   gpc615_5 gpc6183 (
      {stage1_11[282], stage1_11[283], stage1_11[284], stage1_11[285], stage1_11[286]},
      {stage1_12[154]},
      {stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158]},
      {stage2_15[43],stage2_14[44],stage2_13[62],stage2_12[78],stage2_11[120]}
   );
   gpc615_5 gpc6184 (
      {stage1_11[287], stage1_11[288], stage1_11[289], stage1_11[290], stage1_11[291]},
      {stage1_12[155]},
      {stage1_13[159], stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage2_15[44],stage2_14[45],stage2_13[63],stage2_12[79],stage2_11[121]}
   );
   gpc615_5 gpc6185 (
      {stage1_11[292], stage1_11[293], stage1_11[294], stage1_11[295], stage1_11[296]},
      {stage1_12[156]},
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170]},
      {stage2_15[45],stage2_14[46],stage2_13[64],stage2_12[80],stage2_11[122]}
   );
   gpc615_5 gpc6186 (
      {stage1_11[297], stage1_11[298], stage1_11[299], stage1_11[300], stage1_11[301]},
      {stage1_12[157]},
      {stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage2_15[46],stage2_14[47],stage2_13[65],stage2_12[81],stage2_11[123]}
   );
   gpc615_5 gpc6187 (
      {stage1_11[302], stage1_11[303], stage1_11[304], stage1_11[305], stage1_11[306]},
      {stage1_12[158]},
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181], stage1_13[182]},
      {stage2_15[47],stage2_14[48],stage2_13[66],stage2_12[82],stage2_11[124]}
   );
   gpc606_5 gpc6188 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26]},
      {stage2_16[0],stage2_15[48],stage2_14[49],stage2_13[67],stage2_12[83]}
   );
   gpc606_5 gpc6189 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31], stage1_14[32]},
      {stage2_16[1],stage2_15[49],stage2_14[50],stage2_13[68],stage2_12[84]}
   );
   gpc606_5 gpc6190 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37], stage1_14[38]},
      {stage2_16[2],stage2_15[50],stage2_14[51],stage2_13[69],stage2_12[85]}
   );
   gpc1163_5 gpc6191 (
      {stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[0],stage2_16[3],stage2_15[51],stage2_14[52]}
   );
   gpc1163_5 gpc6192 (
      {stage1_14[42], stage1_14[43], stage1_14[44]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[1]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[1],stage2_16[4],stage2_15[52],stage2_14[53]}
   );
   gpc1163_5 gpc6193 (
      {stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[2]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[2],stage2_16[5],stage2_15[53],stage2_14[54]}
   );
   gpc1163_5 gpc6194 (
      {stage1_14[48], stage1_14[49], stage1_14[50]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[3]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[3],stage2_16[6],stage2_15[54],stage2_14[55]}
   );
   gpc1163_5 gpc6195 (
      {stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[4]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[4],stage2_16[7],stage2_15[55],stage2_14[56]}
   );
   gpc1163_5 gpc6196 (
      {stage1_14[54], stage1_14[55], stage1_14[56]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[5]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[5],stage2_16[8],stage2_15[56],stage2_14[57]}
   );
   gpc1163_5 gpc6197 (
      {stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage1_16[6]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[6],stage2_16[9],stage2_15[57],stage2_14[58]}
   );
   gpc1163_5 gpc6198 (
      {stage1_14[60], stage1_14[61], stage1_14[62]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[7]},
      {stage1_17[7]},
      {stage2_18[7],stage2_17[7],stage2_16[10],stage2_15[58],stage2_14[59]}
   );
   gpc1163_5 gpc6199 (
      {stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[8]},
      {stage1_17[8]},
      {stage2_18[8],stage2_17[8],stage2_16[11],stage2_15[59],stage2_14[60]}
   );
   gpc1163_5 gpc6200 (
      {stage1_14[66], stage1_14[67], stage1_14[68]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage1_16[9]},
      {stage1_17[9]},
      {stage2_18[9],stage2_17[9],stage2_16[12],stage2_15[60],stage2_14[61]}
   );
   gpc1163_5 gpc6201 (
      {stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_16[10]},
      {stage1_17[10]},
      {stage2_18[10],stage2_17[10],stage2_16[13],stage2_15[61],stage2_14[62]}
   );
   gpc1163_5 gpc6202 (
      {stage1_14[72], stage1_14[73], stage1_14[74]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage1_16[11]},
      {stage1_17[11]},
      {stage2_18[11],stage2_17[11],stage2_16[14],stage2_15[62],stage2_14[63]}
   );
   gpc1163_5 gpc6203 (
      {stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[12]},
      {stage1_17[12]},
      {stage2_18[12],stage2_17[12],stage2_16[15],stage2_15[63],stage2_14[64]}
   );
   gpc1163_5 gpc6204 (
      {stage1_14[78], stage1_14[79], stage1_14[80]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[13]},
      {stage1_17[13]},
      {stage2_18[13],stage2_17[13],stage2_16[16],stage2_15[64],stage2_14[65]}
   );
   gpc1163_5 gpc6205 (
      {stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage1_16[14]},
      {stage1_17[14]},
      {stage2_18[14],stage2_17[14],stage2_16[17],stage2_15[65],stage2_14[66]}
   );
   gpc1163_5 gpc6206 (
      {stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage1_16[15]},
      {stage1_17[15]},
      {stage2_18[15],stage2_17[15],stage2_16[18],stage2_15[66],stage2_14[67]}
   );
   gpc1163_5 gpc6207 (
      {stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage1_16[16]},
      {stage1_17[16]},
      {stage2_18[16],stage2_17[16],stage2_16[19],stage2_15[67],stage2_14[68]}
   );
   gpc1163_5 gpc6208 (
      {stage1_14[90], stage1_14[91], stage1_14[92]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[17]},
      {stage1_17[17]},
      {stage2_18[17],stage2_17[17],stage2_16[20],stage2_15[68],stage2_14[69]}
   );
   gpc1163_5 gpc6209 (
      {stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage1_16[18]},
      {stage1_17[18]},
      {stage2_18[18],stage2_17[18],stage2_16[21],stage2_15[69],stage2_14[70]}
   );
   gpc1163_5 gpc6210 (
      {stage1_14[96], stage1_14[97], stage1_14[98]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage1_16[19]},
      {stage1_17[19]},
      {stage2_18[19],stage2_17[19],stage2_16[22],stage2_15[70],stage2_14[71]}
   );
   gpc1163_5 gpc6211 (
      {stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage1_16[20]},
      {stage1_17[20]},
      {stage2_18[20],stage2_17[20],stage2_16[23],stage2_15[71],stage2_14[72]}
   );
   gpc1163_5 gpc6212 (
      {stage1_14[102], stage1_14[103], stage1_14[104]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage1_16[21]},
      {stage1_17[21]},
      {stage2_18[21],stage2_17[21],stage2_16[24],stage2_15[72],stage2_14[73]}
   );
   gpc1163_5 gpc6213 (
      {stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage1_16[22]},
      {stage1_17[22]},
      {stage2_18[22],stage2_17[22],stage2_16[25],stage2_15[73],stage2_14[74]}
   );
   gpc1163_5 gpc6214 (
      {stage1_14[108], stage1_14[109], stage1_14[110]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage1_16[23]},
      {stage1_17[23]},
      {stage2_18[23],stage2_17[23],stage2_16[26],stage2_15[74],stage2_14[75]}
   );
   gpc1163_5 gpc6215 (
      {stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage1_16[24]},
      {stage1_17[24]},
      {stage2_18[24],stage2_17[24],stage2_16[27],stage2_15[75],stage2_14[76]}
   );
   gpc1163_5 gpc6216 (
      {stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage1_16[25]},
      {stage1_17[25]},
      {stage2_18[25],stage2_17[25],stage2_16[28],stage2_15[76],stage2_14[77]}
   );
   gpc1163_5 gpc6217 (
      {stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[26]},
      {stage1_17[26]},
      {stage2_18[26],stage2_17[26],stage2_16[29],stage2_15[77],stage2_14[78]}
   );
   gpc1163_5 gpc6218 (
      {stage1_14[120], stage1_14[121], stage1_14[122]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage1_16[27]},
      {stage1_17[27]},
      {stage2_18[27],stage2_17[27],stage2_16[30],stage2_15[78],stage2_14[79]}
   );
   gpc1163_5 gpc6219 (
      {stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage1_16[28]},
      {stage1_17[28]},
      {stage2_18[28],stage2_17[28],stage2_16[31],stage2_15[79],stage2_14[80]}
   );
   gpc1163_5 gpc6220 (
      {stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage1_16[29]},
      {stage1_17[29]},
      {stage2_18[29],stage2_17[29],stage2_16[32],stage2_15[80],stage2_14[81]}
   );
   gpc1163_5 gpc6221 (
      {stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage1_16[30]},
      {stage1_17[30]},
      {stage2_18[30],stage2_17[30],stage2_16[33],stage2_15[81],stage2_14[82]}
   );
   gpc1163_5 gpc6222 (
      {stage1_14[132], stage1_14[133], stage1_14[134]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[31]},
      {stage1_17[31]},
      {stage2_18[31],stage2_17[31],stage2_16[34],stage2_15[82],stage2_14[83]}
   );
   gpc606_5 gpc6223 (
      {stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140]},
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage2_18[32],stage2_17[32],stage2_16[35],stage2_15[83],stage2_14[84]}
   );
   gpc606_5 gpc6224 (
      {stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage2_18[33],stage2_17[33],stage2_16[36],stage2_15[84],stage2_14[85]}
   );
   gpc606_5 gpc6225 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152]},
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage2_18[34],stage2_17[34],stage2_16[37],stage2_15[85],stage2_14[86]}
   );
   gpc606_5 gpc6226 (
      {stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage2_18[35],stage2_17[35],stage2_16[38],stage2_15[86],stage2_14[87]}
   );
   gpc606_5 gpc6227 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163], stage1_14[164]},
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage2_18[36],stage2_17[36],stage2_16[39],stage2_15[87],stage2_14[88]}
   );
   gpc606_5 gpc6228 (
      {stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170]},
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage2_18[37],stage2_17[37],stage2_16[40],stage2_15[88],stage2_14[89]}
   );
   gpc615_5 gpc6229 (
      {stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_15[192]},
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage2_18[38],stage2_17[38],stage2_16[41],stage2_15[89],stage2_14[90]}
   );
   gpc615_5 gpc6230 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180]},
      {stage1_15[193]},
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage2_18[39],stage2_17[39],stage2_16[42],stage2_15[90],stage2_14[91]}
   );
   gpc615_5 gpc6231 (
      {stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage1_15[194]},
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage2_18[40],stage2_17[40],stage2_16[43],stage2_15[91],stage2_14[92]}
   );
   gpc615_5 gpc6232 (
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190]},
      {stage1_15[195]},
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage2_18[41],stage2_17[41],stage2_16[44],stage2_15[92],stage2_14[93]}
   );
   gpc615_5 gpc6233 (
      {stage1_14[191], stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195]},
      {stage1_15[196]},
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage2_18[42],stage2_17[42],stage2_16[45],stage2_15[93],stage2_14[94]}
   );
   gpc615_5 gpc6234 (
      {stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200]},
      {stage1_15[197]},
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage2_18[43],stage2_17[43],stage2_16[46],stage2_15[94],stage2_14[95]}
   );
   gpc615_5 gpc6235 (
      {stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_15[198]},
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage2_18[44],stage2_17[44],stage2_16[47],stage2_15[95],stage2_14[96]}
   );
   gpc615_5 gpc6236 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[199]},
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage2_18[45],stage2_17[45],stage2_16[48],stage2_15[96],stage2_14[97]}
   );
   gpc615_5 gpc6237 (
      {stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage1_15[200]},
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage2_18[46],stage2_17[46],stage2_16[49],stage2_15[97],stage2_14[98]}
   );
   gpc615_5 gpc6238 (
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220]},
      {stage1_15[201]},
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage2_18[47],stage2_17[47],stage2_16[50],stage2_15[98],stage2_14[99]}
   );
   gpc615_5 gpc6239 (
      {stage1_14[221], stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225]},
      {stage1_15[202]},
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage2_18[48],stage2_17[48],stage2_16[51],stage2_15[99],stage2_14[100]}
   );
   gpc615_5 gpc6240 (
      {stage1_14[226], stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230]},
      {stage1_15[203]},
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage2_18[49],stage2_17[49],stage2_16[52],stage2_15[100],stage2_14[101]}
   );
   gpc615_5 gpc6241 (
      {stage1_14[231], stage1_14[232], stage1_14[233], stage1_14[234], stage1_14[235]},
      {stage1_15[204]},
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage2_18[50],stage2_17[50],stage2_16[53],stage2_15[101],stage2_14[102]}
   );
   gpc615_5 gpc6242 (
      {stage1_14[236], stage1_14[237], stage1_14[238], stage1_14[239], stage1_14[240]},
      {stage1_15[205]},
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage2_18[51],stage2_17[51],stage2_16[54],stage2_15[102],stage2_14[103]}
   );
   gpc615_5 gpc6243 (
      {stage1_14[241], stage1_14[242], stage1_14[243], stage1_14[244], stage1_14[245]},
      {stage1_15[206]},
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage2_18[52],stage2_17[52],stage2_16[55],stage2_15[103],stage2_14[104]}
   );
   gpc1406_5 gpc6244 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211], stage1_15[212]},
      {stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[53],stage2_17[53],stage2_16[56],stage2_15[104]}
   );
   gpc1406_5 gpc6245 (
      {stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216], stage1_15[217], stage1_15[218]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39]},
      {stage1_18[1]},
      {stage2_19[1],stage2_18[54],stage2_17[54],stage2_16[57],stage2_15[105]}
   );
   gpc606_5 gpc6246 (
      {stage1_15[219], stage1_15[220], stage1_15[221], stage1_15[222], stage1_15[223], stage1_15[224]},
      {stage1_17[40], stage1_17[41], stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45]},
      {stage2_19[2],stage2_18[55],stage2_17[55],stage2_16[58],stage2_15[106]}
   );
   gpc606_5 gpc6247 (
      {stage1_15[225], stage1_15[226], stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230]},
      {stage1_17[46], stage1_17[47], stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51]},
      {stage2_19[3],stage2_18[56],stage2_17[56],stage2_16[59],stage2_15[107]}
   );
   gpc606_5 gpc6248 (
      {stage1_15[231], stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_17[52], stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage2_19[4],stage2_18[57],stage2_17[57],stage2_16[60],stage2_15[108]}
   );
   gpc606_5 gpc6249 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241], stage1_15[242]},
      {stage1_17[58], stage1_17[59], stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63]},
      {stage2_19[5],stage2_18[58],stage2_17[58],stage2_16[61],stage2_15[109]}
   );
   gpc606_5 gpc6250 (
      {stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246], stage1_15[247], stage1_15[248]},
      {stage1_17[64], stage1_17[65], stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69]},
      {stage2_19[6],stage2_18[59],stage2_17[59],stage2_16[62],stage2_15[110]}
   );
   gpc606_5 gpc6251 (
      {stage1_15[249], stage1_15[250], stage1_15[251], stage1_15[252], stage1_15[253], stage1_15[254]},
      {stage1_17[70], stage1_17[71], stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75]},
      {stage2_19[7],stage2_18[60],stage2_17[60],stage2_16[63],stage2_15[111]}
   );
   gpc606_5 gpc6252 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6], stage1_18[7]},
      {stage2_20[0],stage2_19[8],stage2_18[61],stage2_17[61],stage2_16[64]}
   );
   gpc606_5 gpc6253 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12], stage1_18[13]},
      {stage2_20[1],stage2_19[9],stage2_18[62],stage2_17[62],stage2_16[65]}
   );
   gpc606_5 gpc6254 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18], stage1_18[19]},
      {stage2_20[2],stage2_19[10],stage2_18[63],stage2_17[63],stage2_16[66]}
   );
   gpc606_5 gpc6255 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180], stage1_16[181]},
      {stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25]},
      {stage2_20[3],stage2_19[11],stage2_18[64],stage2_17[64],stage2_16[67]}
   );
   gpc606_5 gpc6256 (
      {stage1_17[76], stage1_17[77], stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[4],stage2_19[12],stage2_18[65],stage2_17[65]}
   );
   gpc606_5 gpc6257 (
      {stage1_17[82], stage1_17[83], stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[5],stage2_19[13],stage2_18[66],stage2_17[66]}
   );
   gpc606_5 gpc6258 (
      {stage1_17[88], stage1_17[89], stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[6],stage2_19[14],stage2_18[67],stage2_17[67]}
   );
   gpc606_5 gpc6259 (
      {stage1_17[94], stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[7],stage2_19[15],stage2_18[68],stage2_17[68]}
   );
   gpc606_5 gpc6260 (
      {stage1_17[100], stage1_17[101], stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[8],stage2_19[16],stage2_18[69],stage2_17[69]}
   );
   gpc606_5 gpc6261 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[9],stage2_19[17],stage2_18[70],stage2_17[70]}
   );
   gpc606_5 gpc6262 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[10],stage2_19[18],stage2_18[71],stage2_17[71]}
   );
   gpc606_5 gpc6263 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[11],stage2_19[19],stage2_18[72],stage2_17[72]}
   );
   gpc606_5 gpc6264 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[12],stage2_19[20],stage2_18[73],stage2_17[73]}
   );
   gpc606_5 gpc6265 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[13],stage2_19[21],stage2_18[74],stage2_17[74]}
   );
   gpc606_5 gpc6266 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[14],stage2_19[22],stage2_18[75],stage2_17[75]}
   );
   gpc606_5 gpc6267 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[15],stage2_19[23],stage2_18[76],stage2_17[76]}
   );
   gpc606_5 gpc6268 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[16],stage2_19[24],stage2_18[77],stage2_17[77]}
   );
   gpc606_5 gpc6269 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[17],stage2_19[25],stage2_18[78],stage2_17[78]}
   );
   gpc606_5 gpc6270 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[18],stage2_19[26],stage2_18[79],stage2_17[79]}
   );
   gpc606_5 gpc6271 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[19],stage2_19[27],stage2_18[80],stage2_17[80]}
   );
   gpc606_5 gpc6272 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[20],stage2_19[28],stage2_18[81],stage2_17[81]}
   );
   gpc606_5 gpc6273 (
      {stage1_17[178], stage1_17[179], stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[21],stage2_19[29],stage2_18[82],stage2_17[82]}
   );
   gpc606_5 gpc6274 (
      {stage1_17[184], stage1_17[185], stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[22],stage2_19[30],stage2_18[83],stage2_17[83]}
   );
   gpc606_5 gpc6275 (
      {stage1_17[190], stage1_17[191], stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[23],stage2_19[31],stage2_18[84],stage2_17[84]}
   );
   gpc606_5 gpc6276 (
      {stage1_17[196], stage1_17[197], stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[24],stage2_19[32],stage2_18[85],stage2_17[85]}
   );
   gpc606_5 gpc6277 (
      {stage1_17[202], stage1_17[203], stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[25],stage2_19[33],stage2_18[86],stage2_17[86]}
   );
   gpc606_5 gpc6278 (
      {stage1_17[208], stage1_17[209], stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[26],stage2_19[34],stage2_18[87],stage2_17[87]}
   );
   gpc606_5 gpc6279 (
      {stage1_17[214], stage1_17[215], stage1_17[216], stage1_17[217], 1'b0, 1'b0},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[27],stage2_19[35],stage2_18[88],stage2_17[88]}
   );
   gpc606_5 gpc6280 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[28],stage2_19[36],stage2_18[89],stage2_17[89]}
   );
   gpc606_5 gpc6281 (
      {stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[25],stage2_20[29],stage2_19[37],stage2_18[90]}
   );
   gpc606_5 gpc6282 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36], stage1_18[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[26],stage2_20[30],stage2_19[38],stage2_18[91]}
   );
   gpc606_5 gpc6283 (
      {stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42], stage1_18[43]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[27],stage2_20[31],stage2_19[39],stage2_18[92]}
   );
   gpc606_5 gpc6284 (
      {stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48], stage1_18[49]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[28],stage2_20[32],stage2_19[40],stage2_18[93]}
   );
   gpc606_5 gpc6285 (
      {stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54], stage1_18[55]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[29],stage2_20[33],stage2_19[41],stage2_18[94]}
   );
   gpc606_5 gpc6286 (
      {stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[30],stage2_20[34],stage2_19[42],stage2_18[95]}
   );
   gpc606_5 gpc6287 (
      {stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[31],stage2_20[35],stage2_19[43],stage2_18[96]}
   );
   gpc606_5 gpc6288 (
      {stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[32],stage2_20[36],stage2_19[44],stage2_18[97]}
   );
   gpc615_5 gpc6289 (
      {stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77], stage1_18[78]},
      {stage1_19[150]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[33],stage2_20[37],stage2_19[45],stage2_18[98]}
   );
   gpc615_5 gpc6290 (
      {stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_19[151]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[34],stage2_20[38],stage2_19[46],stage2_18[99]}
   );
   gpc615_5 gpc6291 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[152]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[35],stage2_20[39],stage2_19[47],stage2_18[100]}
   );
   gpc615_5 gpc6292 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[153]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[36],stage2_20[40],stage2_19[48],stage2_18[101]}
   );
   gpc615_5 gpc6293 (
      {stage1_18[94], stage1_18[95], stage1_18[96], stage1_18[97], stage1_18[98]},
      {stage1_19[154]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[37],stage2_20[41],stage2_19[49],stage2_18[102]}
   );
   gpc615_5 gpc6294 (
      {stage1_18[99], stage1_18[100], stage1_18[101], stage1_18[102], stage1_18[103]},
      {stage1_19[155]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[38],stage2_20[42],stage2_19[50],stage2_18[103]}
   );
   gpc615_5 gpc6295 (
      {stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107], stage1_18[108]},
      {stage1_19[156]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[39],stage2_20[43],stage2_19[51],stage2_18[104]}
   );
   gpc615_5 gpc6296 (
      {stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_19[157]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[40],stage2_20[44],stage2_19[52],stage2_18[105]}
   );
   gpc615_5 gpc6297 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118]},
      {stage1_19[158]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[41],stage2_20[45],stage2_19[53],stage2_18[106]}
   );
   gpc615_5 gpc6298 (
      {stage1_18[119], stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123]},
      {stage1_19[159]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[42],stage2_20[46],stage2_19[54],stage2_18[107]}
   );
   gpc615_5 gpc6299 (
      {stage1_18[124], stage1_18[125], stage1_18[126], stage1_18[127], stage1_18[128]},
      {stage1_19[160]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[43],stage2_20[47],stage2_19[55],stage2_18[108]}
   );
   gpc615_5 gpc6300 (
      {stage1_18[129], stage1_18[130], stage1_18[131], stage1_18[132], stage1_18[133]},
      {stage1_19[161]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[44],stage2_20[48],stage2_19[56],stage2_18[109]}
   );
   gpc615_5 gpc6301 (
      {stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137], stage1_18[138]},
      {stage1_19[162]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[45],stage2_20[49],stage2_19[57],stage2_18[110]}
   );
   gpc615_5 gpc6302 (
      {stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_19[163]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[46],stage2_20[50],stage2_19[58],stage2_18[111]}
   );
   gpc615_5 gpc6303 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148]},
      {stage1_19[164]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[47],stage2_20[51],stage2_19[59],stage2_18[112]}
   );
   gpc615_5 gpc6304 (
      {stage1_18[149], stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153]},
      {stage1_19[165]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[48],stage2_20[52],stage2_19[60],stage2_18[113]}
   );
   gpc615_5 gpc6305 (
      {stage1_18[154], stage1_18[155], stage1_18[156], stage1_18[157], stage1_18[158]},
      {stage1_19[166]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[49],stage2_20[53],stage2_19[61],stage2_18[114]}
   );
   gpc615_5 gpc6306 (
      {stage1_18[159], stage1_18[160], stage1_18[161], stage1_18[162], stage1_18[163]},
      {stage1_19[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[50],stage2_20[54],stage2_19[62],stage2_18[115]}
   );
   gpc615_5 gpc6307 (
      {stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167], stage1_18[168]},
      {stage1_19[168]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[51],stage2_20[55],stage2_19[63],stage2_18[116]}
   );
   gpc615_5 gpc6308 (
      {stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_19[169]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[52],stage2_20[56],stage2_19[64],stage2_18[117]}
   );
   gpc615_5 gpc6309 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[170]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[53],stage2_20[57],stage2_19[65],stage2_18[118]}
   );
   gpc615_5 gpc6310 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[171]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[54],stage2_20[58],stage2_19[66],stage2_18[119]}
   );
   gpc615_5 gpc6311 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[172]},
      {stage1_20[180], stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185]},
      {stage2_22[30],stage2_21[55],stage2_20[59],stage2_19[67],stage2_18[120]}
   );
   gpc615_5 gpc6312 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[173]},
      {stage1_20[186], stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage2_22[31],stage2_21[56],stage2_20[60],stage2_19[68],stage2_18[121]}
   );
   gpc615_5 gpc6313 (
      {stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197], stage1_18[198]},
      {stage1_19[174]},
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197]},
      {stage2_22[32],stage2_21[57],stage2_20[61],stage2_19[69],stage2_18[122]}
   );
   gpc615_5 gpc6314 (
      {stage1_18[199], stage1_18[200], stage1_18[201], stage1_18[202], stage1_18[203]},
      {stage1_19[175]},
      {stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203]},
      {stage2_22[33],stage2_21[58],stage2_20[62],stage2_19[70],stage2_18[123]}
   );
   gpc615_5 gpc6315 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[204]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[34],stage2_21[59],stage2_20[63],stage2_19[71]}
   );
   gpc615_5 gpc6316 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[205]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[35],stage2_21[60],stage2_20[64],stage2_19[72]}
   );
   gpc615_5 gpc6317 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[206]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[36],stage2_21[61],stage2_20[65],stage2_19[73]}
   );
   gpc615_5 gpc6318 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[207]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[37],stage2_21[62],stage2_20[66],stage2_19[74]}
   );
   gpc615_5 gpc6319 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[208]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[38],stage2_21[63],stage2_20[67],stage2_19[75]}
   );
   gpc606_5 gpc6320 (
      {stage1_20[209], stage1_20[210], stage1_20[211], stage1_20[212], stage1_20[213], stage1_20[214]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[39],stage2_21[64],stage2_20[68]}
   );
   gpc606_5 gpc6321 (
      {stage1_20[215], stage1_20[216], stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[40],stage2_21[65],stage2_20[69]}
   );
   gpc606_5 gpc6322 (
      {stage1_20[221], stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[41],stage2_21[66],stage2_20[70]}
   );
   gpc606_5 gpc6323 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[3],stage2_23[8],stage2_22[42],stage2_21[67]}
   );
   gpc606_5 gpc6324 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[4],stage2_23[9],stage2_22[43],stage2_21[68]}
   );
   gpc606_5 gpc6325 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[5],stage2_23[10],stage2_22[44],stage2_21[69]}
   );
   gpc606_5 gpc6326 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[6],stage2_23[11],stage2_22[45],stage2_21[70]}
   );
   gpc606_5 gpc6327 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[7],stage2_23[12],stage2_22[46],stage2_21[71]}
   );
   gpc606_5 gpc6328 (
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[8],stage2_23[13],stage2_22[47],stage2_21[72]}
   );
   gpc606_5 gpc6329 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[9],stage2_23[14],stage2_22[48],stage2_21[73]}
   );
   gpc606_5 gpc6330 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[10],stage2_23[15],stage2_22[49],stage2_21[74]}
   );
   gpc606_5 gpc6331 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[11],stage2_23[16],stage2_22[50],stage2_21[75]}
   );
   gpc606_5 gpc6332 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[12],stage2_23[17],stage2_22[51],stage2_21[76]}
   );
   gpc606_5 gpc6333 (
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[13],stage2_23[18],stage2_22[52],stage2_21[77]}
   );
   gpc606_5 gpc6334 (
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[14],stage2_23[19],stage2_22[53],stage2_21[78]}
   );
   gpc606_5 gpc6335 (
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[15],stage2_23[20],stage2_22[54],stage2_21[79]}
   );
   gpc606_5 gpc6336 (
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[16],stage2_23[21],stage2_22[55],stage2_21[80]}
   );
   gpc606_5 gpc6337 (
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[17],stage2_23[22],stage2_22[56],stage2_21[81]}
   );
   gpc606_5 gpc6338 (
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[18],stage2_23[23],stage2_22[57],stage2_21[82]}
   );
   gpc606_5 gpc6339 (
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[19],stage2_23[24],stage2_22[58],stage2_21[83]}
   );
   gpc606_5 gpc6340 (
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[20],stage2_23[25],stage2_22[59],stage2_21[84]}
   );
   gpc606_5 gpc6341 (
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[21],stage2_23[26],stage2_22[60],stage2_21[85]}
   );
   gpc606_5 gpc6342 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[22],stage2_23[27],stage2_22[61],stage2_21[86]}
   );
   gpc606_5 gpc6343 (
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[23],stage2_23[28],stage2_22[62],stage2_21[87]}
   );
   gpc606_5 gpc6344 (
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[24],stage2_23[29],stage2_22[63],stage2_21[88]}
   );
   gpc606_5 gpc6345 (
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[25],stage2_23[30],stage2_22[64],stage2_21[89]}
   );
   gpc606_5 gpc6346 (
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[26],stage2_23[31],stage2_22[65],stage2_21[90]}
   );
   gpc606_5 gpc6347 (
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[27],stage2_23[32],stage2_22[66],stage2_21[91]}
   );
   gpc606_5 gpc6348 (
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[28],stage2_23[33],stage2_22[67],stage2_21[92]}
   );
   gpc606_5 gpc6349 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[26],stage2_24[29],stage2_23[34],stage2_22[68]}
   );
   gpc615_5 gpc6350 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[156]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[27],stage2_24[30],stage2_23[35],stage2_22[69]}
   );
   gpc615_5 gpc6351 (
      {stage1_22[29], stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33]},
      {stage1_23[157]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[28],stage2_24[31],stage2_23[36],stage2_22[70]}
   );
   gpc615_5 gpc6352 (
      {stage1_22[34], stage1_22[35], stage1_22[36], stage1_22[37], stage1_22[38]},
      {stage1_23[158]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[29],stage2_24[32],stage2_23[37],stage2_22[71]}
   );
   gpc615_5 gpc6353 (
      {stage1_22[39], stage1_22[40], stage1_22[41], stage1_22[42], stage1_22[43]},
      {stage1_23[159]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[30],stage2_24[33],stage2_23[38],stage2_22[72]}
   );
   gpc615_5 gpc6354 (
      {stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47], stage1_22[48]},
      {stage1_23[160]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[31],stage2_24[34],stage2_23[39],stage2_22[73]}
   );
   gpc615_5 gpc6355 (
      {stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_23[161]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[32],stage2_24[35],stage2_23[40],stage2_22[74]}
   );
   gpc615_5 gpc6356 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58]},
      {stage1_23[162]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[33],stage2_24[36],stage2_23[41],stage2_22[75]}
   );
   gpc615_5 gpc6357 (
      {stage1_22[59], stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63]},
      {stage1_23[163]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[34],stage2_24[37],stage2_23[42],stage2_22[76]}
   );
   gpc615_5 gpc6358 (
      {stage1_22[64], stage1_22[65], stage1_22[66], stage1_22[67], stage1_22[68]},
      {stage1_23[164]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[35],stage2_24[38],stage2_23[43],stage2_22[77]}
   );
   gpc615_5 gpc6359 (
      {stage1_22[69], stage1_22[70], stage1_22[71], stage1_22[72], stage1_22[73]},
      {stage1_23[165]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[36],stage2_24[39],stage2_23[44],stage2_22[78]}
   );
   gpc615_5 gpc6360 (
      {stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77], stage1_22[78]},
      {stage1_23[166]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[37],stage2_24[40],stage2_23[45],stage2_22[79]}
   );
   gpc615_5 gpc6361 (
      {stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage1_23[167]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[38],stage2_24[41],stage2_23[46],stage2_22[80]}
   );
   gpc615_5 gpc6362 (
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88]},
      {stage1_23[168]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[39],stage2_24[42],stage2_23[47],stage2_22[81]}
   );
   gpc615_5 gpc6363 (
      {stage1_22[89], stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93]},
      {stage1_23[169]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[40],stage2_24[43],stage2_23[48],stage2_22[82]}
   );
   gpc615_5 gpc6364 (
      {stage1_22[94], stage1_22[95], stage1_22[96], stage1_22[97], stage1_22[98]},
      {stage1_23[170]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[41],stage2_24[44],stage2_23[49],stage2_22[83]}
   );
   gpc615_5 gpc6365 (
      {stage1_22[99], stage1_22[100], stage1_22[101], stage1_22[102], stage1_22[103]},
      {stage1_23[171]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[42],stage2_24[45],stage2_23[50],stage2_22[84]}
   );
   gpc615_5 gpc6366 (
      {stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108]},
      {stage1_23[172]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[43],stage2_24[46],stage2_23[51],stage2_22[85]}
   );
   gpc615_5 gpc6367 (
      {stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage1_23[173]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[44],stage2_24[47],stage2_23[52],stage2_22[86]}
   );
   gpc615_5 gpc6368 (
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118]},
      {stage1_23[174]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[45],stage2_24[48],stage2_23[53],stage2_22[87]}
   );
   gpc615_5 gpc6369 (
      {stage1_22[119], stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123]},
      {stage1_23[175]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[46],stage2_24[49],stage2_23[54],stage2_22[88]}
   );
   gpc615_5 gpc6370 (
      {stage1_22[124], stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128]},
      {stage1_23[176]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[47],stage2_24[50],stage2_23[55],stage2_22[89]}
   );
   gpc615_5 gpc6371 (
      {stage1_22[129], stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133]},
      {stage1_23[177]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[48],stage2_24[51],stage2_23[56],stage2_22[90]}
   );
   gpc615_5 gpc6372 (
      {stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138]},
      {stage1_23[178]},
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage2_26[23],stage2_25[49],stage2_24[52],stage2_23[57],stage2_22[91]}
   );
   gpc615_5 gpc6373 (
      {stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage1_23[179]},
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage2_26[24],stage2_25[50],stage2_24[53],stage2_23[58],stage2_22[92]}
   );
   gpc615_5 gpc6374 (
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148]},
      {stage1_23[180]},
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage2_26[25],stage2_25[51],stage2_24[54],stage2_23[59],stage2_22[93]}
   );
   gpc615_5 gpc6375 (
      {stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153]},
      {stage1_23[181]},
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage2_26[26],stage2_25[52],stage2_24[55],stage2_23[60],stage2_22[94]}
   );
   gpc615_5 gpc6376 (
      {stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157], stage1_22[158]},
      {stage1_23[182]},
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage2_26[27],stage2_25[53],stage2_24[56],stage2_23[61],stage2_22[95]}
   );
   gpc615_5 gpc6377 (
      {stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162], stage1_22[163]},
      {stage1_23[183]},
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage2_26[28],stage2_25[54],stage2_24[57],stage2_23[62],stage2_22[96]}
   );
   gpc615_5 gpc6378 (
      {stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167], stage1_22[168]},
      {stage1_23[184]},
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage2_26[29],stage2_25[55],stage2_24[58],stage2_23[63],stage2_22[97]}
   );
   gpc615_5 gpc6379 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173]},
      {stage1_23[185]},
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage2_26[30],stage2_25[56],stage2_24[59],stage2_23[64],stage2_22[98]}
   );
   gpc615_5 gpc6380 (
      {stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178]},
      {stage1_23[186]},
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage2_26[31],stage2_25[57],stage2_24[60],stage2_23[65],stage2_22[99]}
   );
   gpc615_5 gpc6381 (
      {stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182], stage1_22[183]},
      {stage1_23[187]},
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage2_26[32],stage2_25[58],stage2_24[61],stage2_23[66],stage2_22[100]}
   );
   gpc615_5 gpc6382 (
      {stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187], stage1_22[188]},
      {stage1_23[188]},
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage2_26[33],stage2_25[59],stage2_24[62],stage2_23[67],stage2_22[101]}
   );
   gpc615_5 gpc6383 (
      {stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192], stage1_22[193]},
      {stage1_23[189]},
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage2_26[34],stage2_25[60],stage2_24[63],stage2_23[68],stage2_22[102]}
   );
   gpc615_5 gpc6384 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[210]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[35],stage2_25[61],stage2_24[64],stage2_23[69]}
   );
   gpc615_5 gpc6385 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[211]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[36],stage2_25[62],stage2_24[65],stage2_23[70]}
   );
   gpc615_5 gpc6386 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[212]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[37],stage2_25[63],stage2_24[66],stage2_23[71]}
   );
   gpc615_5 gpc6387 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[213]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[38],stage2_25[64],stage2_24[67],stage2_23[72]}
   );
   gpc615_5 gpc6388 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[214]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[39],stage2_25[65],stage2_24[68],stage2_23[73]}
   );
   gpc615_5 gpc6389 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[215]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[40],stage2_25[66],stage2_24[69],stage2_23[74]}
   );
   gpc615_5 gpc6390 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[216]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[41],stage2_25[67],stage2_24[70],stage2_23[75]}
   );
   gpc615_5 gpc6391 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[217]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[42],stage2_25[68],stage2_24[71],stage2_23[76]}
   );
   gpc615_5 gpc6392 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[218]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[43],stage2_25[69],stage2_24[72],stage2_23[77]}
   );
   gpc615_5 gpc6393 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[219]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[44],stage2_25[70],stage2_24[73],stage2_23[78]}
   );
   gpc615_5 gpc6394 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[220]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[45],stage2_25[71],stage2_24[74],stage2_23[79]}
   );
   gpc615_5 gpc6395 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[221]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[46],stage2_25[72],stage2_24[75],stage2_23[80]}
   );
   gpc615_5 gpc6396 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[222]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[47],stage2_25[73],stage2_24[76],stage2_23[81]}
   );
   gpc615_5 gpc6397 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[223]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[48],stage2_25[74],stage2_24[77],stage2_23[82]}
   );
   gpc615_5 gpc6398 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[224]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[49],stage2_25[75],stage2_24[78],stage2_23[83]}
   );
   gpc615_5 gpc6399 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[225]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[50],stage2_25[76],stage2_24[79],stage2_23[84]}
   );
   gpc615_5 gpc6400 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[226]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[51],stage2_25[77],stage2_24[80],stage2_23[85]}
   );
   gpc615_5 gpc6401 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[227]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[52],stage2_25[78],stage2_24[81],stage2_23[86]}
   );
   gpc615_5 gpc6402 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[228]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[53],stage2_25[79],stage2_24[82],stage2_23[87]}
   );
   gpc615_5 gpc6403 (
      {stage1_23[285], stage1_23[286], stage1_23[287], stage1_23[288], stage1_23[289]},
      {stage1_24[229]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[54],stage2_25[80],stage2_24[83],stage2_23[88]}
   );
   gpc606_5 gpc6404 (
      {stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233], stage1_24[234], 1'b0},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[20],stage2_26[55],stage2_25[81],stage2_24[84]}
   );
   gpc606_5 gpc6405 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[1],stage2_27[21],stage2_26[56],stage2_25[82]}
   );
   gpc606_5 gpc6406 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[2],stage2_27[22],stage2_26[57],stage2_25[83]}
   );
   gpc606_5 gpc6407 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[3],stage2_27[23],stage2_26[58],stage2_25[84]}
   );
   gpc606_5 gpc6408 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[4],stage2_27[24],stage2_26[59],stage2_25[85]}
   );
   gpc606_5 gpc6409 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[5],stage2_27[25],stage2_26[60],stage2_25[86]}
   );
   gpc606_5 gpc6410 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[6],stage2_27[26],stage2_26[61],stage2_25[87]}
   );
   gpc606_5 gpc6411 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[7],stage2_27[27],stage2_26[62],stage2_25[88]}
   );
   gpc606_5 gpc6412 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[8],stage2_27[28],stage2_26[63],stage2_25[89]}
   );
   gpc606_5 gpc6413 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[9],stage2_27[29],stage2_26[64],stage2_25[90]}
   );
   gpc606_5 gpc6414 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[10],stage2_27[30],stage2_26[65],stage2_25[91]}
   );
   gpc615_5 gpc6415 (
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10]},
      {stage1_27[60]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[10],stage2_28[11],stage2_27[31],stage2_26[66]}
   );
   gpc615_5 gpc6416 (
      {stage1_26[11], stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15]},
      {stage1_27[61]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[11],stage2_28[12],stage2_27[32],stage2_26[67]}
   );
   gpc615_5 gpc6417 (
      {stage1_26[16], stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20]},
      {stage1_27[62]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[12],stage2_28[13],stage2_27[33],stage2_26[68]}
   );
   gpc615_5 gpc6418 (
      {stage1_26[21], stage1_26[22], stage1_26[23], stage1_26[24], stage1_26[25]},
      {stage1_27[63]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[13],stage2_28[14],stage2_27[34],stage2_26[69]}
   );
   gpc615_5 gpc6419 (
      {stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29], stage1_26[30]},
      {stage1_27[64]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[14],stage2_28[15],stage2_27[35],stage2_26[70]}
   );
   gpc615_5 gpc6420 (
      {stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[65]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[15],stage2_28[16],stage2_27[36],stage2_26[71]}
   );
   gpc615_5 gpc6421 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40]},
      {stage1_27[66]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[16],stage2_28[17],stage2_27[37],stage2_26[72]}
   );
   gpc615_5 gpc6422 (
      {stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45]},
      {stage1_27[67]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[17],stage2_28[18],stage2_27[38],stage2_26[73]}
   );
   gpc615_5 gpc6423 (
      {stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49], stage1_26[50]},
      {stage1_27[68]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[18],stage2_28[19],stage2_27[39],stage2_26[74]}
   );
   gpc615_5 gpc6424 (
      {stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54], stage1_26[55]},
      {stage1_27[69]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[19],stage2_28[20],stage2_27[40],stage2_26[75]}
   );
   gpc615_5 gpc6425 (
      {stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59], stage1_26[60]},
      {stage1_27[70]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[20],stage2_28[21],stage2_27[41],stage2_26[76]}
   );
   gpc615_5 gpc6426 (
      {stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage1_27[71]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[21],stage2_28[22],stage2_27[42],stage2_26[77]}
   );
   gpc615_5 gpc6427 (
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70]},
      {stage1_27[72]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[22],stage2_28[23],stage2_27[43],stage2_26[78]}
   );
   gpc615_5 gpc6428 (
      {stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75]},
      {stage1_27[73]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[23],stage2_28[24],stage2_27[44],stage2_26[79]}
   );
   gpc615_5 gpc6429 (
      {stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79], stage1_26[80]},
      {stage1_27[74]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[24],stage2_28[25],stage2_27[45],stage2_26[80]}
   );
   gpc615_5 gpc6430 (
      {stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84], stage1_26[85]},
      {stage1_27[75]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[25],stage2_28[26],stage2_27[46],stage2_26[81]}
   );
   gpc615_5 gpc6431 (
      {stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89], stage1_26[90]},
      {stage1_27[76]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[26],stage2_28[27],stage2_27[47],stage2_26[82]}
   );
   gpc615_5 gpc6432 (
      {stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage1_27[77]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[27],stage2_28[28],stage2_27[48],stage2_26[83]}
   );
   gpc615_5 gpc6433 (
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100]},
      {stage1_27[78]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[28],stage2_28[29],stage2_27[49],stage2_26[84]}
   );
   gpc615_5 gpc6434 (
      {stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105]},
      {stage1_27[79]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[29],stage2_28[30],stage2_27[50],stage2_26[85]}
   );
   gpc615_5 gpc6435 (
      {stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109], stage1_26[110]},
      {stage1_27[80]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[30],stage2_28[31],stage2_27[51],stage2_26[86]}
   );
   gpc615_5 gpc6436 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[81]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[31],stage2_28[32],stage2_27[52],stage2_26[87]}
   );
   gpc615_5 gpc6437 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[82]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[32],stage2_28[33],stage2_27[53],stage2_26[88]}
   );
   gpc615_5 gpc6438 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[83]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[33],stage2_28[34],stage2_27[54],stage2_26[89]}
   );
   gpc615_5 gpc6439 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[84]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[34],stage2_28[35],stage2_27[55],stage2_26[90]}
   );
   gpc615_5 gpc6440 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[85]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[35],stage2_28[36],stage2_27[56],stage2_26[91]}
   );
   gpc615_5 gpc6441 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[86]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[36],stage2_28[37],stage2_27[57],stage2_26[92]}
   );
   gpc615_5 gpc6442 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[87]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[37],stage2_28[38],stage2_27[58],stage2_26[93]}
   );
   gpc615_5 gpc6443 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[88]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[38],stage2_28[39],stage2_27[59],stage2_26[94]}
   );
   gpc623_5 gpc6444 (
      {stage1_26[151], stage1_26[152], stage1_26[153]},
      {stage1_27[89], stage1_27[90]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[39],stage2_28[40],stage2_27[60],stage2_26[95]}
   );
   gpc615_5 gpc6445 (
      {stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage1_28[180]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[30],stage2_29[40],stage2_28[41],stage2_27[61]}
   );
   gpc615_5 gpc6446 (
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100]},
      {stage1_28[181]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[31],stage2_29[41],stage2_28[42],stage2_27[62]}
   );
   gpc615_5 gpc6447 (
      {stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105]},
      {stage1_28[182]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[32],stage2_29[42],stage2_28[43],stage2_27[63]}
   );
   gpc615_5 gpc6448 (
      {stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109], stage1_27[110]},
      {stage1_28[183]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[33],stage2_29[43],stage2_28[44],stage2_27[64]}
   );
   gpc615_5 gpc6449 (
      {stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114], stage1_27[115]},
      {stage1_28[184]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[34],stage2_29[44],stage2_28[45],stage2_27[65]}
   );
   gpc615_5 gpc6450 (
      {stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119], stage1_27[120]},
      {stage1_28[185]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[35],stage2_29[45],stage2_28[46],stage2_27[66]}
   );
   gpc615_5 gpc6451 (
      {stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage1_28[186]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[36],stage2_29[46],stage2_28[47],stage2_27[67]}
   );
   gpc615_5 gpc6452 (
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130]},
      {stage1_28[187]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[37],stage2_29[47],stage2_28[48],stage2_27[68]}
   );
   gpc615_5 gpc6453 (
      {stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135]},
      {stage1_28[188]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[38],stage2_29[48],stage2_28[49],stage2_27[69]}
   );
   gpc615_5 gpc6454 (
      {stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139], stage1_27[140]},
      {stage1_28[189]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[39],stage2_29[49],stage2_28[50],stage2_27[70]}
   );
   gpc615_5 gpc6455 (
      {stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144], stage1_27[145]},
      {stage1_28[190]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[40],stage2_29[50],stage2_28[51],stage2_27[71]}
   );
   gpc615_5 gpc6456 (
      {stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149], stage1_27[150]},
      {stage1_28[191]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[41],stage2_29[51],stage2_28[52],stage2_27[72]}
   );
   gpc615_5 gpc6457 (
      {stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage1_28[192]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[42],stage2_29[52],stage2_28[53],stage2_27[73]}
   );
   gpc615_5 gpc6458 (
      {stage1_27[156], stage1_27[157], stage1_27[158], stage1_27[159], stage1_27[160]},
      {stage1_28[193]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[43],stage2_29[53],stage2_28[54],stage2_27[74]}
   );
   gpc615_5 gpc6459 (
      {stage1_27[161], stage1_27[162], stage1_27[163], stage1_27[164], stage1_27[165]},
      {stage1_28[194]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[44],stage2_29[54],stage2_28[55],stage2_27[75]}
   );
   gpc615_5 gpc6460 (
      {stage1_27[166], stage1_27[167], stage1_27[168], stage1_27[169], stage1_27[170]},
      {stage1_28[195]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[45],stage2_29[55],stage2_28[56],stage2_27[76]}
   );
   gpc615_5 gpc6461 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[196]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[46],stage2_29[56],stage2_28[57],stage2_27[77]}
   );
   gpc615_5 gpc6462 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[197]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[47],stage2_29[57],stage2_28[58],stage2_27[78]}
   );
   gpc615_5 gpc6463 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[198]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[48],stage2_29[58],stage2_28[59],stage2_27[79]}
   );
   gpc615_5 gpc6464 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[199]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[49],stage2_29[59],stage2_28[60],stage2_27[80]}
   );
   gpc615_5 gpc6465 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[200]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[50],stage2_29[60],stage2_28[61],stage2_27[81]}
   );
   gpc615_5 gpc6466 (
      {stage1_27[196], stage1_27[197], stage1_27[198], stage1_27[199], stage1_27[200]},
      {stage1_28[201]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[51],stage2_29[61],stage2_28[62],stage2_27[82]}
   );
   gpc615_5 gpc6467 (
      {stage1_27[201], stage1_27[202], stage1_27[203], stage1_27[204], stage1_27[205]},
      {stage1_28[202]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[52],stage2_29[62],stage2_28[63],stage2_27[83]}
   );
   gpc615_5 gpc6468 (
      {stage1_27[206], stage1_27[207], stage1_27[208], stage1_27[209], stage1_27[210]},
      {stage1_28[203]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[53],stage2_29[63],stage2_28[64],stage2_27[84]}
   );
   gpc606_5 gpc6469 (
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[24],stage2_30[54],stage2_29[64],stage2_28[65]}
   );
   gpc606_5 gpc6470 (
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[25],stage2_30[55],stage2_29[65],stage2_28[66]}
   );
   gpc606_5 gpc6471 (
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[26],stage2_30[56],stage2_29[66],stage2_28[67]}
   );
   gpc606_5 gpc6472 (
      {stage1_28[222], stage1_28[223], stage1_28[224], stage1_28[225], stage1_28[226], stage1_28[227]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[27],stage2_30[57],stage2_29[67],stage2_28[68]}
   );
   gpc606_5 gpc6473 (
      {stage1_28[228], stage1_28[229], stage1_28[230], stage1_28[231], stage1_28[232], stage1_28[233]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[28],stage2_30[58],stage2_29[68],stage2_28[69]}
   );
   gpc606_5 gpc6474 (
      {stage1_28[234], stage1_28[235], stage1_28[236], stage1_28[237], stage1_28[238], stage1_28[239]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[29],stage2_30[59],stage2_29[69],stage2_28[70]}
   );
   gpc606_5 gpc6475 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[6],stage2_31[30],stage2_30[60],stage2_29[70]}
   );
   gpc606_5 gpc6476 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[7],stage2_31[31],stage2_30[61],stage2_29[71]}
   );
   gpc606_5 gpc6477 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[8],stage2_31[32],stage2_30[62],stage2_29[72]}
   );
   gpc606_5 gpc6478 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[9],stage2_31[33],stage2_30[63],stage2_29[73]}
   );
   gpc606_5 gpc6479 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[10],stage2_31[34],stage2_30[64],stage2_29[74]}
   );
   gpc606_5 gpc6480 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[11],stage2_31[35],stage2_30[65],stage2_29[75]}
   );
   gpc606_5 gpc6481 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[12],stage2_31[36],stage2_30[66],stage2_29[76]}
   );
   gpc2135_5 gpc6482 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40]},
      {stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_32[0]},
      {stage1_33[0], stage1_33[1]},
      {stage2_34[0],stage2_33[7],stage2_32[13],stage2_31[37],stage2_30[67]}
   );
   gpc207_4 gpc6483 (
      {stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[1], stage1_32[2]},
      {stage2_33[8],stage2_32[14],stage2_31[38],stage2_30[68]}
   );
   gpc207_4 gpc6484 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_32[3], stage1_32[4]},
      {stage2_33[9],stage2_32[15],stage2_31[39],stage2_30[69]}
   );
   gpc207_4 gpc6485 (
      {stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_32[5], stage1_32[6]},
      {stage2_33[10],stage2_32[16],stage2_31[40],stage2_30[70]}
   );
   gpc207_4 gpc6486 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66], stage1_30[67], stage1_30[68]},
      {stage1_32[7], stage1_32[8]},
      {stage2_33[11],stage2_32[17],stage2_31[41],stage2_30[71]}
   );
   gpc207_4 gpc6487 (
      {stage1_30[69], stage1_30[70], stage1_30[71], stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75]},
      {stage1_32[9], stage1_32[10]},
      {stage2_33[12],stage2_32[18],stage2_31[42],stage2_30[72]}
   );
   gpc606_5 gpc6488 (
      {stage1_30[76], stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16]},
      {stage2_34[1],stage2_33[13],stage2_32[19],stage2_31[43],stage2_30[73]}
   );
   gpc606_5 gpc6489 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87]},
      {stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22]},
      {stage2_34[2],stage2_33[14],stage2_32[20],stage2_31[44],stage2_30[74]}
   );
   gpc606_5 gpc6490 (
      {stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93]},
      {stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28]},
      {stage2_34[3],stage2_33[15],stage2_32[21],stage2_31[45],stage2_30[75]}
   );
   gpc606_5 gpc6491 (
      {stage1_30[94], stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34]},
      {stage2_34[4],stage2_33[16],stage2_32[22],stage2_31[46],stage2_30[76]}
   );
   gpc606_5 gpc6492 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105]},
      {stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40]},
      {stage2_34[5],stage2_33[17],stage2_32[23],stage2_31[47],stage2_30[77]}
   );
   gpc606_5 gpc6493 (
      {stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111]},
      {stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46]},
      {stage2_34[6],stage2_33[18],stage2_32[24],stage2_31[48],stage2_30[78]}
   );
   gpc606_5 gpc6494 (
      {stage1_30[112], stage1_30[113], stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117]},
      {stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52]},
      {stage2_34[7],stage2_33[19],stage2_32[25],stage2_31[49],stage2_30[79]}
   );
   gpc606_5 gpc6495 (
      {stage1_30[118], stage1_30[119], stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123]},
      {stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58]},
      {stage2_34[8],stage2_33[20],stage2_32[26],stage2_31[50],stage2_30[80]}
   );
   gpc606_5 gpc6496 (
      {stage1_30[124], stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64]},
      {stage2_34[9],stage2_33[21],stage2_32[27],stage2_31[51],stage2_30[81]}
   );
   gpc606_5 gpc6497 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135]},
      {stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70]},
      {stage2_34[10],stage2_33[22],stage2_32[28],stage2_31[52],stage2_30[82]}
   );
   gpc606_5 gpc6498 (
      {stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141]},
      {stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76]},
      {stage2_34[11],stage2_33[23],stage2_32[29],stage2_31[53],stage2_30[83]}
   );
   gpc606_5 gpc6499 (
      {stage1_30[142], stage1_30[143], stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147]},
      {stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82]},
      {stage2_34[12],stage2_33[24],stage2_32[30],stage2_31[54],stage2_30[84]}
   );
   gpc606_5 gpc6500 (
      {stage1_30[148], stage1_30[149], stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153]},
      {stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88]},
      {stage2_34[13],stage2_33[25],stage2_32[31],stage2_31[55],stage2_30[85]}
   );
   gpc606_5 gpc6501 (
      {stage1_30[154], stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94]},
      {stage2_34[14],stage2_33[26],stage2_32[32],stage2_31[56],stage2_30[86]}
   );
   gpc606_5 gpc6502 (
      {stage1_30[160], stage1_30[161], stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165]},
      {stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100]},
      {stage2_34[15],stage2_33[27],stage2_32[33],stage2_31[57],stage2_30[87]}
   );
   gpc606_5 gpc6503 (
      {stage1_30[166], stage1_30[167], stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171]},
      {stage1_32[101], stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106]},
      {stage2_34[16],stage2_33[28],stage2_32[34],stage2_31[58],stage2_30[88]}
   );
   gpc606_5 gpc6504 (
      {stage1_30[172], stage1_30[173], stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177]},
      {stage1_32[107], stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112]},
      {stage2_34[17],stage2_33[29],stage2_32[35],stage2_31[59],stage2_30[89]}
   );
   gpc606_5 gpc6505 (
      {stage1_30[178], stage1_30[179], stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183]},
      {stage1_32[113], stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118]},
      {stage2_34[18],stage2_33[30],stage2_32[36],stage2_31[60],stage2_30[90]}
   );
   gpc606_5 gpc6506 (
      {stage1_30[184], stage1_30[185], stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189]},
      {stage1_32[119], stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124]},
      {stage2_34[19],stage2_33[31],stage2_32[37],stage2_31[61],stage2_30[91]}
   );
   gpc606_5 gpc6507 (
      {stage1_30[190], stage1_30[191], stage1_30[192], stage1_30[193], stage1_30[194], stage1_30[195]},
      {stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130]},
      {stage2_34[20],stage2_33[32],stage2_32[38],stage2_31[62],stage2_30[92]}
   );
   gpc606_5 gpc6508 (
      {stage1_30[196], stage1_30[197], stage1_30[198], stage1_30[199], stage1_30[200], stage1_30[201]},
      {stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136]},
      {stage2_34[21],stage2_33[33],stage2_32[39],stage2_31[63],stage2_30[93]}
   );
   gpc606_5 gpc6509 (
      {stage1_30[202], stage1_30[203], stage1_30[204], stage1_30[205], stage1_30[206], stage1_30[207]},
      {stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140], stage1_32[141], stage1_32[142]},
      {stage2_34[22],stage2_33[34],stage2_32[40],stage2_31[64],stage2_30[94]}
   );
   gpc606_5 gpc6510 (
      {stage1_30[208], stage1_30[209], stage1_30[210], stage1_30[211], stage1_30[212], stage1_30[213]},
      {stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146], stage1_32[147], stage1_32[148]},
      {stage2_34[23],stage2_33[35],stage2_32[41],stage2_31[65],stage2_30[95]}
   );
   gpc606_5 gpc6511 (
      {stage1_30[214], stage1_30[215], stage1_30[216], stage1_30[217], stage1_30[218], stage1_30[219]},
      {stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152], stage1_32[153], stage1_32[154]},
      {stage2_34[24],stage2_33[36],stage2_32[42],stage2_31[66],stage2_30[96]}
   );
   gpc606_5 gpc6512 (
      {stage1_30[220], stage1_30[221], stage1_30[222], stage1_30[223], stage1_30[224], stage1_30[225]},
      {stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158], stage1_32[159], stage1_32[160]},
      {stage2_34[25],stage2_33[37],stage2_32[43],stage2_31[67],stage2_30[97]}
   );
   gpc606_5 gpc6513 (
      {stage1_30[226], stage1_30[227], stage1_30[228], stage1_30[229], stage1_30[230], stage1_30[231]},
      {stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164], stage1_32[165], stage1_32[166]},
      {stage2_34[26],stage2_33[38],stage2_32[44],stage2_31[68],stage2_30[98]}
   );
   gpc615_5 gpc6514 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49]},
      {stage1_32[167]},
      {stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6], stage1_33[7]},
      {stage2_35[0],stage2_34[27],stage2_33[39],stage2_32[45],stage2_31[69]}
   );
   gpc615_5 gpc6515 (
      {stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54]},
      {stage1_32[168]},
      {stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12], stage1_33[13]},
      {stage2_35[1],stage2_34[28],stage2_33[40],stage2_32[46],stage2_31[70]}
   );
   gpc615_5 gpc6516 (
      {stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage1_32[169]},
      {stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18], stage1_33[19]},
      {stage2_35[2],stage2_34[29],stage2_33[41],stage2_32[47],stage2_31[71]}
   );
   gpc615_5 gpc6517 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64]},
      {stage1_32[170]},
      {stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24], stage1_33[25]},
      {stage2_35[3],stage2_34[30],stage2_33[42],stage2_32[48],stage2_31[72]}
   );
   gpc615_5 gpc6518 (
      {stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69]},
      {stage1_32[171]},
      {stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30], stage1_33[31]},
      {stage2_35[4],stage2_34[31],stage2_33[43],stage2_32[49],stage2_31[73]}
   );
   gpc615_5 gpc6519 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[172]},
      {stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36], stage1_33[37]},
      {stage2_35[5],stage2_34[32],stage2_33[44],stage2_32[50],stage2_31[74]}
   );
   gpc615_5 gpc6520 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79]},
      {stage1_32[173]},
      {stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42], stage1_33[43]},
      {stage2_35[6],stage2_34[33],stage2_33[45],stage2_32[51],stage2_31[75]}
   );
   gpc615_5 gpc6521 (
      {stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84]},
      {stage1_32[174]},
      {stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48], stage1_33[49]},
      {stage2_35[7],stage2_34[34],stage2_33[46],stage2_32[52],stage2_31[76]}
   );
   gpc615_5 gpc6522 (
      {stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_32[175]},
      {stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54], stage1_33[55]},
      {stage2_35[8],stage2_34[35],stage2_33[47],stage2_32[53],stage2_31[77]}
   );
   gpc615_5 gpc6523 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94]},
      {stage1_32[176]},
      {stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60], stage1_33[61]},
      {stage2_35[9],stage2_34[36],stage2_33[48],stage2_32[54],stage2_31[78]}
   );
   gpc615_5 gpc6524 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99]},
      {stage1_32[177]},
      {stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66], stage1_33[67]},
      {stage2_35[10],stage2_34[37],stage2_33[49],stage2_32[55],stage2_31[79]}
   );
   gpc615_5 gpc6525 (
      {stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_32[178]},
      {stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72], stage1_33[73]},
      {stage2_35[11],stage2_34[38],stage2_33[50],stage2_32[56],stage2_31[80]}
   );
   gpc615_5 gpc6526 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[179]},
      {stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78], stage1_33[79]},
      {stage2_35[12],stage2_34[39],stage2_33[51],stage2_32[57],stage2_31[81]}
   );
   gpc615_5 gpc6527 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[180]},
      {stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84], stage1_33[85]},
      {stage2_35[13],stage2_34[40],stage2_33[52],stage2_32[58],stage2_31[82]}
   );
   gpc615_5 gpc6528 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[181]},
      {stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90], stage1_33[91]},
      {stage2_35[14],stage2_34[41],stage2_33[53],stage2_32[59],stage2_31[83]}
   );
   gpc615_5 gpc6529 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[182]},
      {stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96], stage1_33[97]},
      {stage2_35[15],stage2_34[42],stage2_33[54],stage2_32[60],stage2_31[84]}
   );
   gpc615_5 gpc6530 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[183]},
      {stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102], stage1_33[103]},
      {stage2_35[16],stage2_34[43],stage2_33[55],stage2_32[61],stage2_31[85]}
   );
   gpc615_5 gpc6531 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[184]},
      {stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108], stage1_33[109]},
      {stage2_35[17],stage2_34[44],stage2_33[56],stage2_32[62],stage2_31[86]}
   );
   gpc615_5 gpc6532 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[185]},
      {stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114], stage1_33[115]},
      {stage2_35[18],stage2_34[45],stage2_33[57],stage2_32[63],stage2_31[87]}
   );
   gpc615_5 gpc6533 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[186]},
      {stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120], stage1_33[121]},
      {stage2_35[19],stage2_34[46],stage2_33[58],stage2_32[64],stage2_31[88]}
   );
   gpc615_5 gpc6534 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[187]},
      {stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126], stage1_33[127]},
      {stage2_35[20],stage2_34[47],stage2_33[59],stage2_32[65],stage2_31[89]}
   );
   gpc615_5 gpc6535 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[188]},
      {stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132], stage1_33[133]},
      {stage2_35[21],stage2_34[48],stage2_33[60],stage2_32[66],stage2_31[90]}
   );
   gpc615_5 gpc6536 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[189]},
      {stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138], stage1_33[139]},
      {stage2_35[22],stage2_34[49],stage2_33[61],stage2_32[67],stage2_31[91]}
   );
   gpc615_5 gpc6537 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[190]},
      {stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144], stage1_33[145]},
      {stage2_35[23],stage2_34[50],stage2_33[62],stage2_32[68],stage2_31[92]}
   );
   gpc615_5 gpc6538 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[191]},
      {stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150], stage1_33[151]},
      {stage2_35[24],stage2_34[51],stage2_33[63],stage2_32[69],stage2_31[93]}
   );
   gpc615_5 gpc6539 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[192]},
      {stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156], stage1_33[157]},
      {stage2_35[25],stage2_34[52],stage2_33[64],stage2_32[70],stage2_31[94]}
   );
   gpc615_5 gpc6540 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[193]},
      {stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162], stage1_33[163]},
      {stage2_35[26],stage2_34[53],stage2_33[65],stage2_32[71],stage2_31[95]}
   );
   gpc606_5 gpc6541 (
      {stage1_32[194], stage1_32[195], stage1_32[196], stage1_32[197], stage1_32[198], stage1_32[199]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[27],stage2_34[54],stage2_33[66],stage2_32[72]}
   );
   gpc606_5 gpc6542 (
      {stage1_32[200], stage1_32[201], stage1_32[202], stage1_32[203], stage1_32[204], stage1_32[205]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[28],stage2_34[55],stage2_33[67],stage2_32[73]}
   );
   gpc606_5 gpc6543 (
      {stage1_32[206], stage1_32[207], stage1_32[208], stage1_32[209], stage1_32[210], stage1_32[211]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[29],stage2_34[56],stage2_33[68],stage2_32[74]}
   );
   gpc606_5 gpc6544 (
      {stage1_32[212], stage1_32[213], stage1_32[214], stage1_32[215], stage1_32[216], stage1_32[217]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[30],stage2_34[57],stage2_33[69],stage2_32[75]}
   );
   gpc606_5 gpc6545 (
      {stage1_32[218], stage1_32[219], stage1_32[220], stage1_32[221], stage1_32[222], stage1_32[223]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[31],stage2_34[58],stage2_33[70],stage2_32[76]}
   );
   gpc606_5 gpc6546 (
      {stage1_32[224], stage1_32[225], stage1_32[226], stage1_32[227], stage1_32[228], stage1_32[229]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[32],stage2_34[59],stage2_33[71],stage2_32[77]}
   );
   gpc606_5 gpc6547 (
      {stage1_32[230], stage1_32[231], stage1_32[232], stage1_32[233], stage1_32[234], stage1_32[235]},
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage2_36[6],stage2_35[33],stage2_34[60],stage2_33[72],stage2_32[78]}
   );
   gpc606_5 gpc6548 (
      {stage1_32[236], stage1_32[237], stage1_32[238], stage1_32[239], stage1_32[240], stage1_32[241]},
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage2_36[7],stage2_35[34],stage2_34[61],stage2_33[73],stage2_32[79]}
   );
   gpc606_5 gpc6549 (
      {stage1_32[242], stage1_32[243], stage1_32[244], stage1_32[245], stage1_32[246], stage1_32[247]},
      {stage1_34[48], stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53]},
      {stage2_36[8],stage2_35[35],stage2_34[62],stage2_33[74],stage2_32[80]}
   );
   gpc606_5 gpc6550 (
      {stage1_32[248], stage1_32[249], stage1_32[250], stage1_32[251], stage1_32[252], stage1_32[253]},
      {stage1_34[54], stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59]},
      {stage2_36[9],stage2_35[36],stage2_34[63],stage2_33[75],stage2_32[81]}
   );
   gpc606_5 gpc6551 (
      {stage1_32[254], stage1_32[255], stage1_32[256], stage1_32[257], stage1_32[258], stage1_32[259]},
      {stage1_34[60], stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage2_36[10],stage2_35[37],stage2_34[64],stage2_33[76],stage2_32[82]}
   );
   gpc606_5 gpc6552 (
      {stage1_32[260], stage1_32[261], stage1_32[262], stage1_32[263], stage1_32[264], stage1_32[265]},
      {stage1_34[66], stage1_34[67], stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71]},
      {stage2_36[11],stage2_35[38],stage2_34[65],stage2_33[77],stage2_32[83]}
   );
   gpc606_5 gpc6553 (
      {stage1_32[266], stage1_32[267], stage1_32[268], stage1_32[269], stage1_32[270], stage1_32[271]},
      {stage1_34[72], stage1_34[73], stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77]},
      {stage2_36[12],stage2_35[39],stage2_34[66],stage2_33[78],stage2_32[84]}
   );
   gpc606_5 gpc6554 (
      {stage1_32[272], stage1_32[273], stage1_32[274], stage1_32[275], stage1_32[276], stage1_32[277]},
      {stage1_34[78], stage1_34[79], stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83]},
      {stage2_36[13],stage2_35[40],stage2_34[67],stage2_33[79],stage2_32[85]}
   );
   gpc606_5 gpc6555 (
      {stage1_32[278], stage1_32[279], stage1_32[280], stage1_32[281], stage1_32[282], stage1_32[283]},
      {stage1_34[84], stage1_34[85], stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89]},
      {stage2_36[14],stage2_35[41],stage2_34[68],stage2_33[80],stage2_32[86]}
   );
   gpc606_5 gpc6556 (
      {stage1_32[284], stage1_32[285], stage1_32[286], stage1_32[287], stage1_32[288], stage1_32[289]},
      {stage1_34[90], stage1_34[91], stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95]},
      {stage2_36[15],stage2_35[42],stage2_34[69],stage2_33[81],stage2_32[87]}
   );
   gpc606_5 gpc6557 (
      {stage1_32[290], stage1_32[291], stage1_32[292], stage1_32[293], stage1_32[294], stage1_32[295]},
      {stage1_34[96], stage1_34[97], stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101]},
      {stage2_36[16],stage2_35[43],stage2_34[70],stage2_33[82],stage2_32[88]}
   );
   gpc606_5 gpc6558 (
      {stage1_32[296], stage1_32[297], stage1_32[298], stage1_32[299], stage1_32[300], stage1_32[301]},
      {stage1_34[102], stage1_34[103], stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107]},
      {stage2_36[17],stage2_35[44],stage2_34[71],stage2_33[83],stage2_32[89]}
   );
   gpc606_5 gpc6559 (
      {stage1_32[302], stage1_32[303], stage1_32[304], stage1_32[305], stage1_32[306], stage1_32[307]},
      {stage1_34[108], stage1_34[109], stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113]},
      {stage2_36[18],stage2_35[45],stage2_34[72],stage2_33[84],stage2_32[90]}
   );
   gpc606_5 gpc6560 (
      {stage1_32[308], stage1_32[309], stage1_32[310], stage1_32[311], stage1_32[312], stage1_32[313]},
      {stage1_34[114], stage1_34[115], stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119]},
      {stage2_36[19],stage2_35[46],stage2_34[73],stage2_33[85],stage2_32[91]}
   );
   gpc606_5 gpc6561 (
      {stage1_32[314], stage1_32[315], stage1_32[316], stage1_32[317], stage1_32[318], stage1_32[319]},
      {stage1_34[120], stage1_34[121], stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125]},
      {stage2_36[20],stage2_35[47],stage2_34[74],stage2_33[86],stage2_32[92]}
   );
   gpc606_5 gpc6562 (
      {stage1_32[320], stage1_32[321], stage1_32[322], stage1_32[323], stage1_32[324], stage1_32[325]},
      {stage1_34[126], stage1_34[127], stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131]},
      {stage2_36[21],stage2_35[48],stage2_34[75],stage2_33[87],stage2_32[93]}
   );
   gpc606_5 gpc6563 (
      {stage1_32[326], stage1_32[327], stage1_32[328], stage1_32[329], stage1_32[330], stage1_32[331]},
      {stage1_34[132], stage1_34[133], stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137]},
      {stage2_36[22],stage2_35[49],stage2_34[76],stage2_33[88],stage2_32[94]}
   );
   gpc606_5 gpc6564 (
      {stage1_32[332], stage1_32[333], stage1_32[334], stage1_32[335], stage1_32[336], stage1_32[337]},
      {stage1_34[138], stage1_34[139], stage1_34[140], stage1_34[141], stage1_34[142], stage1_34[143]},
      {stage2_36[23],stage2_35[50],stage2_34[77],stage2_33[89],stage2_32[95]}
   );
   gpc606_5 gpc6565 (
      {stage1_32[338], stage1_32[339], stage1_32[340], stage1_32[341], stage1_32[342], stage1_32[343]},
      {stage1_34[144], stage1_34[145], stage1_34[146], stage1_34[147], stage1_34[148], stage1_34[149]},
      {stage2_36[24],stage2_35[51],stage2_34[78],stage2_33[90],stage2_32[96]}
   );
   gpc606_5 gpc6566 (
      {stage1_32[344], stage1_32[345], stage1_32[346], stage1_32[347], stage1_32[348], stage1_32[349]},
      {stage1_34[150], stage1_34[151], stage1_34[152], stage1_34[153], stage1_34[154], stage1_34[155]},
      {stage2_36[25],stage2_35[52],stage2_34[79],stage2_33[91],stage2_32[97]}
   );
   gpc606_5 gpc6567 (
      {stage1_32[350], stage1_32[351], stage1_32[352], stage1_32[353], stage1_32[354], stage1_32[355]},
      {stage1_34[156], stage1_34[157], stage1_34[158], stage1_34[159], stage1_34[160], stage1_34[161]},
      {stage2_36[26],stage2_35[53],stage2_34[80],stage2_33[92],stage2_32[98]}
   );
   gpc606_5 gpc6568 (
      {stage1_32[356], stage1_32[357], stage1_32[358], stage1_32[359], stage1_32[360], stage1_32[361]},
      {stage1_34[162], stage1_34[163], stage1_34[164], stage1_34[165], stage1_34[166], stage1_34[167]},
      {stage2_36[27],stage2_35[54],stage2_34[81],stage2_33[93],stage2_32[99]}
   );
   gpc606_5 gpc6569 (
      {stage1_32[362], stage1_32[363], stage1_32[364], stage1_32[365], stage1_32[366], stage1_32[367]},
      {stage1_34[168], stage1_34[169], stage1_34[170], stage1_34[171], stage1_34[172], stage1_34[173]},
      {stage2_36[28],stage2_35[55],stage2_34[82],stage2_33[94],stage2_32[100]}
   );
   gpc606_5 gpc6570 (
      {stage1_32[368], stage1_32[369], stage1_32[370], stage1_32[371], stage1_32[372], stage1_32[373]},
      {stage1_34[174], stage1_34[175], stage1_34[176], stage1_34[177], stage1_34[178], stage1_34[179]},
      {stage2_36[29],stage2_35[56],stage2_34[83],stage2_33[95],stage2_32[101]}
   );
   gpc606_5 gpc6571 (
      {stage1_32[374], stage1_32[375], stage1_32[376], stage1_32[377], stage1_32[378], stage1_32[379]},
      {stage1_34[180], stage1_34[181], stage1_34[182], stage1_34[183], stage1_34[184], stage1_34[185]},
      {stage2_36[30],stage2_35[57],stage2_34[84],stage2_33[96],stage2_32[102]}
   );
   gpc606_5 gpc6572 (
      {stage1_32[380], stage1_32[381], stage1_32[382], stage1_32[383], stage1_32[384], stage1_32[385]},
      {stage1_34[186], stage1_34[187], stage1_34[188], stage1_34[189], stage1_34[190], stage1_34[191]},
      {stage2_36[31],stage2_35[58],stage2_34[85],stage2_33[97],stage2_32[103]}
   );
   gpc606_5 gpc6573 (
      {stage1_32[386], stage1_32[387], stage1_32[388], stage1_32[389], stage1_32[390], stage1_32[391]},
      {stage1_34[192], stage1_34[193], stage1_34[194], stage1_34[195], stage1_34[196], stage1_34[197]},
      {stage2_36[32],stage2_35[59],stage2_34[86],stage2_33[98],stage2_32[104]}
   );
   gpc606_5 gpc6574 (
      {stage1_32[392], stage1_32[393], stage1_32[394], stage1_32[395], stage1_32[396], stage1_32[397]},
      {stage1_34[198], stage1_34[199], stage1_34[200], stage1_34[201], stage1_34[202], stage1_34[203]},
      {stage2_36[33],stage2_35[60],stage2_34[87],stage2_33[99],stage2_32[105]}
   );
   gpc606_5 gpc6575 (
      {stage1_32[398], stage1_32[399], stage1_32[400], stage1_32[401], stage1_32[402], stage1_32[403]},
      {stage1_34[204], stage1_34[205], stage1_34[206], stage1_34[207], stage1_34[208], stage1_34[209]},
      {stage2_36[34],stage2_35[61],stage2_34[88],stage2_33[100],stage2_32[106]}
   );
   gpc606_5 gpc6576 (
      {stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168], stage1_33[169]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[35],stage2_35[62],stage2_34[89],stage2_33[101]}
   );
   gpc606_5 gpc6577 (
      {stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174], stage1_33[175]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[36],stage2_35[63],stage2_34[90],stage2_33[102]}
   );
   gpc606_5 gpc6578 (
      {stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180], stage1_33[181]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[37],stage2_35[64],stage2_34[91],stage2_33[103]}
   );
   gpc606_5 gpc6579 (
      {stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186], stage1_33[187]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[38],stage2_35[65],stage2_34[92],stage2_33[104]}
   );
   gpc606_5 gpc6580 (
      {stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192], stage1_33[193]},
      {stage1_35[24], stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29]},
      {stage2_37[4],stage2_36[39],stage2_35[66],stage2_34[93],stage2_33[105]}
   );
   gpc606_5 gpc6581 (
      {stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198], stage1_33[199]},
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage2_37[5],stage2_36[40],stage2_35[67],stage2_34[94],stage2_33[106]}
   );
   gpc615_5 gpc6582 (
      {stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage1_34[210]},
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage2_37[6],stage2_36[41],stage2_35[68],stage2_34[95],stage2_33[107]}
   );
   gpc615_5 gpc6583 (
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209]},
      {stage1_34[211]},
      {stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage2_37[7],stage2_36[42],stage2_35[69],stage2_34[96],stage2_33[108]}
   );
   gpc606_5 gpc6584 (
      {stage1_34[212], stage1_34[213], stage1_34[214], stage1_34[215], stage1_34[216], stage1_34[217]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[8],stage2_36[43],stage2_35[70],stage2_34[97]}
   );
   gpc606_5 gpc6585 (
      {stage1_34[218], stage1_34[219], stage1_34[220], stage1_34[221], stage1_34[222], stage1_34[223]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[9],stage2_36[44],stage2_35[71],stage2_34[98]}
   );
   gpc606_5 gpc6586 (
      {stage1_34[224], stage1_34[225], stage1_34[226], stage1_34[227], stage1_34[228], stage1_34[229]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[10],stage2_36[45],stage2_35[72],stage2_34[99]}
   );
   gpc606_5 gpc6587 (
      {stage1_34[230], stage1_34[231], stage1_34[232], stage1_34[233], stage1_34[234], stage1_34[235]},
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23]},
      {stage2_38[3],stage2_37[11],stage2_36[46],stage2_35[73],stage2_34[100]}
   );
   gpc606_5 gpc6588 (
      {stage1_34[236], stage1_34[237], stage1_34[238], stage1_34[239], stage1_34[240], stage1_34[241]},
      {stage1_36[24], stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29]},
      {stage2_38[4],stage2_37[12],stage2_36[47],stage2_35[74],stage2_34[101]}
   );
   gpc615_5 gpc6589 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[30]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[5],stage2_37[13],stage2_36[48],stage2_35[75]}
   );
   gpc615_5 gpc6590 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[31]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[6],stage2_37[14],stage2_36[49],stage2_35[76]}
   );
   gpc615_5 gpc6591 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[32]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[7],stage2_37[15],stage2_36[50],stage2_35[77]}
   );
   gpc615_5 gpc6592 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[33]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[8],stage2_37[16],stage2_36[51],stage2_35[78]}
   );
   gpc615_5 gpc6593 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[34]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[9],stage2_37[17],stage2_36[52],stage2_35[79]}
   );
   gpc615_5 gpc6594 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[35]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[10],stage2_37[18],stage2_36[53],stage2_35[80]}
   );
   gpc615_5 gpc6595 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[36]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[11],stage2_37[19],stage2_36[54],stage2_35[81]}
   );
   gpc615_5 gpc6596 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[37]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[12],stage2_37[20],stage2_36[55],stage2_35[82]}
   );
   gpc615_5 gpc6597 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[38]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[13],stage2_37[21],stage2_36[56],stage2_35[83]}
   );
   gpc615_5 gpc6598 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[39]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[14],stage2_37[22],stage2_36[57],stage2_35[84]}
   );
   gpc615_5 gpc6599 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[40]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[15],stage2_37[23],stage2_36[58],stage2_35[85]}
   );
   gpc615_5 gpc6600 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[41]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[16],stage2_37[24],stage2_36[59],stage2_35[86]}
   );
   gpc615_5 gpc6601 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[42]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[17],stage2_37[25],stage2_36[60],stage2_35[87]}
   );
   gpc615_5 gpc6602 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[43]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[18],stage2_37[26],stage2_36[61],stage2_35[88]}
   );
   gpc615_5 gpc6603 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[44]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[19],stage2_37[27],stage2_36[62],stage2_35[89]}
   );
   gpc615_5 gpc6604 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[45]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[20],stage2_37[28],stage2_36[63],stage2_35[90]}
   );
   gpc615_5 gpc6605 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[46]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[21],stage2_37[29],stage2_36[64],stage2_35[91]}
   );
   gpc615_5 gpc6606 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[47]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[22],stage2_37[30],stage2_36[65],stage2_35[92]}
   );
   gpc615_5 gpc6607 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[48]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[23],stage2_37[31],stage2_36[66],stage2_35[93]}
   );
   gpc615_5 gpc6608 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[49]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[24],stage2_37[32],stage2_36[67],stage2_35[94]}
   );
   gpc615_5 gpc6609 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[50]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[25],stage2_37[33],stage2_36[68],stage2_35[95]}
   );
   gpc615_5 gpc6610 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[51]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[26],stage2_37[34],stage2_36[69],stage2_35[96]}
   );
   gpc615_5 gpc6611 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[52]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[27],stage2_37[35],stage2_36[70],stage2_35[97]}
   );
   gpc615_5 gpc6612 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[53]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[28],stage2_37[36],stage2_36[71],stage2_35[98]}
   );
   gpc615_5 gpc6613 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[54]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[29],stage2_37[37],stage2_36[72],stage2_35[99]}
   );
   gpc1163_5 gpc6614 (
      {stage1_36[55], stage1_36[56], stage1_36[57]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage1_38[0]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[25],stage2_38[30],stage2_37[38],stage2_36[73]}
   );
   gpc606_5 gpc6615 (
      {stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61], stage1_36[62], stage1_36[63]},
      {stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6]},
      {stage2_40[1],stage2_39[26],stage2_38[31],stage2_37[39],stage2_36[74]}
   );
   gpc606_5 gpc6616 (
      {stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67], stage1_36[68], stage1_36[69]},
      {stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12]},
      {stage2_40[2],stage2_39[27],stage2_38[32],stage2_37[40],stage2_36[75]}
   );
   gpc606_5 gpc6617 (
      {stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73], stage1_36[74], stage1_36[75]},
      {stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18]},
      {stage2_40[3],stage2_39[28],stage2_38[33],stage2_37[41],stage2_36[76]}
   );
   gpc606_5 gpc6618 (
      {stage1_36[76], stage1_36[77], stage1_36[78], stage1_36[79], stage1_36[80], stage1_36[81]},
      {stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24]},
      {stage2_40[4],stage2_39[29],stage2_38[34],stage2_37[42],stage2_36[77]}
   );
   gpc606_5 gpc6619 (
      {stage1_36[82], stage1_36[83], stage1_36[84], stage1_36[85], stage1_36[86], stage1_36[87]},
      {stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30]},
      {stage2_40[5],stage2_39[30],stage2_38[35],stage2_37[43],stage2_36[78]}
   );
   gpc606_5 gpc6620 (
      {stage1_36[88], stage1_36[89], stage1_36[90], stage1_36[91], stage1_36[92], stage1_36[93]},
      {stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36]},
      {stage2_40[6],stage2_39[31],stage2_38[36],stage2_37[44],stage2_36[79]}
   );
   gpc606_5 gpc6621 (
      {stage1_36[94], stage1_36[95], stage1_36[96], stage1_36[97], stage1_36[98], stage1_36[99]},
      {stage1_38[37], stage1_38[38], stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42]},
      {stage2_40[7],stage2_39[32],stage2_38[37],stage2_37[45],stage2_36[80]}
   );
   gpc606_5 gpc6622 (
      {stage1_36[100], stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105]},
      {stage1_38[43], stage1_38[44], stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48]},
      {stage2_40[8],stage2_39[33],stage2_38[38],stage2_37[46],stage2_36[81]}
   );
   gpc606_5 gpc6623 (
      {stage1_36[106], stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111]},
      {stage1_38[49], stage1_38[50], stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54]},
      {stage2_40[9],stage2_39[34],stage2_38[39],stage2_37[47],stage2_36[82]}
   );
   gpc606_5 gpc6624 (
      {stage1_36[112], stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117]},
      {stage1_38[55], stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage2_40[10],stage2_39[35],stage2_38[40],stage2_37[48],stage2_36[83]}
   );
   gpc606_5 gpc6625 (
      {stage1_36[118], stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123]},
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65], stage1_38[66]},
      {stage2_40[11],stage2_39[36],stage2_38[41],stage2_37[49],stage2_36[84]}
   );
   gpc606_5 gpc6626 (
      {stage1_36[124], stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129]},
      {stage1_38[67], stage1_38[68], stage1_38[69], stage1_38[70], stage1_38[71], stage1_38[72]},
      {stage2_40[12],stage2_39[37],stage2_38[42],stage2_37[50],stage2_36[85]}
   );
   gpc606_5 gpc6627 (
      {stage1_36[130], stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135]},
      {stage1_38[73], stage1_38[74], stage1_38[75], stage1_38[76], stage1_38[77], stage1_38[78]},
      {stage2_40[13],stage2_39[38],stage2_38[43],stage2_37[51],stage2_36[86]}
   );
   gpc606_5 gpc6628 (
      {stage1_36[136], stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141]},
      {stage1_38[79], stage1_38[80], stage1_38[81], stage1_38[82], stage1_38[83], stage1_38[84]},
      {stage2_40[14],stage2_39[39],stage2_38[44],stage2_37[52],stage2_36[87]}
   );
   gpc606_5 gpc6629 (
      {stage1_36[142], stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147]},
      {stage1_38[85], stage1_38[86], stage1_38[87], stage1_38[88], stage1_38[89], stage1_38[90]},
      {stage2_40[15],stage2_39[40],stage2_38[45],stage2_37[53],stage2_36[88]}
   );
   gpc606_5 gpc6630 (
      {stage1_36[148], stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153]},
      {stage1_38[91], stage1_38[92], stage1_38[93], stage1_38[94], stage1_38[95], stage1_38[96]},
      {stage2_40[16],stage2_39[41],stage2_38[46],stage2_37[54],stage2_36[89]}
   );
   gpc606_5 gpc6631 (
      {stage1_36[154], stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159]},
      {stage1_38[97], stage1_38[98], stage1_38[99], stage1_38[100], stage1_38[101], stage1_38[102]},
      {stage2_40[17],stage2_39[42],stage2_38[47],stage2_37[55],stage2_36[90]}
   );
   gpc606_5 gpc6632 (
      {stage1_36[160], stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165]},
      {stage1_38[103], stage1_38[104], stage1_38[105], stage1_38[106], stage1_38[107], stage1_38[108]},
      {stage2_40[18],stage2_39[43],stage2_38[48],stage2_37[56],stage2_36[91]}
   );
   gpc606_5 gpc6633 (
      {stage1_36[166], stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171]},
      {stage1_38[109], stage1_38[110], stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114]},
      {stage2_40[19],stage2_39[44],stage2_38[49],stage2_37[57],stage2_36[92]}
   );
   gpc606_5 gpc6634 (
      {stage1_36[172], stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177]},
      {stage1_38[115], stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage2_40[20],stage2_39[45],stage2_38[50],stage2_37[58],stage2_36[93]}
   );
   gpc606_5 gpc6635 (
      {stage1_36[178], stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183]},
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125], stage1_38[126]},
      {stage2_40[21],stage2_39[46],stage2_38[51],stage2_37[59],stage2_36[94]}
   );
   gpc606_5 gpc6636 (
      {stage1_36[184], stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189]},
      {stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130], stage1_38[131], stage1_38[132]},
      {stage2_40[22],stage2_39[47],stage2_38[52],stage2_37[60],stage2_36[95]}
   );
   gpc606_5 gpc6637 (
      {stage1_36[190], stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195]},
      {stage1_38[133], stage1_38[134], stage1_38[135], stage1_38[136], stage1_38[137], stage1_38[138]},
      {stage2_40[23],stage2_39[48],stage2_38[53],stage2_37[61],stage2_36[96]}
   );
   gpc606_5 gpc6638 (
      {stage1_36[196], stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201]},
      {stage1_38[139], stage1_38[140], stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144]},
      {stage2_40[24],stage2_39[49],stage2_38[54],stage2_37[62],stage2_36[97]}
   );
   gpc606_5 gpc6639 (
      {stage1_36[202], stage1_36[203], stage1_36[204], stage1_36[205], stage1_36[206], stage1_36[207]},
      {stage1_38[145], stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage2_40[25],stage2_39[50],stage2_38[55],stage2_37[63],stage2_36[98]}
   );
   gpc606_5 gpc6640 (
      {stage1_36[208], stage1_36[209], stage1_36[210], stage1_36[211], stage1_36[212], stage1_36[213]},
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155], stage1_38[156]},
      {stage2_40[26],stage2_39[51],stage2_38[56],stage2_37[64],stage2_36[99]}
   );
   gpc606_5 gpc6641 (
      {stage1_36[214], stage1_36[215], stage1_36[216], stage1_36[217], stage1_36[218], stage1_36[219]},
      {stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160], stage1_38[161], stage1_38[162]},
      {stage2_40[27],stage2_39[52],stage2_38[57],stage2_37[65],stage2_36[100]}
   );
   gpc606_5 gpc6642 (
      {stage1_36[220], stage1_36[221], stage1_36[222], stage1_36[223], stage1_36[224], stage1_36[225]},
      {stage1_38[163], stage1_38[164], stage1_38[165], stage1_38[166], stage1_38[167], stage1_38[168]},
      {stage2_40[28],stage2_39[53],stage2_38[58],stage2_37[66],stage2_36[101]}
   );
   gpc606_5 gpc6643 (
      {stage1_36[226], stage1_36[227], stage1_36[228], stage1_36[229], stage1_36[230], stage1_36[231]},
      {stage1_38[169], stage1_38[170], stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174]},
      {stage2_40[29],stage2_39[54],stage2_38[59],stage2_37[67],stage2_36[102]}
   );
   gpc606_5 gpc6644 (
      {stage1_36[232], stage1_36[233], stage1_36[234], stage1_36[235], stage1_36[236], stage1_36[237]},
      {stage1_38[175], stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage2_40[30],stage2_39[55],stage2_38[60],stage2_37[68],stage2_36[103]}
   );
   gpc606_5 gpc6645 (
      {stage1_36[238], stage1_36[239], stage1_36[240], stage1_36[241], stage1_36[242], stage1_36[243]},
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185], stage1_38[186]},
      {stage2_40[31],stage2_39[56],stage2_38[61],stage2_37[69],stage2_36[104]}
   );
   gpc606_5 gpc6646 (
      {stage1_36[244], stage1_36[245], stage1_36[246], stage1_36[247], stage1_36[248], stage1_36[249]},
      {stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190], stage1_38[191], stage1_38[192]},
      {stage2_40[32],stage2_39[57],stage2_38[62],stage2_37[70],stage2_36[105]}
   );
   gpc606_5 gpc6647 (
      {stage1_36[250], stage1_36[251], stage1_36[252], stage1_36[253], stage1_36[254], stage1_36[255]},
      {stage1_38[193], stage1_38[194], stage1_38[195], stage1_38[196], stage1_38[197], stage1_38[198]},
      {stage2_40[33],stage2_39[58],stage2_38[63],stage2_37[71],stage2_36[106]}
   );
   gpc606_5 gpc6648 (
      {stage1_36[256], stage1_36[257], stage1_36[258], stage1_36[259], stage1_36[260], stage1_36[261]},
      {stage1_38[199], stage1_38[200], stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204]},
      {stage2_40[34],stage2_39[59],stage2_38[64],stage2_37[72],stage2_36[107]}
   );
   gpc606_5 gpc6649 (
      {stage1_36[262], stage1_36[263], stage1_36[264], stage1_36[265], stage1_36[266], stage1_36[267]},
      {stage1_38[205], stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage2_40[35],stage2_39[60],stage2_38[65],stage2_37[73],stage2_36[108]}
   );
   gpc606_5 gpc6650 (
      {stage1_36[268], stage1_36[269], stage1_36[270], stage1_36[271], stage1_36[272], stage1_36[273]},
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215], stage1_38[216]},
      {stage2_40[36],stage2_39[61],stage2_38[66],stage2_37[74],stage2_36[109]}
   );
   gpc606_5 gpc6651 (
      {stage1_36[274], stage1_36[275], stage1_36[276], stage1_36[277], stage1_36[278], stage1_36[279]},
      {stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220], stage1_38[221], stage1_38[222]},
      {stage2_40[37],stage2_39[62],stage2_38[67],stage2_37[75],stage2_36[110]}
   );
   gpc606_5 gpc6652 (
      {stage1_36[280], stage1_36[281], stage1_36[282], stage1_36[283], stage1_36[284], stage1_36[285]},
      {stage1_38[223], stage1_38[224], stage1_38[225], stage1_38[226], stage1_38[227], stage1_38[228]},
      {stage2_40[38],stage2_39[63],stage2_38[68],stage2_37[76],stage2_36[111]}
   );
   gpc606_5 gpc6653 (
      {stage1_36[286], stage1_36[287], stage1_36[288], stage1_36[289], stage1_36[290], stage1_36[291]},
      {stage1_38[229], stage1_38[230], stage1_38[231], stage1_38[232], stage1_38[233], stage1_38[234]},
      {stage2_40[39],stage2_39[64],stage2_38[69],stage2_37[77],stage2_36[112]}
   );
   gpc606_5 gpc6654 (
      {stage1_36[292], stage1_36[293], stage1_36[294], stage1_36[295], stage1_36[296], stage1_36[297]},
      {stage1_38[235], stage1_38[236], stage1_38[237], stage1_38[238], stage1_38[239], stage1_38[240]},
      {stage2_40[40],stage2_39[65],stage2_38[70],stage2_37[78],stage2_36[113]}
   );
   gpc606_5 gpc6655 (
      {stage1_36[298], stage1_36[299], stage1_36[300], stage1_36[301], stage1_36[302], stage1_36[303]},
      {stage1_38[241], stage1_38[242], stage1_38[243], stage1_38[244], stage1_38[245], stage1_38[246]},
      {stage2_40[41],stage2_39[66],stage2_38[71],stage2_37[79],stage2_36[114]}
   );
   gpc606_5 gpc6656 (
      {stage1_36[304], stage1_36[305], stage1_36[306], stage1_36[307], stage1_36[308], stage1_36[309]},
      {stage1_38[247], stage1_38[248], stage1_38[249], stage1_38[250], stage1_38[251], stage1_38[252]},
      {stage2_40[42],stage2_39[67],stage2_38[72],stage2_37[80],stage2_36[115]}
   );
   gpc606_5 gpc6657 (
      {stage1_36[310], stage1_36[311], stage1_36[312], stage1_36[313], stage1_36[314], stage1_36[315]},
      {stage1_38[253], stage1_38[254], stage1_38[255], stage1_38[256], stage1_38[257], stage1_38[258]},
      {stage2_40[43],stage2_39[68],stage2_38[73],stage2_37[81],stage2_36[116]}
   );
   gpc615_5 gpc6658 (
      {stage1_36[316], stage1_36[317], stage1_36[318], stage1_36[319], stage1_36[320]},
      {stage1_37[156]},
      {stage1_38[259], stage1_38[260], stage1_38[261], stage1_38[262], stage1_38[263], stage1_38[264]},
      {stage2_40[44],stage2_39[69],stage2_38[74],stage2_37[82],stage2_36[117]}
   );
   gpc615_5 gpc6659 (
      {stage1_36[321], stage1_36[322], stage1_36[323], stage1_36[324], stage1_36[325]},
      {stage1_37[157]},
      {stage1_38[265], stage1_38[266], stage1_38[267], stage1_38[268], stage1_38[269], stage1_38[270]},
      {stage2_40[45],stage2_39[70],stage2_38[75],stage2_37[83],stage2_36[118]}
   );
   gpc615_5 gpc6660 (
      {stage1_36[326], stage1_36[327], stage1_36[328], stage1_36[329], stage1_36[330]},
      {stage1_37[158]},
      {stage1_38[271], stage1_38[272], stage1_38[273], stage1_38[274], stage1_38[275], stage1_38[276]},
      {stage2_40[46],stage2_39[71],stage2_38[76],stage2_37[84],stage2_36[119]}
   );
   gpc606_5 gpc6661 (
      {stage1_37[159], stage1_37[160], stage1_37[161], stage1_37[162], stage1_37[163], stage1_37[164]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[47],stage2_39[72],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc6662 (
      {stage1_37[165], stage1_37[166], stage1_37[167], stage1_37[168], stage1_37[169], stage1_37[170]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[48],stage2_39[73],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc6663 (
      {stage1_37[171], stage1_37[172], stage1_37[173], stage1_37[174], stage1_37[175], stage1_37[176]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[49],stage2_39[74],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc6664 (
      {stage1_37[177], stage1_37[178], stage1_37[179], stage1_37[180], stage1_37[181], stage1_37[182]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[50],stage2_39[75],stage2_38[80],stage2_37[88]}
   );
   gpc606_5 gpc6665 (
      {stage1_37[183], stage1_37[184], stage1_37[185], stage1_37[186], stage1_37[187], stage1_37[188]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[51],stage2_39[76],stage2_38[81],stage2_37[89]}
   );
   gpc606_5 gpc6666 (
      {stage1_37[189], stage1_37[190], stage1_37[191], stage1_37[192], stage1_37[193], stage1_37[194]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[52],stage2_39[77],stage2_38[82],stage2_37[90]}
   );
   gpc606_5 gpc6667 (
      {stage1_37[195], stage1_37[196], stage1_37[197], stage1_37[198], stage1_37[199], stage1_37[200]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[53],stage2_39[78],stage2_38[83],stage2_37[91]}
   );
   gpc606_5 gpc6668 (
      {stage1_37[201], stage1_37[202], stage1_37[203], stage1_37[204], stage1_37[205], stage1_37[206]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[54],stage2_39[79],stage2_38[84],stage2_37[92]}
   );
   gpc606_5 gpc6669 (
      {stage1_37[207], stage1_37[208], stage1_37[209], stage1_37[210], stage1_37[211], stage1_37[212]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[55],stage2_39[80],stage2_38[85],stage2_37[93]}
   );
   gpc606_5 gpc6670 (
      {stage1_37[213], stage1_37[214], stage1_37[215], stage1_37[216], stage1_37[217], stage1_37[218]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[56],stage2_39[81],stage2_38[86],stage2_37[94]}
   );
   gpc606_5 gpc6671 (
      {stage1_37[219], stage1_37[220], stage1_37[221], stage1_37[222], stage1_37[223], stage1_37[224]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[57],stage2_39[82],stage2_38[87],stage2_37[95]}
   );
   gpc606_5 gpc6672 (
      {stage1_37[225], stage1_37[226], stage1_37[227], stage1_37[228], stage1_37[229], stage1_37[230]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[58],stage2_39[83],stage2_38[88],stage2_37[96]}
   );
   gpc606_5 gpc6673 (
      {stage1_37[231], stage1_37[232], stage1_37[233], stage1_37[234], stage1_37[235], stage1_37[236]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[59],stage2_39[84],stage2_38[89],stage2_37[97]}
   );
   gpc606_5 gpc6674 (
      {stage1_37[237], stage1_37[238], stage1_37[239], stage1_37[240], stage1_37[241], stage1_37[242]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[60],stage2_39[85],stage2_38[90],stage2_37[98]}
   );
   gpc606_5 gpc6675 (
      {stage1_37[243], stage1_37[244], stage1_37[245], stage1_37[246], stage1_37[247], stage1_37[248]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[61],stage2_39[86],stage2_38[91],stage2_37[99]}
   );
   gpc606_5 gpc6676 (
      {stage1_37[249], stage1_37[250], stage1_37[251], stage1_37[252], stage1_37[253], stage1_37[254]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[62],stage2_39[87],stage2_38[92],stage2_37[100]}
   );
   gpc606_5 gpc6677 (
      {stage1_37[255], stage1_37[256], stage1_37[257], stage1_37[258], stage1_37[259], stage1_37[260]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[63],stage2_39[88],stage2_38[93],stage2_37[101]}
   );
   gpc606_5 gpc6678 (
      {stage1_37[261], stage1_37[262], stage1_37[263], stage1_37[264], stage1_37[265], stage1_37[266]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[64],stage2_39[89],stage2_38[94],stage2_37[102]}
   );
   gpc606_5 gpc6679 (
      {stage1_37[267], stage1_37[268], stage1_37[269], stage1_37[270], stage1_37[271], stage1_37[272]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[65],stage2_39[90],stage2_38[95],stage2_37[103]}
   );
   gpc606_5 gpc6680 (
      {stage1_37[273], stage1_37[274], stage1_37[275], stage1_37[276], stage1_37[277], stage1_37[278]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[66],stage2_39[91],stage2_38[96],stage2_37[104]}
   );
   gpc606_5 gpc6681 (
      {stage1_37[279], stage1_37[280], stage1_37[281], stage1_37[282], stage1_37[283], stage1_37[284]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[67],stage2_39[92],stage2_38[97],stage2_37[105]}
   );
   gpc606_5 gpc6682 (
      {stage1_37[285], stage1_37[286], stage1_37[287], stage1_37[288], stage1_37[289], stage1_37[290]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[68],stage2_39[93],stage2_38[98],stage2_37[106]}
   );
   gpc606_5 gpc6683 (
      {stage1_37[291], stage1_37[292], stage1_37[293], stage1_37[294], stage1_37[295], stage1_37[296]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[69],stage2_39[94],stage2_38[99],stage2_37[107]}
   );
   gpc606_5 gpc6684 (
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[0],stage2_41[23],stage2_40[70],stage2_39[95]}
   );
   gpc606_5 gpc6685 (
      {stage1_39[145], stage1_39[146], stage1_39[147], stage1_39[148], stage1_39[149], stage1_39[150]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage2_43[1],stage2_42[1],stage2_41[24],stage2_40[71],stage2_39[96]}
   );
   gpc606_5 gpc6686 (
      {stage1_39[151], stage1_39[152], stage1_39[153], stage1_39[154], stage1_39[155], stage1_39[156]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage2_43[2],stage2_42[2],stage2_41[25],stage2_40[72],stage2_39[97]}
   );
   gpc606_5 gpc6687 (
      {stage1_39[157], stage1_39[158], stage1_39[159], stage1_39[160], stage1_39[161], stage1_39[162]},
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage2_43[3],stage2_42[3],stage2_41[26],stage2_40[73],stage2_39[98]}
   );
   gpc606_5 gpc6688 (
      {stage1_39[163], stage1_39[164], stage1_39[165], stage1_39[166], stage1_39[167], stage1_39[168]},
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage2_43[4],stage2_42[4],stage2_41[27],stage2_40[74],stage2_39[99]}
   );
   gpc615_5 gpc6689 (
      {stage1_39[169], stage1_39[170], stage1_39[171], stage1_39[172], stage1_39[173]},
      {stage1_40[0]},
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage2_43[5],stage2_42[5],stage2_41[28],stage2_40[75],stage2_39[100]}
   );
   gpc615_5 gpc6690 (
      {stage1_39[174], stage1_39[175], stage1_39[176], stage1_39[177], stage1_39[178]},
      {stage1_40[1]},
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage2_43[6],stage2_42[6],stage2_41[29],stage2_40[76],stage2_39[101]}
   );
   gpc615_5 gpc6691 (
      {stage1_39[179], stage1_39[180], stage1_39[181], stage1_39[182], stage1_39[183]},
      {stage1_40[2]},
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage2_43[7],stage2_42[7],stage2_41[30],stage2_40[77],stage2_39[102]}
   );
   gpc615_5 gpc6692 (
      {stage1_39[184], stage1_39[185], stage1_39[186], stage1_39[187], stage1_39[188]},
      {stage1_40[3]},
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52], stage1_41[53]},
      {stage2_43[8],stage2_42[8],stage2_41[31],stage2_40[78],stage2_39[103]}
   );
   gpc615_5 gpc6693 (
      {stage1_39[189], stage1_39[190], stage1_39[191], stage1_39[192], stage1_39[193]},
      {stage1_40[4]},
      {stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57], stage1_41[58], stage1_41[59]},
      {stage2_43[9],stage2_42[9],stage2_41[32],stage2_40[79],stage2_39[104]}
   );
   gpc606_5 gpc6694 (
      {stage1_40[5], stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[10],stage2_42[10],stage2_41[33],stage2_40[80]}
   );
   gpc606_5 gpc6695 (
      {stage1_40[11], stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[11],stage2_42[11],stage2_41[34],stage2_40[81]}
   );
   gpc606_5 gpc6696 (
      {stage1_40[17], stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[12],stage2_42[12],stage2_41[35],stage2_40[82]}
   );
   gpc606_5 gpc6697 (
      {stage1_40[23], stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[13],stage2_42[13],stage2_41[36],stage2_40[83]}
   );
   gpc606_5 gpc6698 (
      {stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[14],stage2_42[14],stage2_41[37],stage2_40[84]}
   );
   gpc606_5 gpc6699 (
      {stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[15],stage2_42[15],stage2_41[38],stage2_40[85]}
   );
   gpc606_5 gpc6700 (
      {stage1_40[41], stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[16],stage2_42[16],stage2_41[39],stage2_40[86]}
   );
   gpc606_5 gpc6701 (
      {stage1_40[47], stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[17],stage2_42[17],stage2_41[40],stage2_40[87]}
   );
   gpc606_5 gpc6702 (
      {stage1_40[53], stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[18],stage2_42[18],stage2_41[41],stage2_40[88]}
   );
   gpc606_5 gpc6703 (
      {stage1_40[59], stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[19],stage2_42[19],stage2_41[42],stage2_40[89]}
   );
   gpc606_5 gpc6704 (
      {stage1_40[65], stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[20],stage2_42[20],stage2_41[43],stage2_40[90]}
   );
   gpc606_5 gpc6705 (
      {stage1_40[71], stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[21],stage2_42[21],stage2_41[44],stage2_40[91]}
   );
   gpc606_5 gpc6706 (
      {stage1_40[77], stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[22],stage2_42[22],stage2_41[45],stage2_40[92]}
   );
   gpc606_5 gpc6707 (
      {stage1_40[83], stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[23],stage2_42[23],stage2_41[46],stage2_40[93]}
   );
   gpc606_5 gpc6708 (
      {stage1_40[89], stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[24],stage2_42[24],stage2_41[47],stage2_40[94]}
   );
   gpc606_5 gpc6709 (
      {stage1_40[95], stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[25],stage2_42[25],stage2_41[48],stage2_40[95]}
   );
   gpc606_5 gpc6710 (
      {stage1_40[101], stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[26],stage2_42[26],stage2_41[49],stage2_40[96]}
   );
   gpc606_5 gpc6711 (
      {stage1_40[107], stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[27],stage2_42[27],stage2_41[50],stage2_40[97]}
   );
   gpc606_5 gpc6712 (
      {stage1_40[113], stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[28],stage2_42[28],stage2_41[51],stage2_40[98]}
   );
   gpc606_5 gpc6713 (
      {stage1_40[119], stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[29],stage2_42[29],stage2_41[52],stage2_40[99]}
   );
   gpc606_5 gpc6714 (
      {stage1_40[125], stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[30],stage2_42[30],stage2_41[53],stage2_40[100]}
   );
   gpc606_5 gpc6715 (
      {stage1_40[131], stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[31],stage2_42[31],stage2_41[54],stage2_40[101]}
   );
   gpc606_5 gpc6716 (
      {stage1_40[137], stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[32],stage2_42[32],stage2_41[55],stage2_40[102]}
   );
   gpc606_5 gpc6717 (
      {stage1_40[143], stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148]},
      {stage1_42[138], stage1_42[139], stage1_42[140], stage1_42[141], stage1_42[142], stage1_42[143]},
      {stage2_44[23],stage2_43[33],stage2_42[33],stage2_41[56],stage2_40[103]}
   );
   gpc606_5 gpc6718 (
      {stage1_40[149], stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154]},
      {stage1_42[144], stage1_42[145], stage1_42[146], stage1_42[147], stage1_42[148], stage1_42[149]},
      {stage2_44[24],stage2_43[34],stage2_42[34],stage2_41[57],stage2_40[104]}
   );
   gpc606_5 gpc6719 (
      {stage1_40[155], stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160]},
      {stage1_42[150], stage1_42[151], stage1_42[152], stage1_42[153], stage1_42[154], stage1_42[155]},
      {stage2_44[25],stage2_43[35],stage2_42[35],stage2_41[58],stage2_40[105]}
   );
   gpc606_5 gpc6720 (
      {stage1_40[161], stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166]},
      {stage1_42[156], stage1_42[157], stage1_42[158], stage1_42[159], stage1_42[160], stage1_42[161]},
      {stage2_44[26],stage2_43[36],stage2_42[36],stage2_41[59],stage2_40[106]}
   );
   gpc606_5 gpc6721 (
      {stage1_40[167], stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172]},
      {stage1_42[162], stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage2_44[27],stage2_43[37],stage2_42[37],stage2_41[60],stage2_40[107]}
   );
   gpc606_5 gpc6722 (
      {stage1_40[173], stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178]},
      {stage1_42[168], stage1_42[169], stage1_42[170], stage1_42[171], stage1_42[172], stage1_42[173]},
      {stage2_44[28],stage2_43[38],stage2_42[38],stage2_41[61],stage2_40[108]}
   );
   gpc606_5 gpc6723 (
      {stage1_40[179], stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184]},
      {stage1_42[174], stage1_42[175], stage1_42[176], stage1_42[177], stage1_42[178], stage1_42[179]},
      {stage2_44[29],stage2_43[39],stage2_42[39],stage2_41[62],stage2_40[109]}
   );
   gpc606_5 gpc6724 (
      {stage1_40[185], stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190]},
      {stage1_42[180], stage1_42[181], stage1_42[182], stage1_42[183], stage1_42[184], stage1_42[185]},
      {stage2_44[30],stage2_43[40],stage2_42[40],stage2_41[63],stage2_40[110]}
   );
   gpc606_5 gpc6725 (
      {stage1_40[191], stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196]},
      {stage1_42[186], stage1_42[187], stage1_42[188], stage1_42[189], stage1_42[190], stage1_42[191]},
      {stage2_44[31],stage2_43[41],stage2_42[41],stage2_41[64],stage2_40[111]}
   );
   gpc606_5 gpc6726 (
      {stage1_40[197], stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202]},
      {stage1_42[192], stage1_42[193], stage1_42[194], stage1_42[195], stage1_42[196], stage1_42[197]},
      {stage2_44[32],stage2_43[42],stage2_42[42],stage2_41[65],stage2_40[112]}
   );
   gpc606_5 gpc6727 (
      {stage1_41[60], stage1_41[61], stage1_41[62], stage1_41[63], stage1_41[64], stage1_41[65]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[33],stage2_43[43],stage2_42[43],stage2_41[66]}
   );
   gpc606_5 gpc6728 (
      {stage1_41[66], stage1_41[67], stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[34],stage2_43[44],stage2_42[44],stage2_41[67]}
   );
   gpc606_5 gpc6729 (
      {stage1_41[72], stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[35],stage2_43[45],stage2_42[45],stage2_41[68]}
   );
   gpc606_5 gpc6730 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82], stage1_41[83]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[36],stage2_43[46],stage2_42[46],stage2_41[69]}
   );
   gpc606_5 gpc6731 (
      {stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87], stage1_41[88], stage1_41[89]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[37],stage2_43[47],stage2_42[47],stage2_41[70]}
   );
   gpc606_5 gpc6732 (
      {stage1_41[90], stage1_41[91], stage1_41[92], stage1_41[93], stage1_41[94], stage1_41[95]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[38],stage2_43[48],stage2_42[48],stage2_41[71]}
   );
   gpc606_5 gpc6733 (
      {stage1_41[96], stage1_41[97], stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[39],stage2_43[49],stage2_42[49],stage2_41[72]}
   );
   gpc606_5 gpc6734 (
      {stage1_41[102], stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[40],stage2_43[50],stage2_42[50],stage2_41[73]}
   );
   gpc606_5 gpc6735 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112], stage1_41[113]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[41],stage2_43[51],stage2_42[51],stage2_41[74]}
   );
   gpc606_5 gpc6736 (
      {stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117], stage1_41[118], stage1_41[119]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[42],stage2_43[52],stage2_42[52],stage2_41[75]}
   );
   gpc606_5 gpc6737 (
      {stage1_41[120], stage1_41[121], stage1_41[122], stage1_41[123], stage1_41[124], stage1_41[125]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[43],stage2_43[53],stage2_42[53],stage2_41[76]}
   );
   gpc606_5 gpc6738 (
      {stage1_41[126], stage1_41[127], stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[44],stage2_43[54],stage2_42[54],stage2_41[77]}
   );
   gpc606_5 gpc6739 (
      {stage1_41[132], stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[45],stage2_43[55],stage2_42[55],stage2_41[78]}
   );
   gpc606_5 gpc6740 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142], stage1_41[143]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[46],stage2_43[56],stage2_42[56],stage2_41[79]}
   );
   gpc606_5 gpc6741 (
      {stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147], stage1_41[148], stage1_41[149]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[47],stage2_43[57],stage2_42[57],stage2_41[80]}
   );
   gpc606_5 gpc6742 (
      {stage1_41[150], stage1_41[151], stage1_41[152], stage1_41[153], stage1_41[154], stage1_41[155]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[48],stage2_43[58],stage2_42[58],stage2_41[81]}
   );
   gpc606_5 gpc6743 (
      {stage1_41[156], stage1_41[157], stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[49],stage2_43[59],stage2_42[59],stage2_41[82]}
   );
   gpc606_5 gpc6744 (
      {stage1_41[162], stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[50],stage2_43[60],stage2_42[60],stage2_41[83]}
   );
   gpc606_5 gpc6745 (
      {stage1_41[168], stage1_41[169], stage1_41[170], stage1_41[171], stage1_41[172], stage1_41[173]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[51],stage2_43[61],stage2_42[61],stage2_41[84]}
   );
   gpc606_5 gpc6746 (
      {stage1_41[174], stage1_41[175], stage1_41[176], stage1_41[177], stage1_41[178], stage1_41[179]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[52],stage2_43[62],stage2_42[62],stage2_41[85]}
   );
   gpc606_5 gpc6747 (
      {stage1_41[180], stage1_41[181], stage1_41[182], stage1_41[183], stage1_41[184], stage1_41[185]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[53],stage2_43[63],stage2_42[63],stage2_41[86]}
   );
   gpc606_5 gpc6748 (
      {stage1_41[186], stage1_41[187], stage1_41[188], stage1_41[189], stage1_41[190], stage1_41[191]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[54],stage2_43[64],stage2_42[64],stage2_41[87]}
   );
   gpc606_5 gpc6749 (
      {stage1_41[192], stage1_41[193], stage1_41[194], stage1_41[195], stage1_41[196], stage1_41[197]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[55],stage2_43[65],stage2_42[65],stage2_41[88]}
   );
   gpc606_5 gpc6750 (
      {stage1_41[198], stage1_41[199], stage1_41[200], stage1_41[201], stage1_41[202], stage1_41[203]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[56],stage2_43[66],stage2_42[66],stage2_41[89]}
   );
   gpc606_5 gpc6751 (
      {stage1_41[204], stage1_41[205], stage1_41[206], stage1_41[207], stage1_41[208], stage1_41[209]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[57],stage2_43[67],stage2_42[67],stage2_41[90]}
   );
   gpc606_5 gpc6752 (
      {stage1_41[210], stage1_41[211], stage1_41[212], stage1_41[213], stage1_41[214], stage1_41[215]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[58],stage2_43[68],stage2_42[68],stage2_41[91]}
   );
   gpc606_5 gpc6753 (
      {stage1_41[216], stage1_41[217], stage1_41[218], stage1_41[219], stage1_41[220], stage1_41[221]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[59],stage2_43[69],stage2_42[69],stage2_41[92]}
   );
   gpc606_5 gpc6754 (
      {stage1_41[222], stage1_41[223], stage1_41[224], stage1_41[225], stage1_41[226], stage1_41[227]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[60],stage2_43[70],stage2_42[70],stage2_41[93]}
   );
   gpc606_5 gpc6755 (
      {stage1_41[228], stage1_41[229], stage1_41[230], stage1_41[231], stage1_41[232], stage1_41[233]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[61],stage2_43[71],stage2_42[71],stage2_41[94]}
   );
   gpc606_5 gpc6756 (
      {stage1_41[234], stage1_41[235], stage1_41[236], stage1_41[237], stage1_41[238], stage1_41[239]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[62],stage2_43[72],stage2_42[72],stage2_41[95]}
   );
   gpc606_5 gpc6757 (
      {stage1_41[240], stage1_41[241], stage1_41[242], stage1_41[243], stage1_41[244], stage1_41[245]},
      {stage1_43[180], stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage2_45[30],stage2_44[63],stage2_43[73],stage2_42[73],stage2_41[96]}
   );
   gpc606_5 gpc6758 (
      {stage1_41[246], stage1_41[247], stage1_41[248], stage1_41[249], stage1_41[250], stage1_41[251]},
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190], stage1_43[191]},
      {stage2_45[31],stage2_44[64],stage2_43[74],stage2_42[74],stage2_41[97]}
   );
   gpc615_5 gpc6759 (
      {stage1_42[198], stage1_42[199], stage1_42[200], stage1_42[201], stage1_42[202]},
      {stage1_43[192]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[32],stage2_44[65],stage2_43[75],stage2_42[75]}
   );
   gpc615_5 gpc6760 (
      {stage1_42[203], stage1_42[204], stage1_42[205], stage1_42[206], stage1_42[207]},
      {stage1_43[193]},
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage2_46[1],stage2_45[33],stage2_44[66],stage2_43[76],stage2_42[76]}
   );
   gpc615_5 gpc6761 (
      {stage1_42[208], stage1_42[209], stage1_42[210], stage1_42[211], stage1_42[212]},
      {stage1_43[194]},
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage2_46[2],stage2_45[34],stage2_44[67],stage2_43[77],stage2_42[77]}
   );
   gpc615_5 gpc6762 (
      {stage1_42[213], stage1_42[214], stage1_42[215], stage1_42[216], stage1_42[217]},
      {stage1_43[195]},
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage2_46[3],stage2_45[35],stage2_44[68],stage2_43[78],stage2_42[78]}
   );
   gpc615_5 gpc6763 (
      {stage1_42[218], stage1_42[219], stage1_42[220], stage1_42[221], stage1_42[222]},
      {stage1_43[196]},
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage2_46[4],stage2_45[36],stage2_44[69],stage2_43[79],stage2_42[79]}
   );
   gpc615_5 gpc6764 (
      {stage1_42[223], stage1_42[224], stage1_42[225], stage1_42[226], stage1_42[227]},
      {stage1_43[197]},
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage2_46[5],stage2_45[37],stage2_44[70],stage2_43[80],stage2_42[80]}
   );
   gpc1415_5 gpc6765 (
      {stage1_43[198], stage1_43[199], stage1_43[200], stage1_43[201], stage1_43[202]},
      {stage1_44[36]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3]},
      {stage1_46[0]},
      {stage2_47[0],stage2_46[6],stage2_45[38],stage2_44[71],stage2_43[81]}
   );
   gpc1415_5 gpc6766 (
      {stage1_43[203], stage1_43[204], stage1_43[205], stage1_43[206], stage1_43[207]},
      {stage1_44[37]},
      {stage1_45[4], stage1_45[5], stage1_45[6], stage1_45[7]},
      {stage1_46[1]},
      {stage2_47[1],stage2_46[7],stage2_45[39],stage2_44[72],stage2_43[82]}
   );
   gpc1415_5 gpc6767 (
      {stage1_43[208], stage1_43[209], stage1_43[210], stage1_43[211], stage1_43[212]},
      {stage1_44[38]},
      {stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage1_46[2]},
      {stage2_47[2],stage2_46[8],stage2_45[40],stage2_44[73],stage2_43[83]}
   );
   gpc1415_5 gpc6768 (
      {stage1_43[213], stage1_43[214], stage1_43[215], stage1_43[216], stage1_43[217]},
      {stage1_44[39]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15]},
      {stage1_46[3]},
      {stage2_47[3],stage2_46[9],stage2_45[41],stage2_44[74],stage2_43[84]}
   );
   gpc606_5 gpc6769 (
      {stage1_44[40], stage1_44[41], stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45]},
      {stage1_46[4], stage1_46[5], stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9]},
      {stage2_48[0],stage2_47[4],stage2_46[10],stage2_45[42],stage2_44[75]}
   );
   gpc606_5 gpc6770 (
      {stage1_44[46], stage1_44[47], stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51]},
      {stage1_46[10], stage1_46[11], stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15]},
      {stage2_48[1],stage2_47[5],stage2_46[11],stage2_45[43],stage2_44[76]}
   );
   gpc606_5 gpc6771 (
      {stage1_44[52], stage1_44[53], stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57]},
      {stage1_46[16], stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage2_48[2],stage2_47[6],stage2_46[12],stage2_45[44],stage2_44[77]}
   );
   gpc606_5 gpc6772 (
      {stage1_44[58], stage1_44[59], stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63]},
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27]},
      {stage2_48[3],stage2_47[7],stage2_46[13],stage2_45[45],stage2_44[78]}
   );
   gpc606_5 gpc6773 (
      {stage1_44[64], stage1_44[65], stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69]},
      {stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33]},
      {stage2_48[4],stage2_47[8],stage2_46[14],stage2_45[46],stage2_44[79]}
   );
   gpc606_5 gpc6774 (
      {stage1_44[70], stage1_44[71], stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75]},
      {stage1_46[34], stage1_46[35], stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39]},
      {stage2_48[5],stage2_47[9],stage2_46[15],stage2_45[47],stage2_44[80]}
   );
   gpc606_5 gpc6775 (
      {stage1_44[76], stage1_44[77], stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81]},
      {stage1_46[40], stage1_46[41], stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45]},
      {stage2_48[6],stage2_47[10],stage2_46[16],stage2_45[48],stage2_44[81]}
   );
   gpc606_5 gpc6776 (
      {stage1_44[82], stage1_44[83], stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87]},
      {stage1_46[46], stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage2_48[7],stage2_47[11],stage2_46[17],stage2_45[49],stage2_44[82]}
   );
   gpc606_5 gpc6777 (
      {stage1_44[88], stage1_44[89], stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93]},
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57]},
      {stage2_48[8],stage2_47[12],stage2_46[18],stage2_45[50],stage2_44[83]}
   );
   gpc606_5 gpc6778 (
      {stage1_44[94], stage1_44[95], stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99]},
      {stage1_46[58], stage1_46[59], stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63]},
      {stage2_48[9],stage2_47[13],stage2_46[19],stage2_45[51],stage2_44[84]}
   );
   gpc606_5 gpc6779 (
      {stage1_44[100], stage1_44[101], stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105]},
      {stage1_46[64], stage1_46[65], stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69]},
      {stage2_48[10],stage2_47[14],stage2_46[20],stage2_45[52],stage2_44[85]}
   );
   gpc606_5 gpc6780 (
      {stage1_44[106], stage1_44[107], stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111]},
      {stage1_46[70], stage1_46[71], stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75]},
      {stage2_48[11],stage2_47[15],stage2_46[21],stage2_45[53],stage2_44[86]}
   );
   gpc606_5 gpc6781 (
      {stage1_44[112], stage1_44[113], stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117]},
      {stage1_46[76], stage1_46[77], stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81]},
      {stage2_48[12],stage2_47[16],stage2_46[22],stage2_45[54],stage2_44[87]}
   );
   gpc606_5 gpc6782 (
      {stage1_44[118], stage1_44[119], stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123]},
      {stage1_46[82], stage1_46[83], stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87]},
      {stage2_48[13],stage2_47[17],stage2_46[23],stage2_45[55],stage2_44[88]}
   );
   gpc615_5 gpc6783 (
      {stage1_44[124], stage1_44[125], stage1_44[126], stage1_44[127], stage1_44[128]},
      {stage1_45[16]},
      {stage1_46[88], stage1_46[89], stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93]},
      {stage2_48[14],stage2_47[18],stage2_46[24],stage2_45[56],stage2_44[89]}
   );
   gpc615_5 gpc6784 (
      {stage1_44[129], stage1_44[130], stage1_44[131], stage1_44[132], stage1_44[133]},
      {stage1_45[17]},
      {stage1_46[94], stage1_46[95], stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99]},
      {stage2_48[15],stage2_47[19],stage2_46[25],stage2_45[57],stage2_44[90]}
   );
   gpc615_5 gpc6785 (
      {stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137], stage1_44[138]},
      {stage1_45[18]},
      {stage1_46[100], stage1_46[101], stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105]},
      {stage2_48[16],stage2_47[20],stage2_46[26],stage2_45[58],stage2_44[91]}
   );
   gpc615_5 gpc6786 (
      {stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_45[19]},
      {stage1_46[106], stage1_46[107], stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111]},
      {stage2_48[17],stage2_47[21],stage2_46[27],stage2_45[59],stage2_44[92]}
   );
   gpc615_5 gpc6787 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148]},
      {stage1_45[20]},
      {stage1_46[112], stage1_46[113], stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117]},
      {stage2_48[18],stage2_47[22],stage2_46[28],stage2_45[60],stage2_44[93]}
   );
   gpc615_5 gpc6788 (
      {stage1_44[149], stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153]},
      {stage1_45[21]},
      {stage1_46[118], stage1_46[119], stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123]},
      {stage2_48[19],stage2_47[23],stage2_46[29],stage2_45[61],stage2_44[94]}
   );
   gpc615_5 gpc6789 (
      {stage1_44[154], stage1_44[155], stage1_44[156], stage1_44[157], stage1_44[158]},
      {stage1_45[22]},
      {stage1_46[124], stage1_46[125], stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129]},
      {stage2_48[20],stage2_47[24],stage2_46[30],stage2_45[62],stage2_44[95]}
   );
   gpc615_5 gpc6790 (
      {stage1_44[159], stage1_44[160], stage1_44[161], stage1_44[162], stage1_44[163]},
      {stage1_45[23]},
      {stage1_46[130], stage1_46[131], stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135]},
      {stage2_48[21],stage2_47[25],stage2_46[31],stage2_45[63],stage2_44[96]}
   );
   gpc615_5 gpc6791 (
      {stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167], stage1_44[168]},
      {stage1_45[24]},
      {stage1_46[136], stage1_46[137], stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141]},
      {stage2_48[22],stage2_47[26],stage2_46[32],stage2_45[64],stage2_44[97]}
   );
   gpc615_5 gpc6792 (
      {stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_45[25]},
      {stage1_46[142], stage1_46[143], stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147]},
      {stage2_48[23],stage2_47[27],stage2_46[33],stage2_45[65],stage2_44[98]}
   );
   gpc615_5 gpc6793 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178]},
      {stage1_45[26]},
      {stage1_46[148], stage1_46[149], stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153]},
      {stage2_48[24],stage2_47[28],stage2_46[34],stage2_45[66],stage2_44[99]}
   );
   gpc615_5 gpc6794 (
      {stage1_44[179], stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183]},
      {stage1_45[27]},
      {stage1_46[154], stage1_46[155], stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159]},
      {stage2_48[25],stage2_47[29],stage2_46[35],stage2_45[67],stage2_44[100]}
   );
   gpc615_5 gpc6795 (
      {stage1_44[184], stage1_44[185], stage1_44[186], stage1_44[187], stage1_44[188]},
      {stage1_45[28]},
      {stage1_46[160], stage1_46[161], stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165]},
      {stage2_48[26],stage2_47[30],stage2_46[36],stage2_45[68],stage2_44[101]}
   );
   gpc615_5 gpc6796 (
      {stage1_44[189], stage1_44[190], stage1_44[191], stage1_44[192], stage1_44[193]},
      {stage1_45[29]},
      {stage1_46[166], stage1_46[167], stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171]},
      {stage2_48[27],stage2_47[31],stage2_46[37],stage2_45[69],stage2_44[102]}
   );
   gpc615_5 gpc6797 (
      {stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197], stage1_44[198]},
      {stage1_45[30]},
      {stage1_46[172], stage1_46[173], stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177]},
      {stage2_48[28],stage2_47[32],stage2_46[38],stage2_45[70],stage2_44[103]}
   );
   gpc615_5 gpc6798 (
      {stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_45[31]},
      {stage1_46[178], stage1_46[179], stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183]},
      {stage2_48[29],stage2_47[33],stage2_46[39],stage2_45[71],stage2_44[104]}
   );
   gpc615_5 gpc6799 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208]},
      {stage1_45[32]},
      {stage1_46[184], stage1_46[185], stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189]},
      {stage2_48[30],stage2_47[34],stage2_46[40],stage2_45[72],stage2_44[105]}
   );
   gpc615_5 gpc6800 (
      {stage1_44[209], stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213]},
      {stage1_45[33]},
      {stage1_46[190], stage1_46[191], stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195]},
      {stage2_48[31],stage2_47[35],stage2_46[41],stage2_45[73],stage2_44[106]}
   );
   gpc615_5 gpc6801 (
      {stage1_44[214], stage1_44[215], stage1_44[216], stage1_44[217], stage1_44[218]},
      {stage1_45[34]},
      {stage1_46[196], stage1_46[197], stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201]},
      {stage2_48[32],stage2_47[36],stage2_46[42],stage2_45[74],stage2_44[107]}
   );
   gpc615_5 gpc6802 (
      {stage1_44[219], stage1_44[220], stage1_44[221], stage1_44[222], stage1_44[223]},
      {stage1_45[35]},
      {stage1_46[202], stage1_46[203], stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207]},
      {stage2_48[33],stage2_47[37],stage2_46[43],stage2_45[75],stage2_44[108]}
   );
   gpc615_5 gpc6803 (
      {stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227], stage1_44[228]},
      {stage1_45[36]},
      {stage1_46[208], stage1_46[209], stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213]},
      {stage2_48[34],stage2_47[38],stage2_46[44],stage2_45[76],stage2_44[109]}
   );
   gpc615_5 gpc6804 (
      {stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_45[37]},
      {stage1_46[214], stage1_46[215], stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219]},
      {stage2_48[35],stage2_47[39],stage2_46[45],stage2_45[77],stage2_44[110]}
   );
   gpc615_5 gpc6805 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238]},
      {stage1_45[38]},
      {stage1_46[220], stage1_46[221], stage1_46[222], stage1_46[223], stage1_46[224], stage1_46[225]},
      {stage2_48[36],stage2_47[40],stage2_46[46],stage2_45[78],stage2_44[111]}
   );
   gpc615_5 gpc6806 (
      {stage1_44[239], stage1_44[240], stage1_44[241], stage1_44[242], stage1_44[243]},
      {stage1_45[39]},
      {stage1_46[226], stage1_46[227], stage1_46[228], stage1_46[229], stage1_46[230], stage1_46[231]},
      {stage2_48[37],stage2_47[41],stage2_46[47],stage2_45[79],stage2_44[112]}
   );
   gpc606_5 gpc6807 (
      {stage1_45[40], stage1_45[41], stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[38],stage2_47[42],stage2_46[48],stage2_45[80]}
   );
   gpc606_5 gpc6808 (
      {stage1_45[46], stage1_45[47], stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[39],stage2_47[43],stage2_46[49],stage2_45[81]}
   );
   gpc606_5 gpc6809 (
      {stage1_45[52], stage1_45[53], stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[40],stage2_47[44],stage2_46[50],stage2_45[82]}
   );
   gpc606_5 gpc6810 (
      {stage1_45[58], stage1_45[59], stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[41],stage2_47[45],stage2_46[51],stage2_45[83]}
   );
   gpc606_5 gpc6811 (
      {stage1_45[64], stage1_45[65], stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[42],stage2_47[46],stage2_46[52],stage2_45[84]}
   );
   gpc606_5 gpc6812 (
      {stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[43],stage2_47[47],stage2_46[53],stage2_45[85]}
   );
   gpc606_5 gpc6813 (
      {stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[44],stage2_47[48],stage2_46[54],stage2_45[86]}
   );
   gpc606_5 gpc6814 (
      {stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[45],stage2_47[49],stage2_46[55],stage2_45[87]}
   );
   gpc606_5 gpc6815 (
      {stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[46],stage2_47[50],stage2_46[56],stage2_45[88]}
   );
   gpc606_5 gpc6816 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98], stage1_45[99]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[47],stage2_47[51],stage2_46[57],stage2_45[89]}
   );
   gpc606_5 gpc6817 (
      {stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103], stage1_45[104], stage1_45[105]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[48],stage2_47[52],stage2_46[58],stage2_45[90]}
   );
   gpc606_5 gpc6818 (
      {stage1_45[106], stage1_45[107], stage1_45[108], stage1_45[109], stage1_45[110], stage1_45[111]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[49],stage2_47[53],stage2_46[59],stage2_45[91]}
   );
   gpc606_5 gpc6819 (
      {stage1_45[112], stage1_45[113], stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[50],stage2_47[54],stage2_46[60],stage2_45[92]}
   );
   gpc606_5 gpc6820 (
      {stage1_45[118], stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[51],stage2_47[55],stage2_46[61],stage2_45[93]}
   );
   gpc606_5 gpc6821 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128], stage1_45[129]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[52],stage2_47[56],stage2_46[62],stage2_45[94]}
   );
   gpc606_5 gpc6822 (
      {stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133], stage1_45[134], stage1_45[135]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[53],stage2_47[57],stage2_46[63],stage2_45[95]}
   );
   gpc606_5 gpc6823 (
      {stage1_45[136], stage1_45[137], stage1_45[138], stage1_45[139], stage1_45[140], stage1_45[141]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[54],stage2_47[58],stage2_46[64],stage2_45[96]}
   );
   gpc615_5 gpc6824 (
      {stage1_45[142], stage1_45[143], stage1_45[144], stage1_45[145], stage1_45[146]},
      {stage1_46[232]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[55],stage2_47[59],stage2_46[65],stage2_45[97]}
   );
   gpc615_5 gpc6825 (
      {stage1_45[147], stage1_45[148], stage1_45[149], stage1_45[150], stage1_45[151]},
      {stage1_46[233]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[56],stage2_47[60],stage2_46[66],stage2_45[98]}
   );
   gpc615_5 gpc6826 (
      {stage1_45[152], stage1_45[153], stage1_45[154], stage1_45[155], stage1_45[156]},
      {stage1_46[234]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[57],stage2_47[61],stage2_46[67],stage2_45[99]}
   );
   gpc615_5 gpc6827 (
      {stage1_46[235], stage1_46[236], stage1_46[237], stage1_46[238], stage1_46[239]},
      {stage1_47[120]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[20],stage2_48[58],stage2_47[62],stage2_46[68]}
   );
   gpc615_5 gpc6828 (
      {stage1_46[240], stage1_46[241], stage1_46[242], stage1_46[243], stage1_46[244]},
      {stage1_47[121]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[21],stage2_48[59],stage2_47[63],stage2_46[69]}
   );
   gpc615_5 gpc6829 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[122]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[22],stage2_48[60],stage2_47[64],stage2_46[70]}
   );
   gpc615_5 gpc6830 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[123]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[23],stage2_48[61],stage2_47[65],stage2_46[71]}
   );
   gpc615_5 gpc6831 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[124]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[24],stage2_48[62],stage2_47[66],stage2_46[72]}
   );
   gpc615_5 gpc6832 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[125]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[25],stage2_48[63],stage2_47[67],stage2_46[73]}
   );
   gpc615_5 gpc6833 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[126]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[26],stage2_48[64],stage2_47[68],stage2_46[74]}
   );
   gpc615_5 gpc6834 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[127]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[27],stage2_48[65],stage2_47[69],stage2_46[75]}
   );
   gpc615_5 gpc6835 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[128]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[28],stage2_48[66],stage2_47[70],stage2_46[76]}
   );
   gpc615_5 gpc6836 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[129]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[29],stage2_48[67],stage2_47[71],stage2_46[77]}
   );
   gpc615_5 gpc6837 (
      {stage1_47[130], stage1_47[131], stage1_47[132], stage1_47[133], stage1_47[134]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[30],stage2_48[68],stage2_47[72]}
   );
   gpc615_5 gpc6838 (
      {stage1_47[135], stage1_47[136], stage1_47[137], stage1_47[138], stage1_47[139]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[31],stage2_48[69],stage2_47[73]}
   );
   gpc615_5 gpc6839 (
      {stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143], stage1_47[144]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[32],stage2_48[70],stage2_47[74]}
   );
   gpc615_5 gpc6840 (
      {stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[33],stage2_48[71],stage2_47[75]}
   );
   gpc615_5 gpc6841 (
      {stage1_47[150], stage1_47[151], stage1_47[152], stage1_47[153], stage1_47[154]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[34],stage2_48[72],stage2_47[76]}
   );
   gpc615_5 gpc6842 (
      {stage1_47[155], stage1_47[156], stage1_47[157], stage1_47[158], stage1_47[159]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[35],stage2_48[73],stage2_47[77]}
   );
   gpc615_5 gpc6843 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[36],stage2_48[74],stage2_47[78]}
   );
   gpc615_5 gpc6844 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[37],stage2_48[75],stage2_47[79]}
   );
   gpc615_5 gpc6845 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[38],stage2_48[76],stage2_47[80]}
   );
   gpc615_5 gpc6846 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[39],stage2_48[77],stage2_47[81]}
   );
   gpc615_5 gpc6847 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[40],stage2_48[78],stage2_47[82]}
   );
   gpc615_5 gpc6848 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[41],stage2_48[79],stage2_47[83]}
   );
   gpc615_5 gpc6849 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[42],stage2_48[80],stage2_47[84]}
   );
   gpc615_5 gpc6850 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[43],stage2_48[81],stage2_47[85]}
   );
   gpc615_5 gpc6851 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[74]},
      {stage1_49[84], stage1_49[85], stage1_49[86], stage1_49[87], stage1_49[88], stage1_49[89]},
      {stage2_51[14],stage2_50[24],stage2_49[44],stage2_48[82],stage2_47[86]}
   );
   gpc615_5 gpc6852 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[75]},
      {stage1_49[90], stage1_49[91], stage1_49[92], stage1_49[93], stage1_49[94], stage1_49[95]},
      {stage2_51[15],stage2_50[25],stage2_49[45],stage2_48[83],stage2_47[87]}
   );
   gpc615_5 gpc6853 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[76]},
      {stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99], stage1_49[100], stage1_49[101]},
      {stage2_51[16],stage2_50[26],stage2_49[46],stage2_48[84],stage2_47[88]}
   );
   gpc615_5 gpc6854 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[77]},
      {stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105], stage1_49[106], stage1_49[107]},
      {stage2_51[17],stage2_50[27],stage2_49[47],stage2_48[85],stage2_47[89]}
   );
   gpc615_5 gpc6855 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[78]},
      {stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111], stage1_49[112], stage1_49[113]},
      {stage2_51[18],stage2_50[28],stage2_49[48],stage2_48[86],stage2_47[90]}
   );
   gpc615_5 gpc6856 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[79]},
      {stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117], stage1_49[118], stage1_49[119]},
      {stage2_51[19],stage2_50[29],stage2_49[49],stage2_48[87],stage2_47[91]}
   );
   gpc615_5 gpc6857 (
      {stage1_47[230], stage1_47[231], stage1_47[232], stage1_47[233], stage1_47[234]},
      {stage1_48[80]},
      {stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123], stage1_49[124], stage1_49[125]},
      {stage2_51[20],stage2_50[30],stage2_49[50],stage2_48[88],stage2_47[92]}
   );
   gpc615_5 gpc6858 (
      {stage1_47[235], stage1_47[236], stage1_47[237], stage1_47[238], stage1_47[239]},
      {stage1_48[81]},
      {stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129], stage1_49[130], stage1_49[131]},
      {stage2_51[21],stage2_50[31],stage2_49[51],stage2_48[89],stage2_47[93]}
   );
   gpc615_5 gpc6859 (
      {stage1_47[240], stage1_47[241], stage1_47[242], stage1_47[243], stage1_47[244]},
      {stage1_48[82]},
      {stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135], stage1_49[136], stage1_49[137]},
      {stage2_51[22],stage2_50[32],stage2_49[52],stage2_48[90],stage2_47[94]}
   );
   gpc615_5 gpc6860 (
      {stage1_47[245], stage1_47[246], stage1_47[247], stage1_47[248], stage1_47[249]},
      {stage1_48[83]},
      {stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141], stage1_49[142], stage1_49[143]},
      {stage2_51[23],stage2_50[33],stage2_49[53],stage2_48[91],stage2_47[95]}
   );
   gpc615_5 gpc6861 (
      {stage1_47[250], stage1_47[251], stage1_47[252], stage1_47[253], stage1_47[254]},
      {stage1_48[84]},
      {stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147], stage1_49[148], stage1_49[149]},
      {stage2_51[24],stage2_50[34],stage2_49[54],stage2_48[92],stage2_47[96]}
   );
   gpc615_5 gpc6862 (
      {stage1_47[255], stage1_47[256], stage1_47[257], stage1_47[258], stage1_47[259]},
      {stage1_48[85]},
      {stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153], stage1_49[154], stage1_49[155]},
      {stage2_51[25],stage2_50[35],stage2_49[55],stage2_48[93],stage2_47[97]}
   );
   gpc615_5 gpc6863 (
      {stage1_47[260], stage1_47[261], stage1_47[262], stage1_47[263], stage1_47[264]},
      {stage1_48[86]},
      {stage1_49[156], stage1_49[157], stage1_49[158], stage1_49[159], stage1_49[160], stage1_49[161]},
      {stage2_51[26],stage2_50[36],stage2_49[56],stage2_48[94],stage2_47[98]}
   );
   gpc615_5 gpc6864 (
      {stage1_47[265], stage1_47[266], stage1_47[267], stage1_47[268], stage1_47[269]},
      {stage1_48[87]},
      {stage1_49[162], stage1_49[163], stage1_49[164], stage1_49[165], stage1_49[166], stage1_49[167]},
      {stage2_51[27],stage2_50[37],stage2_49[57],stage2_48[95],stage2_47[99]}
   );
   gpc606_5 gpc6865 (
      {stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91], stage1_48[92], stage1_48[93]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[28],stage2_50[38],stage2_49[58],stage2_48[96]}
   );
   gpc606_5 gpc6866 (
      {stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97], stage1_48[98], stage1_48[99]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[29],stage2_50[39],stage2_49[59],stage2_48[97]}
   );
   gpc606_5 gpc6867 (
      {stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103], stage1_48[104], stage1_48[105]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[30],stage2_50[40],stage2_49[60],stage2_48[98]}
   );
   gpc606_5 gpc6868 (
      {stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109], stage1_48[110], stage1_48[111]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[31],stage2_50[41],stage2_49[61],stage2_48[99]}
   );
   gpc606_5 gpc6869 (
      {stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115], stage1_48[116], stage1_48[117]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[32],stage2_50[42],stage2_49[62],stage2_48[100]}
   );
   gpc606_5 gpc6870 (
      {stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121], stage1_48[122], stage1_48[123]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[33],stage2_50[43],stage2_49[63],stage2_48[101]}
   );
   gpc606_5 gpc6871 (
      {stage1_48[124], stage1_48[125], stage1_48[126], stage1_48[127], stage1_48[128], stage1_48[129]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[34],stage2_50[44],stage2_49[64],stage2_48[102]}
   );
   gpc606_5 gpc6872 (
      {stage1_48[130], stage1_48[131], stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[35],stage2_50[45],stage2_49[65],stage2_48[103]}
   );
   gpc606_5 gpc6873 (
      {stage1_48[136], stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[36],stage2_50[46],stage2_49[66],stage2_48[104]}
   );
   gpc606_5 gpc6874 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146], stage1_48[147]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[37],stage2_50[47],stage2_49[67],stage2_48[105]}
   );
   gpc606_5 gpc6875 (
      {stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151], stage1_48[152], stage1_48[153]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[38],stage2_50[48],stage2_49[68],stage2_48[106]}
   );
   gpc606_5 gpc6876 (
      {stage1_48[154], stage1_48[155], stage1_48[156], stage1_48[157], stage1_48[158], stage1_48[159]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[39],stage2_50[49],stage2_49[69],stage2_48[107]}
   );
   gpc606_5 gpc6877 (
      {stage1_48[160], stage1_48[161], stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[40],stage2_50[50],stage2_49[70],stage2_48[108]}
   );
   gpc606_5 gpc6878 (
      {stage1_49[168], stage1_49[169], stage1_49[170], stage1_49[171], stage1_49[172], stage1_49[173]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[13],stage2_51[41],stage2_50[51],stage2_49[71]}
   );
   gpc606_5 gpc6879 (
      {stage1_49[174], stage1_49[175], stage1_49[176], stage1_49[177], stage1_49[178], stage1_49[179]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[14],stage2_51[42],stage2_50[52],stage2_49[72]}
   );
   gpc606_5 gpc6880 (
      {stage1_49[180], stage1_49[181], stage1_49[182], stage1_49[183], stage1_49[184], stage1_49[185]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[15],stage2_51[43],stage2_50[53],stage2_49[73]}
   );
   gpc606_5 gpc6881 (
      {stage1_49[186], stage1_49[187], stage1_49[188], stage1_49[189], stage1_49[190], stage1_49[191]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[16],stage2_51[44],stage2_50[54],stage2_49[74]}
   );
   gpc606_5 gpc6882 (
      {stage1_49[192], stage1_49[193], stage1_49[194], stage1_49[195], stage1_49[196], stage1_49[197]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[17],stage2_51[45],stage2_50[55],stage2_49[75]}
   );
   gpc615_5 gpc6883 (
      {stage1_49[198], stage1_49[199], stage1_49[200], stage1_49[201], stage1_49[202]},
      {stage1_50[78]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[18],stage2_51[46],stage2_50[56],stage2_49[76]}
   );
   gpc1163_5 gpc6884 (
      {stage1_50[79], stage1_50[80], stage1_50[81]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage1_52[0]},
      {stage1_53[0]},
      {stage2_54[0],stage2_53[6],stage2_52[19],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc6885 (
      {stage1_50[82], stage1_50[83], stage1_50[84]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage1_52[1]},
      {stage1_53[1]},
      {stage2_54[1],stage2_53[7],stage2_52[20],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc6886 (
      {stage1_50[85], stage1_50[86], stage1_50[87]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage1_52[2]},
      {stage1_53[2]},
      {stage2_54[2],stage2_53[8],stage2_52[21],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc6887 (
      {stage1_50[88], stage1_50[89], stage1_50[90]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage1_52[3]},
      {stage1_53[3]},
      {stage2_54[3],stage2_53[9],stage2_52[22],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc6888 (
      {stage1_50[91], stage1_50[92], stage1_50[93]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage1_52[4]},
      {stage1_53[4]},
      {stage2_54[4],stage2_53[10],stage2_52[23],stage2_51[51],stage2_50[61]}
   );
   gpc615_5 gpc6889 (
      {stage1_50[94], stage1_50[95], stage1_50[96], stage1_50[97], stage1_50[98]},
      {stage1_51[66]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[11],stage2_52[24],stage2_51[52],stage2_50[62]}
   );
   gpc615_5 gpc6890 (
      {stage1_50[99], stage1_50[100], stage1_50[101], stage1_50[102], stage1_50[103]},
      {stage1_51[67]},
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage2_54[6],stage2_53[12],stage2_52[25],stage2_51[53],stage2_50[63]}
   );
   gpc615_5 gpc6891 (
      {stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107], stage1_50[108]},
      {stage1_51[68]},
      {stage1_52[17], stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22]},
      {stage2_54[7],stage2_53[13],stage2_52[26],stage2_51[54],stage2_50[64]}
   );
   gpc615_5 gpc6892 (
      {stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112], stage1_50[113]},
      {stage1_51[69]},
      {stage1_52[23], stage1_52[24], stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28]},
      {stage2_54[8],stage2_53[14],stage2_52[27],stage2_51[55],stage2_50[65]}
   );
   gpc615_5 gpc6893 (
      {stage1_50[114], stage1_50[115], stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[70]},
      {stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34]},
      {stage2_54[9],stage2_53[15],stage2_52[28],stage2_51[56],stage2_50[66]}
   );
   gpc615_5 gpc6894 (
      {stage1_50[119], stage1_50[120], stage1_50[121], stage1_50[122], stage1_50[123]},
      {stage1_51[71]},
      {stage1_52[35], stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40]},
      {stage2_54[10],stage2_53[16],stage2_52[29],stage2_51[57],stage2_50[67]}
   );
   gpc615_5 gpc6895 (
      {stage1_50[124], stage1_50[125], stage1_50[126], stage1_50[127], stage1_50[128]},
      {stage1_51[72]},
      {stage1_52[41], stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46]},
      {stage2_54[11],stage2_53[17],stage2_52[30],stage2_51[58],stage2_50[68]}
   );
   gpc615_5 gpc6896 (
      {stage1_50[129], stage1_50[130], stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[73]},
      {stage1_52[47], stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52]},
      {stage2_54[12],stage2_53[18],stage2_52[31],stage2_51[59],stage2_50[69]}
   );
   gpc606_5 gpc6897 (
      {stage1_51[74], stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79]},
      {stage1_53[5], stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10]},
      {stage2_55[0],stage2_54[13],stage2_53[19],stage2_52[32],stage2_51[60]}
   );
   gpc606_5 gpc6898 (
      {stage1_51[80], stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85]},
      {stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16]},
      {stage2_55[1],stage2_54[14],stage2_53[20],stage2_52[33],stage2_51[61]}
   );
   gpc606_5 gpc6899 (
      {stage1_51[86], stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91]},
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22]},
      {stage2_55[2],stage2_54[15],stage2_53[21],stage2_52[34],stage2_51[62]}
   );
   gpc606_5 gpc6900 (
      {stage1_51[92], stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97]},
      {stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28]},
      {stage2_55[3],stage2_54[16],stage2_53[22],stage2_52[35],stage2_51[63]}
   );
   gpc606_5 gpc6901 (
      {stage1_51[98], stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103]},
      {stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage2_55[4],stage2_54[17],stage2_53[23],stage2_52[36],stage2_51[64]}
   );
   gpc606_5 gpc6902 (
      {stage1_51[104], stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109]},
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40]},
      {stage2_55[5],stage2_54[18],stage2_53[24],stage2_52[37],stage2_51[65]}
   );
   gpc606_5 gpc6903 (
      {stage1_51[110], stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115]},
      {stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46]},
      {stage2_55[6],stage2_54[19],stage2_53[25],stage2_52[38],stage2_51[66]}
   );
   gpc606_5 gpc6904 (
      {stage1_51[116], stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121]},
      {stage1_53[47], stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52]},
      {stage2_55[7],stage2_54[20],stage2_53[26],stage2_52[39],stage2_51[67]}
   );
   gpc606_5 gpc6905 (
      {stage1_51[122], stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127]},
      {stage1_53[53], stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58]},
      {stage2_55[8],stage2_54[21],stage2_53[27],stage2_52[40],stage2_51[68]}
   );
   gpc606_5 gpc6906 (
      {stage1_51[128], stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133]},
      {stage1_53[59], stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64]},
      {stage2_55[9],stage2_54[22],stage2_53[28],stage2_52[41],stage2_51[69]}
   );
   gpc606_5 gpc6907 (
      {stage1_51[134], stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139]},
      {stage1_53[65], stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70]},
      {stage2_55[10],stage2_54[23],stage2_53[29],stage2_52[42],stage2_51[70]}
   );
   gpc606_5 gpc6908 (
      {stage1_51[140], stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145]},
      {stage1_53[71], stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76]},
      {stage2_55[11],stage2_54[24],stage2_53[30],stage2_52[43],stage2_51[71]}
   );
   gpc606_5 gpc6909 (
      {stage1_51[146], stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151]},
      {stage1_53[77], stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82]},
      {stage2_55[12],stage2_54[25],stage2_53[31],stage2_52[44],stage2_51[72]}
   );
   gpc606_5 gpc6910 (
      {stage1_51[152], stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157]},
      {stage1_53[83], stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88]},
      {stage2_55[13],stage2_54[26],stage2_53[32],stage2_52[45],stage2_51[73]}
   );
   gpc606_5 gpc6911 (
      {stage1_51[158], stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163]},
      {stage1_53[89], stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94]},
      {stage2_55[14],stage2_54[27],stage2_53[33],stage2_52[46],stage2_51[74]}
   );
   gpc606_5 gpc6912 (
      {stage1_51[164], stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169]},
      {stage1_53[95], stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100]},
      {stage2_55[15],stage2_54[28],stage2_53[34],stage2_52[47],stage2_51[75]}
   );
   gpc606_5 gpc6913 (
      {stage1_51[170], stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175]},
      {stage1_53[101], stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106]},
      {stage2_55[16],stage2_54[29],stage2_53[35],stage2_52[48],stage2_51[76]}
   );
   gpc606_5 gpc6914 (
      {stage1_51[176], stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181]},
      {stage1_53[107], stage1_53[108], stage1_53[109], stage1_53[110], stage1_53[111], stage1_53[112]},
      {stage2_55[17],stage2_54[30],stage2_53[36],stage2_52[49],stage2_51[77]}
   );
   gpc606_5 gpc6915 (
      {stage1_51[182], stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187]},
      {stage1_53[113], stage1_53[114], stage1_53[115], stage1_53[116], stage1_53[117], stage1_53[118]},
      {stage2_55[18],stage2_54[31],stage2_53[37],stage2_52[50],stage2_51[78]}
   );
   gpc606_5 gpc6916 (
      {stage1_51[188], stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193]},
      {stage1_53[119], stage1_53[120], stage1_53[121], stage1_53[122], stage1_53[123], stage1_53[124]},
      {stage2_55[19],stage2_54[32],stage2_53[38],stage2_52[51],stage2_51[79]}
   );
   gpc606_5 gpc6917 (
      {stage1_51[194], stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199]},
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129], stage1_53[130]},
      {stage2_55[20],stage2_54[33],stage2_53[39],stage2_52[52],stage2_51[80]}
   );
   gpc606_5 gpc6918 (
      {stage1_51[200], stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_53[131], stage1_53[132], stage1_53[133], stage1_53[134], stage1_53[135], stage1_53[136]},
      {stage2_55[21],stage2_54[34],stage2_53[40],stage2_52[53],stage2_51[81]}
   );
   gpc606_5 gpc6919 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210], stage1_51[211]},
      {stage1_53[137], stage1_53[138], stage1_53[139], stage1_53[140], stage1_53[141], stage1_53[142]},
      {stage2_55[22],stage2_54[35],stage2_53[41],stage2_52[54],stage2_51[82]}
   );
   gpc606_5 gpc6920 (
      {stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215], stage1_51[216], stage1_51[217]},
      {stage1_53[143], stage1_53[144], stage1_53[145], stage1_53[146], stage1_53[147], stage1_53[148]},
      {stage2_55[23],stage2_54[36],stage2_53[42],stage2_52[55],stage2_51[83]}
   );
   gpc606_5 gpc6921 (
      {stage1_51[218], stage1_51[219], stage1_51[220], stage1_51[221], stage1_51[222], stage1_51[223]},
      {stage1_53[149], stage1_53[150], stage1_53[151], stage1_53[152], stage1_53[153], stage1_53[154]},
      {stage2_55[24],stage2_54[37],stage2_53[43],stage2_52[56],stage2_51[84]}
   );
   gpc606_5 gpc6922 (
      {stage1_52[53], stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[25],stage2_54[38],stage2_53[44],stage2_52[57]}
   );
   gpc606_5 gpc6923 (
      {stage1_52[59], stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[26],stage2_54[39],stage2_53[45],stage2_52[58]}
   );
   gpc606_5 gpc6924 (
      {stage1_52[65], stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[27],stage2_54[40],stage2_53[46],stage2_52[59]}
   );
   gpc606_5 gpc6925 (
      {stage1_52[71], stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[28],stage2_54[41],stage2_53[47],stage2_52[60]}
   );
   gpc606_5 gpc6926 (
      {stage1_52[77], stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[29],stage2_54[42],stage2_53[48],stage2_52[61]}
   );
   gpc606_5 gpc6927 (
      {stage1_52[83], stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[30],stage2_54[43],stage2_53[49],stage2_52[62]}
   );
   gpc606_5 gpc6928 (
      {stage1_52[89], stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[31],stage2_54[44],stage2_53[50],stage2_52[63]}
   );
   gpc606_5 gpc6929 (
      {stage1_52[95], stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[32],stage2_54[45],stage2_53[51],stage2_52[64]}
   );
   gpc606_5 gpc6930 (
      {stage1_52[101], stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[33],stage2_54[46],stage2_53[52],stage2_52[65]}
   );
   gpc606_5 gpc6931 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111], stage1_52[112]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[34],stage2_54[47],stage2_53[53],stage2_52[66]}
   );
   gpc606_5 gpc6932 (
      {stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116], stage1_52[117], stage1_52[118]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[35],stage2_54[48],stage2_53[54],stage2_52[67]}
   );
   gpc606_5 gpc6933 (
      {stage1_52[119], stage1_52[120], stage1_52[121], stage1_52[122], stage1_52[123], stage1_52[124]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[36],stage2_54[49],stage2_53[55],stage2_52[68]}
   );
   gpc606_5 gpc6934 (
      {stage1_52[125], stage1_52[126], stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[37],stage2_54[50],stage2_53[56],stage2_52[69]}
   );
   gpc606_5 gpc6935 (
      {stage1_52[131], stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[38],stage2_54[51],stage2_53[57],stage2_52[70]}
   );
   gpc606_5 gpc6936 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141], stage1_52[142]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[39],stage2_54[52],stage2_53[58],stage2_52[71]}
   );
   gpc606_5 gpc6937 (
      {stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146], stage1_52[147], stage1_52[148]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[40],stage2_54[53],stage2_53[59],stage2_52[72]}
   );
   gpc606_5 gpc6938 (
      {stage1_52[149], stage1_52[150], stage1_52[151], stage1_52[152], stage1_52[153], stage1_52[154]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[41],stage2_54[54],stage2_53[60],stage2_52[73]}
   );
   gpc606_5 gpc6939 (
      {stage1_52[155], stage1_52[156], stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[42],stage2_54[55],stage2_53[61],stage2_52[74]}
   );
   gpc606_5 gpc6940 (
      {stage1_52[161], stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[43],stage2_54[56],stage2_53[62],stage2_52[75]}
   );
   gpc606_5 gpc6941 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171], stage1_52[172]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[44],stage2_54[57],stage2_53[63],stage2_52[76]}
   );
   gpc606_5 gpc6942 (
      {stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176], stage1_52[177], stage1_52[178]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[45],stage2_54[58],stage2_53[64],stage2_52[77]}
   );
   gpc606_5 gpc6943 (
      {stage1_52[179], stage1_52[180], stage1_52[181], stage1_52[182], stage1_52[183], stage1_52[184]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[46],stage2_54[59],stage2_53[65],stage2_52[78]}
   );
   gpc606_5 gpc6944 (
      {stage1_52[185], stage1_52[186], stage1_52[187], stage1_52[188], stage1_52[189], stage1_52[190]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[47],stage2_54[60],stage2_53[66],stage2_52[79]}
   );
   gpc606_5 gpc6945 (
      {stage1_52[191], stage1_52[192], stage1_52[193], stage1_52[194], stage1_52[195], stage1_52[196]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[48],stage2_54[61],stage2_53[67],stage2_52[80]}
   );
   gpc606_5 gpc6946 (
      {stage1_52[197], stage1_52[198], stage1_52[199], stage1_52[200], stage1_52[201], stage1_52[202]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[49],stage2_54[62],stage2_53[68],stage2_52[81]}
   );
   gpc606_5 gpc6947 (
      {stage1_52[203], stage1_52[204], stage1_52[205], stage1_52[206], stage1_52[207], stage1_52[208]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[50],stage2_54[63],stage2_53[69],stage2_52[82]}
   );
   gpc606_5 gpc6948 (
      {stage1_52[209], stage1_52[210], stage1_52[211], stage1_52[212], stage1_52[213], stage1_52[214]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[51],stage2_54[64],stage2_53[70],stage2_52[83]}
   );
   gpc606_5 gpc6949 (
      {stage1_52[215], stage1_52[216], stage1_52[217], stage1_52[218], stage1_52[219], stage1_52[220]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[52],stage2_54[65],stage2_53[71],stage2_52[84]}
   );
   gpc606_5 gpc6950 (
      {stage1_52[221], stage1_52[222], stage1_52[223], stage1_52[224], stage1_52[225], stage1_52[226]},
      {stage1_54[168], stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173]},
      {stage2_56[28],stage2_55[53],stage2_54[66],stage2_53[72],stage2_52[85]}
   );
   gpc606_5 gpc6951 (
      {stage1_52[227], stage1_52[228], stage1_52[229], stage1_52[230], stage1_52[231], stage1_52[232]},
      {stage1_54[174], stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179]},
      {stage2_56[29],stage2_55[54],stage2_54[67],stage2_53[73],stage2_52[86]}
   );
   gpc606_5 gpc6952 (
      {stage1_52[233], stage1_52[234], stage1_52[235], stage1_52[236], stage1_52[237], stage1_52[238]},
      {stage1_54[180], stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185]},
      {stage2_56[30],stage2_55[55],stage2_54[68],stage2_53[74],stage2_52[87]}
   );
   gpc606_5 gpc6953 (
      {stage1_52[239], stage1_52[240], stage1_52[241], stage1_52[242], stage1_52[243], stage1_52[244]},
      {stage1_54[186], stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191]},
      {stage2_56[31],stage2_55[56],stage2_54[69],stage2_53[75],stage2_52[88]}
   );
   gpc606_5 gpc6954 (
      {stage1_52[245], stage1_52[246], stage1_52[247], stage1_52[248], stage1_52[249], stage1_52[250]},
      {stage1_54[192], stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage2_56[32],stage2_55[57],stage2_54[70],stage2_53[76],stage2_52[89]}
   );
   gpc606_5 gpc6955 (
      {stage1_52[251], stage1_52[252], stage1_52[253], stage1_52[254], stage1_52[255], stage1_52[256]},
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202], stage1_54[203]},
      {stage2_56[33],stage2_55[58],stage2_54[71],stage2_53[77],stage2_52[90]}
   );
   gpc606_5 gpc6956 (
      {stage1_52[257], stage1_52[258], stage1_52[259], stage1_52[260], stage1_52[261], stage1_52[262]},
      {stage1_54[204], stage1_54[205], stage1_54[206], stage1_54[207], stage1_54[208], stage1_54[209]},
      {stage2_56[34],stage2_55[59],stage2_54[72],stage2_53[78],stage2_52[91]}
   );
   gpc606_5 gpc6957 (
      {stage1_52[263], stage1_52[264], stage1_52[265], stage1_52[266], stage1_52[267], stage1_52[268]},
      {stage1_54[210], stage1_54[211], stage1_54[212], stage1_54[213], stage1_54[214], stage1_54[215]},
      {stage2_56[35],stage2_55[60],stage2_54[73],stage2_53[79],stage2_52[92]}
   );
   gpc606_5 gpc6958 (
      {stage1_53[155], stage1_53[156], stage1_53[157], stage1_53[158], stage1_53[159], stage1_53[160]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[36],stage2_55[61],stage2_54[74],stage2_53[80]}
   );
   gpc606_5 gpc6959 (
      {stage1_53[161], stage1_53[162], stage1_53[163], stage1_53[164], stage1_53[165], stage1_53[166]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[37],stage2_55[62],stage2_54[75],stage2_53[81]}
   );
   gpc606_5 gpc6960 (
      {stage1_53[167], stage1_53[168], stage1_53[169], stage1_53[170], stage1_53[171], stage1_53[172]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[38],stage2_55[63],stage2_54[76],stage2_53[82]}
   );
   gpc2135_5 gpc6961 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[0], stage1_56[1], stage1_56[2]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[0],stage2_57[3],stage2_56[39],stage2_55[64]}
   );
   gpc2135_5 gpc6962 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[1],stage2_57[4],stage2_56[40],stage2_55[65]}
   );
   gpc2135_5 gpc6963 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[6], stage1_56[7], stage1_56[8]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[2],stage2_57[5],stage2_56[41],stage2_55[66]}
   );
   gpc2135_5 gpc6964 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[3],stage2_57[6],stage2_56[42],stage2_55[67]}
   );
   gpc2135_5 gpc6965 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12], stage1_56[13], stage1_56[14]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[4],stage2_57[7],stage2_56[43],stage2_55[68]}
   );
   gpc2135_5 gpc6966 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[5],stage2_57[8],stage2_56[44],stage2_55[69]}
   );
   gpc2135_5 gpc6967 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[18], stage1_56[19], stage1_56[20]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[6],stage2_57[9],stage2_56[45],stage2_55[70]}
   );
   gpc2135_5 gpc6968 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[7],stage2_57[10],stage2_56[46],stage2_55[71]}
   );
   gpc2135_5 gpc6969 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[24], stage1_56[25], stage1_56[26]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[8],stage2_57[11],stage2_56[47],stage2_55[72]}
   );
   gpc2135_5 gpc6970 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[9],stage2_57[12],stage2_56[48],stage2_55[73]}
   );
   gpc2135_5 gpc6971 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[30], stage1_56[31], stage1_56[32]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[10],stage2_57[13],stage2_56[49],stage2_55[74]}
   );
   gpc2135_5 gpc6972 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[11],stage2_57[14],stage2_56[50],stage2_55[75]}
   );
   gpc2135_5 gpc6973 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[12],stage2_57[15],stage2_56[51],stage2_55[76]}
   );
   gpc2135_5 gpc6974 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[13],stage2_57[16],stage2_56[52],stage2_55[77]}
   );
   gpc2135_5 gpc6975 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[14],stage2_57[17],stage2_56[53],stage2_55[78]}
   );
   gpc2135_5 gpc6976 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[15],stage2_57[18],stage2_56[54],stage2_55[79]}
   );
   gpc2135_5 gpc6977 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[16],stage2_57[19],stage2_56[55],stage2_55[80]}
   );
   gpc2135_5 gpc6978 (
      {stage1_55[103], stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[17],stage2_57[20],stage2_56[56],stage2_55[81]}
   );
   gpc2135_5 gpc6979 (
      {stage1_55[108], stage1_55[109], stage1_55[110], stage1_55[111], stage1_55[112]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[18]},
      {stage1_58[36], stage1_58[37]},
      {stage2_59[18],stage2_58[18],stage2_57[21],stage2_56[57],stage2_55[82]}
   );
   gpc2135_5 gpc6980 (
      {stage1_55[113], stage1_55[114], stage1_55[115], stage1_55[116], stage1_55[117]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[19]},
      {stage1_58[38], stage1_58[39]},
      {stage2_59[19],stage2_58[19],stage2_57[22],stage2_56[58],stage2_55[83]}
   );
   gpc2135_5 gpc6981 (
      {stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121], stage1_55[122]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[20]},
      {stage1_58[40], stage1_58[41]},
      {stage2_59[20],stage2_58[20],stage2_57[23],stage2_56[59],stage2_55[84]}
   );
   gpc2135_5 gpc6982 (
      {stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[21]},
      {stage1_58[42], stage1_58[43]},
      {stage2_59[21],stage2_58[21],stage2_57[24],stage2_56[60],stage2_55[85]}
   );
   gpc2135_5 gpc6983 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[22]},
      {stage1_58[44], stage1_58[45]},
      {stage2_59[22],stage2_58[22],stage2_57[25],stage2_56[61],stage2_55[86]}
   );
   gpc2135_5 gpc6984 (
      {stage1_55[133], stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[23]},
      {stage1_58[46], stage1_58[47]},
      {stage2_59[23],stage2_58[23],stage2_57[26],stage2_56[62],stage2_55[87]}
   );
   gpc2135_5 gpc6985 (
      {stage1_55[138], stage1_55[139], stage1_55[140], stage1_55[141], stage1_55[142]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[24]},
      {stage1_58[48], stage1_58[49]},
      {stage2_59[24],stage2_58[24],stage2_57[27],stage2_56[63],stage2_55[88]}
   );
   gpc2135_5 gpc6986 (
      {stage1_55[143], stage1_55[144], stage1_55[145], stage1_55[146], stage1_55[147]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[25]},
      {stage1_58[50], stage1_58[51]},
      {stage2_59[25],stage2_58[25],stage2_57[28],stage2_56[64],stage2_55[89]}
   );
   gpc2135_5 gpc6987 (
      {stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151], stage1_55[152]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[26]},
      {stage1_58[52], stage1_58[53]},
      {stage2_59[26],stage2_58[26],stage2_57[29],stage2_56[65],stage2_55[90]}
   );
   gpc2135_5 gpc6988 (
      {stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[27]},
      {stage1_58[54], stage1_58[55]},
      {stage2_59[27],stage2_58[27],stage2_57[30],stage2_56[66],stage2_55[91]}
   );
   gpc2135_5 gpc6989 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[28]},
      {stage1_58[56], stage1_58[57]},
      {stage2_59[28],stage2_58[28],stage2_57[31],stage2_56[67],stage2_55[92]}
   );
   gpc2135_5 gpc6990 (
      {stage1_55[163], stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[29]},
      {stage1_58[58], stage1_58[59]},
      {stage2_59[29],stage2_58[29],stage2_57[32],stage2_56[68],stage2_55[93]}
   );
   gpc606_5 gpc6991 (
      {stage1_55[168], stage1_55[169], stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[30],stage2_58[30],stage2_57[33],stage2_56[69],stage2_55[94]}
   );
   gpc615_5 gpc6992 (
      {stage1_55[174], stage1_55[175], stage1_55[176], stage1_55[177], stage1_55[178]},
      {stage1_56[90]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[31],stage2_58[31],stage2_57[34],stage2_56[70],stage2_55[95]}
   );
   gpc615_5 gpc6993 (
      {stage1_55[179], stage1_55[180], stage1_55[181], stage1_55[182], stage1_55[183]},
      {stage1_56[91]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[32],stage2_58[32],stage2_57[35],stage2_56[71],stage2_55[96]}
   );
   gpc615_5 gpc6994 (
      {stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187], stage1_55[188]},
      {stage1_56[92]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[33],stage2_58[33],stage2_57[36],stage2_56[72],stage2_55[97]}
   );
   gpc615_5 gpc6995 (
      {stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_56[93]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[34],stage2_58[34],stage2_57[37],stage2_56[73],stage2_55[98]}
   );
   gpc615_5 gpc6996 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198]},
      {stage1_56[94]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[35],stage2_58[35],stage2_57[38],stage2_56[74],stage2_55[99]}
   );
   gpc615_5 gpc6997 (
      {stage1_55[199], stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203]},
      {stage1_56[95]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[36],stage2_58[36],stage2_57[39],stage2_56[75],stage2_55[100]}
   );
   gpc615_5 gpc6998 (
      {stage1_55[204], stage1_55[205], stage1_55[206], stage1_55[207], stage1_55[208]},
      {stage1_56[96]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[37],stage2_58[37],stage2_57[40],stage2_56[76],stage2_55[101]}
   );
   gpc615_5 gpc6999 (
      {stage1_55[209], stage1_55[210], stage1_55[211], stage1_55[212], stage1_55[213]},
      {stage1_56[97]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[38],stage2_58[38],stage2_57[41],stage2_56[77],stage2_55[102]}
   );
   gpc615_5 gpc7000 (
      {stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217], stage1_55[218]},
      {stage1_56[98]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[39],stage2_58[39],stage2_57[42],stage2_56[78],stage2_55[103]}
   );
   gpc606_5 gpc7001 (
      {stage1_56[99], stage1_56[100], stage1_56[101], stage1_56[102], stage1_56[103], stage1_56[104]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[0],stage2_59[40],stage2_58[40],stage2_57[43],stage2_56[79]}
   );
   gpc606_5 gpc7002 (
      {stage1_56[105], stage1_56[106], stage1_56[107], stage1_56[108], stage1_56[109], stage1_56[110]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[1],stage2_59[41],stage2_58[41],stage2_57[44],stage2_56[80]}
   );
   gpc606_5 gpc7003 (
      {stage1_56[111], stage1_56[112], stage1_56[113], stage1_56[114], stage1_56[115], stage1_56[116]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[2],stage2_59[42],stage2_58[42],stage2_57[45],stage2_56[81]}
   );
   gpc606_5 gpc7004 (
      {stage1_56[117], stage1_56[118], stage1_56[119], stage1_56[120], stage1_56[121], stage1_56[122]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[3],stage2_59[43],stage2_58[43],stage2_57[46],stage2_56[82]}
   );
   gpc606_5 gpc7005 (
      {stage1_56[123], stage1_56[124], stage1_56[125], stage1_56[126], stage1_56[127], stage1_56[128]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[4],stage2_59[44],stage2_58[44],stage2_57[47],stage2_56[83]}
   );
   gpc606_5 gpc7006 (
      {stage1_56[129], stage1_56[130], stage1_56[131], stage1_56[132], stage1_56[133], stage1_56[134]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[5],stage2_59[45],stage2_58[45],stage2_57[48],stage2_56[84]}
   );
   gpc606_5 gpc7007 (
      {stage1_56[135], stage1_56[136], stage1_56[137], stage1_56[138], stage1_56[139], stage1_56[140]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[6],stage2_59[46],stage2_58[46],stage2_57[49],stage2_56[85]}
   );
   gpc606_5 gpc7008 (
      {stage1_56[141], stage1_56[142], stage1_56[143], stage1_56[144], stage1_56[145], stage1_56[146]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[7],stage2_59[47],stage2_58[47],stage2_57[50],stage2_56[86]}
   );
   gpc606_5 gpc7009 (
      {stage1_56[147], stage1_56[148], stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[8],stage2_59[48],stage2_58[48],stage2_57[51],stage2_56[87]}
   );
   gpc606_5 gpc7010 (
      {stage1_56[153], stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_58[114], stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage2_60[9],stage2_59[49],stage2_58[49],stage2_57[52],stage2_56[88]}
   );
   gpc606_5 gpc7011 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163], stage1_56[164]},
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124], stage1_58[125]},
      {stage2_60[10],stage2_59[50],stage2_58[50],stage2_57[53],stage2_56[89]}
   );
   gpc606_5 gpc7012 (
      {stage1_56[165], stage1_56[166], stage1_56[167], stage1_56[168], stage1_56[169], stage1_56[170]},
      {stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129], stage1_58[130], stage1_58[131]},
      {stage2_60[11],stage2_59[51],stage2_58[51],stage2_57[54],stage2_56[90]}
   );
   gpc606_5 gpc7013 (
      {stage1_56[171], stage1_56[172], stage1_56[173], stage1_56[174], stage1_56[175], stage1_56[176]},
      {stage1_58[132], stage1_58[133], stage1_58[134], stage1_58[135], stage1_58[136], stage1_58[137]},
      {stage2_60[12],stage2_59[52],stage2_58[52],stage2_57[55],stage2_56[91]}
   );
   gpc606_5 gpc7014 (
      {stage1_56[177], stage1_56[178], stage1_56[179], stage1_56[180], stage1_56[181], stage1_56[182]},
      {stage1_58[138], stage1_58[139], stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143]},
      {stage2_60[13],stage2_59[53],stage2_58[53],stage2_57[56],stage2_56[92]}
   );
   gpc606_5 gpc7015 (
      {stage1_56[183], stage1_56[184], stage1_56[185], stage1_56[186], stage1_56[187], stage1_56[188]},
      {stage1_58[144], stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage2_60[14],stage2_59[54],stage2_58[54],stage2_57[57],stage2_56[93]}
   );
   gpc606_5 gpc7016 (
      {stage1_56[189], stage1_56[190], stage1_56[191], stage1_56[192], stage1_56[193], stage1_56[194]},
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154], stage1_58[155]},
      {stage2_60[15],stage2_59[55],stage2_58[55],stage2_57[58],stage2_56[94]}
   );
   gpc606_5 gpc7017 (
      {stage1_56[195], stage1_56[196], stage1_56[197], stage1_56[198], stage1_56[199], stage1_56[200]},
      {stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159], stage1_58[160], stage1_58[161]},
      {stage2_60[16],stage2_59[56],stage2_58[56],stage2_57[59],stage2_56[95]}
   );
   gpc606_5 gpc7018 (
      {stage1_56[201], stage1_56[202], stage1_56[203], stage1_56[204], stage1_56[205], stage1_56[206]},
      {stage1_58[162], stage1_58[163], stage1_58[164], stage1_58[165], stage1_58[166], stage1_58[167]},
      {stage2_60[17],stage2_59[57],stage2_58[57],stage2_57[60],stage2_56[96]}
   );
   gpc606_5 gpc7019 (
      {stage1_56[207], stage1_56[208], stage1_56[209], stage1_56[210], stage1_56[211], stage1_56[212]},
      {stage1_58[168], stage1_58[169], stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173]},
      {stage2_60[18],stage2_59[58],stage2_58[58],stage2_57[61],stage2_56[97]}
   );
   gpc606_5 gpc7020 (
      {stage1_56[213], stage1_56[214], stage1_56[215], stage1_56[216], stage1_56[217], stage1_56[218]},
      {stage1_58[174], stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage2_60[19],stage2_59[59],stage2_58[59],stage2_57[62],stage2_56[98]}
   );
   gpc606_5 gpc7021 (
      {stage1_56[219], stage1_56[220], stage1_56[221], stage1_56[222], stage1_56[223], stage1_56[224]},
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184], stage1_58[185]},
      {stage2_60[20],stage2_59[60],stage2_58[60],stage2_57[63],stage2_56[99]}
   );
   gpc606_5 gpc7022 (
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[21],stage2_59[61],stage2_58[61],stage2_57[64]}
   );
   gpc606_5 gpc7023 (
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[22],stage2_59[62],stage2_58[62],stage2_57[65]}
   );
   gpc606_5 gpc7024 (
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[23],stage2_59[63],stage2_58[63],stage2_57[66]}
   );
   gpc606_5 gpc7025 (
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[24],stage2_59[64],stage2_58[64],stage2_57[67]}
   );
   gpc606_5 gpc7026 (
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage2_61[4],stage2_60[25],stage2_59[65],stage2_58[65],stage2_57[68]}
   );
   gpc606_5 gpc7027 (
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage2_61[5],stage2_60[26],stage2_59[66],stage2_58[66],stage2_57[69]}
   );
   gpc606_5 gpc7028 (
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage2_61[6],stage2_60[27],stage2_59[67],stage2_58[67],stage2_57[70]}
   );
   gpc606_5 gpc7029 (
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage1_59[42], stage1_59[43], stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47]},
      {stage2_61[7],stage2_60[28],stage2_59[68],stage2_58[68],stage2_57[71]}
   );
   gpc606_5 gpc7030 (
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage1_59[48], stage1_59[49], stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53]},
      {stage2_61[8],stage2_60[29],stage2_59[69],stage2_58[69],stage2_57[72]}
   );
   gpc606_5 gpc7031 (
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage1_59[54], stage1_59[55], stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59]},
      {stage2_61[9],stage2_60[30],stage2_59[70],stage2_58[70],stage2_57[73]}
   );
   gpc606_5 gpc7032 (
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage1_59[60], stage1_59[61], stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65]},
      {stage2_61[10],stage2_60[31],stage2_59[71],stage2_58[71],stage2_57[74]}
   );
   gpc606_5 gpc7033 (
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage1_59[66], stage1_59[67], stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71]},
      {stage2_61[11],stage2_60[32],stage2_59[72],stage2_58[72],stage2_57[75]}
   );
   gpc606_5 gpc7034 (
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage1_59[72], stage1_59[73], stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77]},
      {stage2_61[12],stage2_60[33],stage2_59[73],stage2_58[73],stage2_57[76]}
   );
   gpc606_5 gpc7035 (
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage1_59[78], stage1_59[79], stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83]},
      {stage2_61[13],stage2_60[34],stage2_59[74],stage2_58[74],stage2_57[77]}
   );
   gpc606_5 gpc7036 (
      {stage1_57[174], stage1_57[175], stage1_57[176], stage1_57[177], stage1_57[178], stage1_57[179]},
      {stage1_59[84], stage1_59[85], stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89]},
      {stage2_61[14],stage2_60[35],stage2_59[75],stage2_58[75],stage2_57[78]}
   );
   gpc117_4 gpc7037 (
      {stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189], stage1_58[190], stage1_58[191], stage1_58[192]},
      {stage1_59[90]},
      {stage1_60[0]},
      {stage2_61[15],stage2_60[36],stage2_59[76],stage2_58[76]}
   );
   gpc117_4 gpc7038 (
      {stage1_58[193], stage1_58[194], stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[91]},
      {stage1_60[1]},
      {stage2_61[16],stage2_60[37],stage2_59[77],stage2_58[77]}
   );
   gpc117_4 gpc7039 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204], stage1_58[205], stage1_58[206]},
      {stage1_59[92]},
      {stage1_60[2]},
      {stage2_61[17],stage2_60[38],stage2_59[78],stage2_58[78]}
   );
   gpc117_4 gpc7040 (
      {stage1_58[207], stage1_58[208], stage1_58[209], stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213]},
      {stage1_59[93]},
      {stage1_60[3]},
      {stage2_61[18],stage2_60[39],stage2_59[79],stage2_58[79]}
   );
   gpc606_5 gpc7041 (
      {stage1_58[214], stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_60[4], stage1_60[5], stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9]},
      {stage2_62[0],stage2_61[19],stage2_60[40],stage2_59[80],stage2_58[80]}
   );
   gpc606_5 gpc7042 (
      {stage1_58[220], stage1_58[221], stage1_58[222], stage1_58[223], stage1_58[224], stage1_58[225]},
      {stage1_60[10], stage1_60[11], stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15]},
      {stage2_62[1],stage2_61[20],stage2_60[41],stage2_59[81],stage2_58[81]}
   );
   gpc606_5 gpc7043 (
      {stage1_58[226], stage1_58[227], stage1_58[228], stage1_58[229], stage1_58[230], stage1_58[231]},
      {stage1_60[16], stage1_60[17], stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21]},
      {stage2_62[2],stage2_61[21],stage2_60[42],stage2_59[82],stage2_58[82]}
   );
   gpc606_5 gpc7044 (
      {stage1_58[232], stage1_58[233], stage1_58[234], stage1_58[235], stage1_58[236], stage1_58[237]},
      {stage1_60[22], stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage2_62[3],stage2_61[22],stage2_60[43],stage2_59[83],stage2_58[83]}
   );
   gpc606_5 gpc7045 (
      {stage1_58[238], stage1_58[239], stage1_58[240], stage1_58[241], stage1_58[242], 1'b0},
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33]},
      {stage2_62[4],stage2_61[23],stage2_60[44],stage2_59[84],stage2_58[84]}
   );
   gpc606_5 gpc7046 (
      {stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97], stage1_59[98], stage1_59[99]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[24],stage2_60[45],stage2_59[85]}
   );
   gpc606_5 gpc7047 (
      {stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103], stage1_59[104], stage1_59[105]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[25],stage2_60[46],stage2_59[86]}
   );
   gpc606_5 gpc7048 (
      {stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109], stage1_59[110], stage1_59[111]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[26],stage2_60[47],stage2_59[87]}
   );
   gpc606_5 gpc7049 (
      {stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115], stage1_59[116], stage1_59[117]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[27],stage2_60[48],stage2_59[88]}
   );
   gpc606_5 gpc7050 (
      {stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121], stage1_59[122], stage1_59[123]},
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage2_63[4],stage2_62[9],stage2_61[28],stage2_60[49],stage2_59[89]}
   );
   gpc606_5 gpc7051 (
      {stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127], stage1_59[128], stage1_59[129]},
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage2_63[5],stage2_62[10],stage2_61[29],stage2_60[50],stage2_59[90]}
   );
   gpc606_5 gpc7052 (
      {stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133], stage1_59[134], stage1_59[135]},
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage2_63[6],stage2_62[11],stage2_61[30],stage2_60[51],stage2_59[91]}
   );
   gpc606_5 gpc7053 (
      {stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139], stage1_59[140], stage1_59[141]},
      {stage1_61[42], stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage2_63[7],stage2_62[12],stage2_61[31],stage2_60[52],stage2_59[92]}
   );
   gpc606_5 gpc7054 (
      {stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145], stage1_59[146], stage1_59[147]},
      {stage1_61[48], stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53]},
      {stage2_63[8],stage2_62[13],stage2_61[32],stage2_60[53],stage2_59[93]}
   );
   gpc606_5 gpc7055 (
      {stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151], stage1_59[152], stage1_59[153]},
      {stage1_61[54], stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59]},
      {stage2_63[9],stage2_62[14],stage2_61[33],stage2_60[54],stage2_59[94]}
   );
   gpc606_5 gpc7056 (
      {stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157], stage1_59[158], stage1_59[159]},
      {stage1_61[60], stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65]},
      {stage2_63[10],stage2_62[15],stage2_61[34],stage2_60[55],stage2_59[95]}
   );
   gpc606_5 gpc7057 (
      {stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163], stage1_59[164], stage1_59[165]},
      {stage1_61[66], stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71]},
      {stage2_63[11],stage2_62[16],stage2_61[35],stage2_60[56],stage2_59[96]}
   );
   gpc606_5 gpc7058 (
      {stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169], stage1_59[170], stage1_59[171]},
      {stage1_61[72], stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77]},
      {stage2_63[12],stage2_62[17],stage2_61[36],stage2_60[57],stage2_59[97]}
   );
   gpc606_5 gpc7059 (
      {stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175], stage1_59[176], stage1_59[177]},
      {stage1_61[78], stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83]},
      {stage2_63[13],stage2_62[18],stage2_61[37],stage2_60[58],stage2_59[98]}
   );
   gpc606_5 gpc7060 (
      {stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181], stage1_59[182], stage1_59[183]},
      {stage1_61[84], stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89]},
      {stage2_63[14],stage2_62[19],stage2_61[38],stage2_60[59],stage2_59[99]}
   );
   gpc606_5 gpc7061 (
      {stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187], stage1_59[188], stage1_59[189]},
      {stage1_61[90], stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95]},
      {stage2_63[15],stage2_62[20],stage2_61[39],stage2_60[60],stage2_59[100]}
   );
   gpc606_5 gpc7062 (
      {stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193], stage1_59[194], stage1_59[195]},
      {stage1_61[96], stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101]},
      {stage2_63[16],stage2_62[21],stage2_61[40],stage2_60[61],stage2_59[101]}
   );
   gpc606_5 gpc7063 (
      {stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199], stage1_59[200], stage1_59[201]},
      {stage1_61[102], stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107]},
      {stage2_63[17],stage2_62[22],stage2_61[41],stage2_60[62],stage2_59[102]}
   );
   gpc606_5 gpc7064 (
      {stage1_59[202], stage1_59[203], stage1_59[204], stage1_59[205], stage1_59[206], stage1_59[207]},
      {stage1_61[108], stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113]},
      {stage2_63[18],stage2_62[23],stage2_61[42],stage2_60[63],stage2_59[103]}
   );
   gpc606_5 gpc7065 (
      {stage1_59[208], stage1_59[209], stage1_59[210], stage1_59[211], stage1_59[212], stage1_59[213]},
      {stage1_61[114], stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119]},
      {stage2_63[19],stage2_62[24],stage2_61[43],stage2_60[64],stage2_59[104]}
   );
   gpc606_5 gpc7066 (
      {stage1_59[214], stage1_59[215], stage1_59[216], stage1_59[217], stage1_59[218], stage1_59[219]},
      {stage1_61[120], stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125]},
      {stage2_63[20],stage2_62[25],stage2_61[44],stage2_60[65],stage2_59[105]}
   );
   gpc606_5 gpc7067 (
      {stage1_59[220], stage1_59[221], stage1_59[222], stage1_59[223], stage1_59[224], stage1_59[225]},
      {stage1_61[126], stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131]},
      {stage2_63[21],stage2_62[26],stage2_61[45],stage2_60[66],stage2_59[106]}
   );
   gpc606_5 gpc7068 (
      {stage1_59[226], stage1_59[227], stage1_59[228], stage1_59[229], stage1_59[230], stage1_59[231]},
      {stage1_61[132], stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137]},
      {stage2_63[22],stage2_62[27],stage2_61[46],stage2_60[67],stage2_59[107]}
   );
   gpc606_5 gpc7069 (
      {stage1_59[232], stage1_59[233], stage1_59[234], stage1_59[235], stage1_59[236], stage1_59[237]},
      {stage1_61[138], stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143]},
      {stage2_63[23],stage2_62[28],stage2_61[47],stage2_60[68],stage2_59[108]}
   );
   gpc606_5 gpc7070 (
      {stage1_59[238], stage1_59[239], stage1_59[240], stage1_59[241], stage1_59[242], stage1_59[243]},
      {stage1_61[144], stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149]},
      {stage2_63[24],stage2_62[29],stage2_61[48],stage2_60[69],stage2_59[109]}
   );
   gpc606_5 gpc7071 (
      {stage1_59[244], stage1_59[245], stage1_59[246], stage1_59[247], stage1_59[248], stage1_59[249]},
      {stage1_61[150], stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155]},
      {stage2_63[25],stage2_62[30],stage2_61[49],stage2_60[70],stage2_59[110]}
   );
   gpc606_5 gpc7072 (
      {stage1_59[250], stage1_59[251], stage1_59[252], stage1_59[253], stage1_59[254], stage1_59[255]},
      {stage1_61[156], stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161]},
      {stage2_63[26],stage2_62[31],stage2_61[50],stage2_60[71],stage2_59[111]}
   );
   gpc606_5 gpc7073 (
      {stage1_59[256], stage1_59[257], stage1_59[258], stage1_59[259], stage1_59[260], stage1_59[261]},
      {stage1_61[162], stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167]},
      {stage2_63[27],stage2_62[32],stage2_61[51],stage2_60[72],stage2_59[112]}
   );
   gpc606_5 gpc7074 (
      {stage1_59[262], stage1_59[263], stage1_59[264], stage1_59[265], stage1_59[266], stage1_59[267]},
      {stage1_61[168], stage1_61[169], stage1_61[170], stage1_61[171], stage1_61[172], stage1_61[173]},
      {stage2_63[28],stage2_62[33],stage2_61[52],stage2_60[73],stage2_59[113]}
   );
   gpc1406_5 gpc7075 (
      {stage1_60[34], stage1_60[35], stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3]},
      {stage1_63[0]},
      {stage2_64[0],stage2_63[29],stage2_62[34],stage2_61[53],stage2_60[74]}
   );
   gpc606_5 gpc7076 (
      {stage1_60[40], stage1_60[41], stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45]},
      {stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9]},
      {stage2_64[1],stage2_63[30],stage2_62[35],stage2_61[54],stage2_60[75]}
   );
   gpc606_5 gpc7077 (
      {stage1_60[46], stage1_60[47], stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51]},
      {stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15]},
      {stage2_64[2],stage2_63[31],stage2_62[36],stage2_61[55],stage2_60[76]}
   );
   gpc606_5 gpc7078 (
      {stage1_60[52], stage1_60[53], stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57]},
      {stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21]},
      {stage2_64[3],stage2_63[32],stage2_62[37],stage2_61[56],stage2_60[77]}
   );
   gpc606_5 gpc7079 (
      {stage1_60[58], stage1_60[59], stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63]},
      {stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27]},
      {stage2_64[4],stage2_63[33],stage2_62[38],stage2_61[57],stage2_60[78]}
   );
   gpc606_5 gpc7080 (
      {stage1_60[64], stage1_60[65], stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69]},
      {stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33]},
      {stage2_64[5],stage2_63[34],stage2_62[39],stage2_61[58],stage2_60[79]}
   );
   gpc606_5 gpc7081 (
      {stage1_60[70], stage1_60[71], stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75]},
      {stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39]},
      {stage2_64[6],stage2_63[35],stage2_62[40],stage2_61[59],stage2_60[80]}
   );
   gpc606_5 gpc7082 (
      {stage1_60[76], stage1_60[77], stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81]},
      {stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage2_64[7],stage2_63[36],stage2_62[41],stage2_61[60],stage2_60[81]}
   );
   gpc606_5 gpc7083 (
      {stage1_60[82], stage1_60[83], stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87]},
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51]},
      {stage2_64[8],stage2_63[37],stage2_62[42],stage2_61[61],stage2_60[82]}
   );
   gpc606_5 gpc7084 (
      {stage1_60[88], stage1_60[89], stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93]},
      {stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57]},
      {stage2_64[9],stage2_63[38],stage2_62[43],stage2_61[62],stage2_60[83]}
   );
   gpc606_5 gpc7085 (
      {stage1_60[94], stage1_60[95], stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99]},
      {stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63]},
      {stage2_64[10],stage2_63[39],stage2_62[44],stage2_61[63],stage2_60[84]}
   );
   gpc606_5 gpc7086 (
      {stage1_60[100], stage1_60[101], stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105]},
      {stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69]},
      {stage2_64[11],stage2_63[40],stage2_62[45],stage2_61[64],stage2_60[85]}
   );
   gpc606_5 gpc7087 (
      {stage1_60[106], stage1_60[107], stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111]},
      {stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75]},
      {stage2_64[12],stage2_63[41],stage2_62[46],stage2_61[65],stage2_60[86]}
   );
   gpc606_5 gpc7088 (
      {stage1_60[112], stage1_60[113], stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117]},
      {stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79], stage1_62[80], stage1_62[81]},
      {stage2_64[13],stage2_63[42],stage2_62[47],stage2_61[66],stage2_60[87]}
   );
   gpc606_5 gpc7089 (
      {stage1_60[118], stage1_60[119], stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123]},
      {stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85], stage1_62[86], stage1_62[87]},
      {stage2_64[14],stage2_63[43],stage2_62[48],stage2_61[67],stage2_60[88]}
   );
   gpc606_5 gpc7090 (
      {stage1_60[124], stage1_60[125], stage1_60[126], stage1_60[127], stage1_60[128], stage1_60[129]},
      {stage1_62[88], stage1_62[89], stage1_62[90], stage1_62[91], stage1_62[92], stage1_62[93]},
      {stage2_64[15],stage2_63[44],stage2_62[49],stage2_61[68],stage2_60[89]}
   );
   gpc606_5 gpc7091 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[94], stage1_62[95], stage1_62[96], stage1_62[97], stage1_62[98], stage1_62[99]},
      {stage2_64[16],stage2_63[45],stage2_62[50],stage2_61[69],stage2_60[90]}
   );
   gpc606_5 gpc7092 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[100], stage1_62[101], stage1_62[102], stage1_62[103], stage1_62[104], stage1_62[105]},
      {stage2_64[17],stage2_63[46],stage2_62[51],stage2_61[70],stage2_60[91]}
   );
   gpc606_5 gpc7093 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[106], stage1_62[107], stage1_62[108], stage1_62[109], stage1_62[110], stage1_62[111]},
      {stage2_64[18],stage2_63[47],stage2_62[52],stage2_61[71],stage2_60[92]}
   );
   gpc606_5 gpc7094 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[112], stage1_62[113], stage1_62[114], stage1_62[115], stage1_62[116], stage1_62[117]},
      {stage2_64[19],stage2_63[48],stage2_62[53],stage2_61[72],stage2_60[93]}
   );
   gpc606_5 gpc7095 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[118], stage1_62[119], stage1_62[120], stage1_62[121], stage1_62[122], stage1_62[123]},
      {stage2_64[20],stage2_63[49],stage2_62[54],stage2_61[73],stage2_60[94]}
   );
   gpc615_5 gpc7096 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164]},
      {stage1_61[174]},
      {stage1_62[124], stage1_62[125], stage1_62[126], stage1_62[127], stage1_62[128], stage1_62[129]},
      {stage2_64[21],stage2_63[50],stage2_62[55],stage2_61[74],stage2_60[95]}
   );
   gpc615_5 gpc7097 (
      {stage1_60[165], stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169]},
      {stage1_61[175]},
      {stage1_62[130], stage1_62[131], stage1_62[132], stage1_62[133], stage1_62[134], stage1_62[135]},
      {stage2_64[22],stage2_63[51],stage2_62[56],stage2_61[75],stage2_60[96]}
   );
   gpc615_5 gpc7098 (
      {stage1_60[170], stage1_60[171], stage1_60[172], stage1_60[173], stage1_60[174]},
      {stage1_61[176]},
      {stage1_62[136], stage1_62[137], stage1_62[138], stage1_62[139], stage1_62[140], stage1_62[141]},
      {stage2_64[23],stage2_63[52],stage2_62[57],stage2_61[76],stage2_60[97]}
   );
   gpc615_5 gpc7099 (
      {stage1_60[175], stage1_60[176], stage1_60[177], stage1_60[178], stage1_60[179]},
      {stage1_61[177]},
      {stage1_62[142], stage1_62[143], stage1_62[144], stage1_62[145], stage1_62[146], stage1_62[147]},
      {stage2_64[24],stage2_63[53],stage2_62[58],stage2_61[77],stage2_60[98]}
   );
   gpc615_5 gpc7100 (
      {stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183], stage1_60[184]},
      {stage1_61[178]},
      {stage1_62[148], stage1_62[149], stage1_62[150], stage1_62[151], stage1_62[152], stage1_62[153]},
      {stage2_64[25],stage2_63[54],stage2_62[59],stage2_61[78],stage2_60[99]}
   );
   gpc615_5 gpc7101 (
      {stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188], stage1_60[189]},
      {stage1_61[179]},
      {stage1_62[154], stage1_62[155], stage1_62[156], stage1_62[157], stage1_62[158], stage1_62[159]},
      {stage2_64[26],stage2_63[55],stage2_62[60],stage2_61[79],stage2_60[100]}
   );
   gpc606_5 gpc7102 (
      {stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183], stage1_61[184], stage1_61[185]},
      {stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6]},
      {stage2_65[0],stage2_64[27],stage2_63[56],stage2_62[61],stage2_61[80]}
   );
   gpc606_5 gpc7103 (
      {stage1_61[186], stage1_61[187], stage1_61[188], stage1_61[189], stage1_61[190], stage1_61[191]},
      {stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12]},
      {stage2_65[1],stage2_64[28],stage2_63[57],stage2_62[62],stage2_61[81]}
   );
   gpc606_5 gpc7104 (
      {stage1_61[192], stage1_61[193], stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197]},
      {stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18]},
      {stage2_65[2],stage2_64[29],stage2_63[58],stage2_62[63],stage2_61[82]}
   );
   gpc1163_5 gpc7105 (
      {stage1_62[160], stage1_62[161], stage1_62[162]},
      {stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[3],stage2_64[30],stage2_63[59],stage2_62[64]}
   );
   gpc1163_5 gpc7106 (
      {stage1_62[163], stage1_62[164], stage1_62[165]},
      {stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29], stage1_63[30]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[4],stage2_64[31],stage2_63[60],stage2_62[65]}
   );
   gpc1163_5 gpc7107 (
      {stage1_62[166], stage1_62[167], stage1_62[168]},
      {stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35], stage1_63[36]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[5],stage2_64[32],stage2_63[61],stage2_62[66]}
   );
   gpc1163_5 gpc7108 (
      {stage1_62[169], stage1_62[170], stage1_62[171]},
      {stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41], stage1_63[42]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[6],stage2_64[33],stage2_63[62],stage2_62[67]}
   );
   gpc1163_5 gpc7109 (
      {stage1_62[172], stage1_62[173], stage1_62[174]},
      {stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47], stage1_63[48]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[7],stage2_64[34],stage2_63[63],stage2_62[68]}
   );
   gpc1163_5 gpc7110 (
      {stage1_62[175], stage1_62[176], stage1_62[177]},
      {stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53], stage1_63[54]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[8],stage2_64[35],stage2_63[64],stage2_62[69]}
   );
   gpc1163_5 gpc7111 (
      {stage1_62[178], stage1_62[179], stage1_62[180]},
      {stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59], stage1_63[60]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[9],stage2_64[36],stage2_63[65],stage2_62[70]}
   );
   gpc1163_5 gpc7112 (
      {stage1_62[181], stage1_62[182], stage1_62[183]},
      {stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65], stage1_63[66]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[10],stage2_64[37],stage2_63[66],stage2_62[71]}
   );
   gpc1163_5 gpc7113 (
      {stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71], stage1_63[72]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[11],stage2_64[38],stage2_63[67],stage2_62[72]}
   );
   gpc1163_5 gpc7114 (
      {stage1_62[187], stage1_62[188], stage1_62[189]},
      {stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77], stage1_63[78]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[12],stage2_64[39],stage2_63[68],stage2_62[73]}
   );
   gpc1163_5 gpc7115 (
      {stage1_62[190], stage1_62[191], stage1_62[192]},
      {stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83], stage1_63[84]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[13],stage2_64[40],stage2_63[69],stage2_62[74]}
   );
   gpc1163_5 gpc7116 (
      {stage1_62[193], stage1_62[194], stage1_62[195]},
      {stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89], stage1_63[90]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[14],stage2_64[41],stage2_63[70],stage2_62[75]}
   );
   gpc1163_5 gpc7117 (
      {stage1_62[196], stage1_62[197], stage1_62[198]},
      {stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95], stage1_63[96]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[15],stage2_64[42],stage2_63[71],stage2_62[76]}
   );
   gpc1163_5 gpc7118 (
      {stage1_62[199], stage1_62[200], stage1_62[201]},
      {stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101], stage1_63[102]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[16],stage2_64[43],stage2_63[72],stage2_62[77]}
   );
   gpc1163_5 gpc7119 (
      {stage1_62[202], stage1_62[203], stage1_62[204]},
      {stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107], stage1_63[108]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[17],stage2_64[44],stage2_63[73],stage2_62[78]}
   );
   gpc1163_5 gpc7120 (
      {stage1_62[205], stage1_62[206], stage1_62[207]},
      {stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113], stage1_63[114]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[18],stage2_64[45],stage2_63[74],stage2_62[79]}
   );
   gpc1163_5 gpc7121 (
      {stage1_62[208], stage1_62[209], stage1_62[210]},
      {stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119], stage1_63[120]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[19],stage2_64[46],stage2_63[75],stage2_62[80]}
   );
   gpc1163_5 gpc7122 (
      {stage1_62[211], stage1_62[212], stage1_62[213]},
      {stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125], stage1_63[126]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[20],stage2_64[47],stage2_63[76],stage2_62[81]}
   );
   gpc1163_5 gpc7123 (
      {stage1_62[214], stage1_62[215], stage1_62[216]},
      {stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131], stage1_63[132]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[21],stage2_64[48],stage2_63[77],stage2_62[82]}
   );
   gpc1163_5 gpc7124 (
      {stage1_62[217], stage1_62[218], stage1_62[219]},
      {stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137], stage1_63[138]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[22],stage2_64[49],stage2_63[78],stage2_62[83]}
   );
   gpc1163_5 gpc7125 (
      {stage1_62[220], stage1_62[221], stage1_62[222]},
      {stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143], stage1_63[144]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[23],stage2_64[50],stage2_63[79],stage2_62[84]}
   );
   gpc1163_5 gpc7126 (
      {stage1_62[223], stage1_62[224], stage1_62[225]},
      {stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149], stage1_63[150]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[24],stage2_64[51],stage2_63[80],stage2_62[85]}
   );
   gpc1163_5 gpc7127 (
      {stage1_62[226], stage1_62[227], stage1_62[228]},
      {stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155], stage1_63[156]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[25],stage2_64[52],stage2_63[81],stage2_62[86]}
   );
   gpc1163_5 gpc7128 (
      {stage1_62[229], stage1_62[230], stage1_62[231]},
      {stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161], stage1_63[162]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[26],stage2_64[53],stage2_63[82],stage2_62[87]}
   );
   gpc1163_5 gpc7129 (
      {stage1_62[232], stage1_62[233], stage1_62[234]},
      {stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167], stage1_63[168]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[27],stage2_64[54],stage2_63[83],stage2_62[88]}
   );
   gpc1163_5 gpc7130 (
      {stage1_62[235], stage1_62[236], stage1_62[237]},
      {stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173], stage1_63[174]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[28],stage2_64[55],stage2_63[84],stage2_62[89]}
   );
   gpc1163_5 gpc7131 (
      {stage1_62[238], stage1_62[239], stage1_62[240]},
      {stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179], stage1_63[180]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[29],stage2_64[56],stage2_63[85],stage2_62[90]}
   );
   gpc1163_5 gpc7132 (
      {stage1_62[241], stage1_62[242], stage1_62[243]},
      {stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185], stage1_63[186]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[30],stage2_64[57],stage2_63[86],stage2_62[91]}
   );
   gpc1163_5 gpc7133 (
      {stage1_62[244], stage1_62[245], stage1_62[246]},
      {stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191], stage1_63[192]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[31],stage2_64[58],stage2_63[87],stage2_62[92]}
   );
   gpc1163_5 gpc7134 (
      {stage1_62[247], stage1_62[248], stage1_62[249]},
      {stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197], stage1_63[198]},
      {stage1_64[29]},
      {stage1_65[29]},
      {stage2_66[29],stage2_65[32],stage2_64[59],stage2_63[88],stage2_62[93]}
   );
   gpc1163_5 gpc7135 (
      {stage1_62[250], stage1_62[251], stage1_62[252]},
      {stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203], stage1_63[204]},
      {stage1_64[30]},
      {stage1_65[30]},
      {stage2_66[30],stage2_65[33],stage2_64[60],stage2_63[89],stage2_62[94]}
   );
   gpc1163_5 gpc7136 (
      {stage1_62[253], stage1_62[254], stage1_62[255]},
      {stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209], stage1_63[210]},
      {stage1_64[31]},
      {stage1_65[31]},
      {stage2_66[31],stage2_65[34],stage2_64[61],stage2_63[90],stage2_62[95]}
   );
   gpc1163_5 gpc7137 (
      {stage1_62[256], stage1_62[257], stage1_62[258]},
      {stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215], stage1_63[216]},
      {stage1_64[32]},
      {stage1_65[32]},
      {stage2_66[32],stage2_65[35],stage2_64[62],stage2_63[91],stage2_62[96]}
   );
   gpc1163_5 gpc7138 (
      {stage1_62[259], stage1_62[260], stage1_62[261]},
      {stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221], stage1_63[222]},
      {stage1_64[33]},
      {stage1_65[33]},
      {stage2_66[33],stage2_65[36],stage2_64[63],stage2_63[92],stage2_62[97]}
   );
   gpc1163_5 gpc7139 (
      {stage1_62[262], stage1_62[263], stage1_62[264]},
      {stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227], stage1_63[228]},
      {stage1_64[34]},
      {stage1_65[34]},
      {stage2_66[34],stage2_65[37],stage2_64[64],stage2_63[93],stage2_62[98]}
   );
   gpc1163_5 gpc7140 (
      {stage1_62[265], stage1_62[266], stage1_62[267]},
      {stage1_63[229], stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[35]},
      {stage1_65[35]},
      {stage2_66[35],stage2_65[38],stage2_64[65],stage2_63[94],stage2_62[99]}
   );
   gpc1163_5 gpc7141 (
      {stage1_62[268], stage1_62[269], stage1_62[270]},
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239], stage1_63[240]},
      {stage1_64[36]},
      {stage1_65[36]},
      {stage2_66[36],stage2_65[39],stage2_64[66],stage2_63[95],stage2_62[100]}
   );
   gpc1163_5 gpc7142 (
      {stage1_62[271], stage1_62[272], stage1_62[273]},
      {stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_64[37]},
      {stage1_65[37]},
      {stage2_66[37],stage2_65[40],stage2_64[67],stage2_63[96],stage2_62[101]}
   );
   gpc1163_5 gpc7143 (
      {stage1_62[274], stage1_62[275], stage1_62[276]},
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252]},
      {stage1_64[38]},
      {stage1_65[38]},
      {stage2_66[38],stage2_65[41],stage2_64[68],stage2_63[97],stage2_62[102]}
   );
   gpc1163_5 gpc7144 (
      {stage1_62[277], stage1_62[278], stage1_62[279]},
      {stage1_63[253], stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258]},
      {stage1_64[39]},
      {stage1_65[39]},
      {stage2_66[39],stage2_65[42],stage2_64[69],stage2_63[98],stage2_62[103]}
   );
   gpc1163_5 gpc7145 (
      {stage1_62[280], stage1_62[281], stage1_62[282]},
      {stage1_63[259], stage1_63[260], stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264]},
      {stage1_64[40]},
      {stage1_65[40]},
      {stage2_66[40],stage2_65[43],stage2_64[70],stage2_63[99],stage2_62[104]}
   );
   gpc1163_5 gpc7146 (
      {stage1_62[283], stage1_62[284], stage1_62[285]},
      {stage1_63[265], stage1_63[266], stage1_63[267], stage1_63[268], stage1_63[269], stage1_63[270]},
      {stage1_64[41]},
      {stage1_65[41]},
      {stage2_66[41],stage2_65[44],stage2_64[71],stage2_63[100],stage2_62[105]}
   );
   gpc1163_5 gpc7147 (
      {stage1_62[286], stage1_62[287], stage1_62[288]},
      {stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274], stage1_63[275], stage1_63[276]},
      {stage1_64[42]},
      {stage1_65[42]},
      {stage2_66[42],stage2_65[45],stage2_64[72],stage2_63[101],stage2_62[106]}
   );
   gpc1163_5 gpc7148 (
      {stage1_62[289], stage1_62[290], stage1_62[291]},
      {stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281], stage1_63[282]},
      {stage1_64[43]},
      {stage1_65[43]},
      {stage2_66[43],stage2_65[46],stage2_64[73],stage2_63[102],stage2_62[107]}
   );
   gpc1163_5 gpc7149 (
      {stage1_62[292], stage1_62[293], stage1_62[294]},
      {stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_64[44]},
      {stage1_65[44]},
      {stage2_66[44],stage2_65[47],stage2_64[74],stage2_63[103],stage2_62[108]}
   );
   gpc1163_5 gpc7150 (
      {stage1_62[295], stage1_62[296], stage1_62[297]},
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294]},
      {stage1_64[45]},
      {stage1_65[45]},
      {stage2_66[45],stage2_65[48],stage2_64[75],stage2_63[104],stage2_62[109]}
   );
   gpc606_5 gpc7151 (
      {stage1_62[298], stage1_62[299], stage1_62[300], stage1_62[301], stage1_62[302], stage1_62[303]},
      {stage1_64[46], stage1_64[47], stage1_64[48], stage1_64[49], stage1_64[50], stage1_64[51]},
      {stage2_66[46],stage2_65[49],stage2_64[76],stage2_63[105],stage2_62[110]}
   );
   gpc606_5 gpc7152 (
      {stage1_62[304], stage1_62[305], stage1_62[306], stage1_62[307], stage1_62[308], stage1_62[309]},
      {stage1_64[52], stage1_64[53], stage1_64[54], stage1_64[55], stage1_64[56], stage1_64[57]},
      {stage2_66[47],stage2_65[50],stage2_64[77],stage2_63[106],stage2_62[111]}
   );
   gpc606_5 gpc7153 (
      {stage1_62[310], stage1_62[311], stage1_62[312], stage1_62[313], stage1_62[314], stage1_62[315]},
      {stage1_64[58], stage1_64[59], stage1_64[60], stage1_64[61], stage1_64[62], stage1_64[63]},
      {stage2_66[48],stage2_65[51],stage2_64[78],stage2_63[107],stage2_62[112]}
   );
   gpc606_5 gpc7154 (
      {stage1_62[316], stage1_62[317], stage1_62[318], stage1_62[319], stage1_62[320], stage1_62[321]},
      {stage1_64[64], stage1_64[65], stage1_64[66], stage1_64[67], stage1_64[68], stage1_64[69]},
      {stage2_66[49],stage2_65[52],stage2_64[79],stage2_63[108],stage2_62[113]}
   );
   gpc606_5 gpc7155 (
      {stage1_62[322], stage1_62[323], stage1_62[324], stage1_62[325], stage1_62[326], stage1_62[327]},
      {stage1_64[70], stage1_64[71], stage1_64[72], stage1_64[73], stage1_64[74], stage1_64[75]},
      {stage2_66[50],stage2_65[53],stage2_64[80],stage2_63[109],stage2_62[114]}
   );
   gpc606_5 gpc7156 (
      {stage1_62[328], stage1_62[329], stage1_62[330], stage1_62[331], stage1_62[332], stage1_62[333]},
      {stage1_64[76], stage1_64[77], stage1_64[78], stage1_64[79], stage1_64[80], stage1_64[81]},
      {stage2_66[51],stage2_65[54],stage2_64[81],stage2_63[110],stage2_62[115]}
   );
   gpc606_5 gpc7157 (
      {stage1_62[334], stage1_62[335], stage1_62[336], stage1_62[337], stage1_62[338], stage1_62[339]},
      {stage1_64[82], stage1_64[83], stage1_64[84], stage1_64[85], stage1_64[86], stage1_64[87]},
      {stage2_66[52],stage2_65[55],stage2_64[82],stage2_63[111],stage2_62[116]}
   );
   gpc606_5 gpc7158 (
      {stage1_62[340], stage1_62[341], stage1_62[342], stage1_62[343], stage1_62[344], stage1_62[345]},
      {stage1_64[88], stage1_64[89], stage1_64[90], stage1_64[91], stage1_64[92], stage1_64[93]},
      {stage2_66[53],stage2_65[56],stage2_64[83],stage2_63[112],stage2_62[117]}
   );
   gpc1_1 gpc7159 (
      {stage1_0[112]},
      {stage2_0[27]}
   );
   gpc1_1 gpc7160 (
      {stage1_0[113]},
      {stage2_0[28]}
   );
   gpc1_1 gpc7161 (
      {stage1_0[114]},
      {stage2_0[29]}
   );
   gpc1_1 gpc7162 (
      {stage1_0[115]},
      {stage2_0[30]}
   );
   gpc1_1 gpc7163 (
      {stage1_0[116]},
      {stage2_0[31]}
   );
   gpc1_1 gpc7164 (
      {stage1_0[117]},
      {stage2_0[32]}
   );
   gpc1_1 gpc7165 (
      {stage1_0[118]},
      {stage2_0[33]}
   );
   gpc1_1 gpc7166 (
      {stage1_2[208]},
      {stage2_2[60]}
   );
   gpc1_1 gpc7167 (
      {stage1_2[209]},
      {stage2_2[61]}
   );
   gpc1_1 gpc7168 (
      {stage1_2[210]},
      {stage2_2[62]}
   );
   gpc1_1 gpc7169 (
      {stage1_2[211]},
      {stage2_2[63]}
   );
   gpc1_1 gpc7170 (
      {stage1_2[212]},
      {stage2_2[64]}
   );
   gpc1_1 gpc7171 (
      {stage1_2[213]},
      {stage2_2[65]}
   );
   gpc1_1 gpc7172 (
      {stage1_2[214]},
      {stage2_2[66]}
   );
   gpc1_1 gpc7173 (
      {stage1_2[215]},
      {stage2_2[67]}
   );
   gpc1_1 gpc7174 (
      {stage1_2[216]},
      {stage2_2[68]}
   );
   gpc1_1 gpc7175 (
      {stage1_2[217]},
      {stage2_2[69]}
   );
   gpc1_1 gpc7176 (
      {stage1_2[218]},
      {stage2_2[70]}
   );
   gpc1_1 gpc7177 (
      {stage1_2[219]},
      {stage2_2[71]}
   );
   gpc1_1 gpc7178 (
      {stage1_2[220]},
      {stage2_2[72]}
   );
   gpc1_1 gpc7179 (
      {stage1_3[139]},
      {stage2_3[71]}
   );
   gpc1_1 gpc7180 (
      {stage1_3[140]},
      {stage2_3[72]}
   );
   gpc1_1 gpc7181 (
      {stage1_3[141]},
      {stage2_3[73]}
   );
   gpc1_1 gpc7182 (
      {stage1_3[142]},
      {stage2_3[74]}
   );
   gpc1_1 gpc7183 (
      {stage1_3[143]},
      {stage2_3[75]}
   );
   gpc1_1 gpc7184 (
      {stage1_3[144]},
      {stage2_3[76]}
   );
   gpc1_1 gpc7185 (
      {stage1_3[145]},
      {stage2_3[77]}
   );
   gpc1_1 gpc7186 (
      {stage1_3[146]},
      {stage2_3[78]}
   );
   gpc1_1 gpc7187 (
      {stage1_3[147]},
      {stage2_3[79]}
   );
   gpc1_1 gpc7188 (
      {stage1_3[148]},
      {stage2_3[80]}
   );
   gpc1_1 gpc7189 (
      {stage1_3[149]},
      {stage2_3[81]}
   );
   gpc1_1 gpc7190 (
      {stage1_3[150]},
      {stage2_3[82]}
   );
   gpc1_1 gpc7191 (
      {stage1_3[151]},
      {stage2_3[83]}
   );
   gpc1_1 gpc7192 (
      {stage1_3[152]},
      {stage2_3[84]}
   );
   gpc1_1 gpc7193 (
      {stage1_3[153]},
      {stage2_3[85]}
   );
   gpc1_1 gpc7194 (
      {stage1_3[154]},
      {stage2_3[86]}
   );
   gpc1_1 gpc7195 (
      {stage1_3[155]},
      {stage2_3[87]}
   );
   gpc1_1 gpc7196 (
      {stage1_3[156]},
      {stage2_3[88]}
   );
   gpc1_1 gpc7197 (
      {stage1_3[157]},
      {stage2_3[89]}
   );
   gpc1_1 gpc7198 (
      {stage1_3[158]},
      {stage2_3[90]}
   );
   gpc1_1 gpc7199 (
      {stage1_3[159]},
      {stage2_3[91]}
   );
   gpc1_1 gpc7200 (
      {stage1_3[160]},
      {stage2_3[92]}
   );
   gpc1_1 gpc7201 (
      {stage1_3[161]},
      {stage2_3[93]}
   );
   gpc1_1 gpc7202 (
      {stage1_3[162]},
      {stage2_3[94]}
   );
   gpc1_1 gpc7203 (
      {stage1_3[163]},
      {stage2_3[95]}
   );
   gpc1_1 gpc7204 (
      {stage1_3[164]},
      {stage2_3[96]}
   );
   gpc1_1 gpc7205 (
      {stage1_3[165]},
      {stage2_3[97]}
   );
   gpc1_1 gpc7206 (
      {stage1_3[166]},
      {stage2_3[98]}
   );
   gpc1_1 gpc7207 (
      {stage1_3[167]},
      {stage2_3[99]}
   );
   gpc1_1 gpc7208 (
      {stage1_3[168]},
      {stage2_3[100]}
   );
   gpc1_1 gpc7209 (
      {stage1_3[169]},
      {stage2_3[101]}
   );
   gpc1_1 gpc7210 (
      {stage1_3[170]},
      {stage2_3[102]}
   );
   gpc1_1 gpc7211 (
      {stage1_3[171]},
      {stage2_3[103]}
   );
   gpc1_1 gpc7212 (
      {stage1_3[172]},
      {stage2_3[104]}
   );
   gpc1_1 gpc7213 (
      {stage1_3[173]},
      {stage2_3[105]}
   );
   gpc1_1 gpc7214 (
      {stage1_3[174]},
      {stage2_3[106]}
   );
   gpc1_1 gpc7215 (
      {stage1_3[175]},
      {stage2_3[107]}
   );
   gpc1_1 gpc7216 (
      {stage1_3[176]},
      {stage2_3[108]}
   );
   gpc1_1 gpc7217 (
      {stage1_3[177]},
      {stage2_3[109]}
   );
   gpc1_1 gpc7218 (
      {stage1_3[178]},
      {stage2_3[110]}
   );
   gpc1_1 gpc7219 (
      {stage1_3[179]},
      {stage2_3[111]}
   );
   gpc1_1 gpc7220 (
      {stage1_3[180]},
      {stage2_3[112]}
   );
   gpc1_1 gpc7221 (
      {stage1_3[181]},
      {stage2_3[113]}
   );
   gpc1_1 gpc7222 (
      {stage1_3[182]},
      {stage2_3[114]}
   );
   gpc1_1 gpc7223 (
      {stage1_3[183]},
      {stage2_3[115]}
   );
   gpc1_1 gpc7224 (
      {stage1_3[184]},
      {stage2_3[116]}
   );
   gpc1_1 gpc7225 (
      {stage1_3[185]},
      {stage2_3[117]}
   );
   gpc1_1 gpc7226 (
      {stage1_3[186]},
      {stage2_3[118]}
   );
   gpc1_1 gpc7227 (
      {stage1_3[187]},
      {stage2_3[119]}
   );
   gpc1_1 gpc7228 (
      {stage1_3[188]},
      {stage2_3[120]}
   );
   gpc1_1 gpc7229 (
      {stage1_3[189]},
      {stage2_3[121]}
   );
   gpc1_1 gpc7230 (
      {stage1_3[190]},
      {stage2_3[122]}
   );
   gpc1_1 gpc7231 (
      {stage1_3[191]},
      {stage2_3[123]}
   );
   gpc1_1 gpc7232 (
      {stage1_3[192]},
      {stage2_3[124]}
   );
   gpc1_1 gpc7233 (
      {stage1_3[193]},
      {stage2_3[125]}
   );
   gpc1_1 gpc7234 (
      {stage1_3[194]},
      {stage2_3[126]}
   );
   gpc1_1 gpc7235 (
      {stage1_3[195]},
      {stage2_3[127]}
   );
   gpc1_1 gpc7236 (
      {stage1_3[196]},
      {stage2_3[128]}
   );
   gpc1_1 gpc7237 (
      {stage1_3[197]},
      {stage2_3[129]}
   );
   gpc1_1 gpc7238 (
      {stage1_3[198]},
      {stage2_3[130]}
   );
   gpc1_1 gpc7239 (
      {stage1_3[199]},
      {stage2_3[131]}
   );
   gpc1_1 gpc7240 (
      {stage1_3[200]},
      {stage2_3[132]}
   );
   gpc1_1 gpc7241 (
      {stage1_3[201]},
      {stage2_3[133]}
   );
   gpc1_1 gpc7242 (
      {stage1_3[202]},
      {stage2_3[134]}
   );
   gpc1_1 gpc7243 (
      {stage1_3[203]},
      {stage2_3[135]}
   );
   gpc1_1 gpc7244 (
      {stage1_3[204]},
      {stage2_3[136]}
   );
   gpc1_1 gpc7245 (
      {stage1_3[205]},
      {stage2_3[137]}
   );
   gpc1_1 gpc7246 (
      {stage1_3[206]},
      {stage2_3[138]}
   );
   gpc1_1 gpc7247 (
      {stage1_3[207]},
      {stage2_3[139]}
   );
   gpc1_1 gpc7248 (
      {stage1_3[208]},
      {stage2_3[140]}
   );
   gpc1_1 gpc7249 (
      {stage1_3[209]},
      {stage2_3[141]}
   );
   gpc1_1 gpc7250 (
      {stage1_3[210]},
      {stage2_3[142]}
   );
   gpc1_1 gpc7251 (
      {stage1_3[211]},
      {stage2_3[143]}
   );
   gpc1_1 gpc7252 (
      {stage1_3[212]},
      {stage2_3[144]}
   );
   gpc1_1 gpc7253 (
      {stage1_3[213]},
      {stage2_3[145]}
   );
   gpc1_1 gpc7254 (
      {stage1_3[214]},
      {stage2_3[146]}
   );
   gpc1_1 gpc7255 (
      {stage1_3[215]},
      {stage2_3[147]}
   );
   gpc1_1 gpc7256 (
      {stage1_3[216]},
      {stage2_3[148]}
   );
   gpc1_1 gpc7257 (
      {stage1_3[217]},
      {stage2_3[149]}
   );
   gpc1_1 gpc7258 (
      {stage1_3[218]},
      {stage2_3[150]}
   );
   gpc1_1 gpc7259 (
      {stage1_3[219]},
      {stage2_3[151]}
   );
   gpc1_1 gpc7260 (
      {stage1_3[220]},
      {stage2_3[152]}
   );
   gpc1_1 gpc7261 (
      {stage1_3[221]},
      {stage2_3[153]}
   );
   gpc1_1 gpc7262 (
      {stage1_3[222]},
      {stage2_3[154]}
   );
   gpc1_1 gpc7263 (
      {stage1_3[223]},
      {stage2_3[155]}
   );
   gpc1_1 gpc7264 (
      {stage1_3[224]},
      {stage2_3[156]}
   );
   gpc1_1 gpc7265 (
      {stage1_3[225]},
      {stage2_3[157]}
   );
   gpc1_1 gpc7266 (
      {stage1_3[226]},
      {stage2_3[158]}
   );
   gpc1_1 gpc7267 (
      {stage1_3[227]},
      {stage2_3[159]}
   );
   gpc1_1 gpc7268 (
      {stage1_3[228]},
      {stage2_3[160]}
   );
   gpc1_1 gpc7269 (
      {stage1_3[229]},
      {stage2_3[161]}
   );
   gpc1_1 gpc7270 (
      {stage1_3[230]},
      {stage2_3[162]}
   );
   gpc1_1 gpc7271 (
      {stage1_3[231]},
      {stage2_3[163]}
   );
   gpc1_1 gpc7272 (
      {stage1_3[232]},
      {stage2_3[164]}
   );
   gpc1_1 gpc7273 (
      {stage1_3[233]},
      {stage2_3[165]}
   );
   gpc1_1 gpc7274 (
      {stage1_3[234]},
      {stage2_3[166]}
   );
   gpc1_1 gpc7275 (
      {stage1_3[235]},
      {stage2_3[167]}
   );
   gpc1_1 gpc7276 (
      {stage1_3[236]},
      {stage2_3[168]}
   );
   gpc1_1 gpc7277 (
      {stage1_3[237]},
      {stage2_3[169]}
   );
   gpc1_1 gpc7278 (
      {stage1_3[238]},
      {stage2_3[170]}
   );
   gpc1_1 gpc7279 (
      {stage1_3[239]},
      {stage2_3[171]}
   );
   gpc1_1 gpc7280 (
      {stage1_3[240]},
      {stage2_3[172]}
   );
   gpc1_1 gpc7281 (
      {stage1_3[241]},
      {stage2_3[173]}
   );
   gpc1_1 gpc7282 (
      {stage1_3[242]},
      {stage2_3[174]}
   );
   gpc1_1 gpc7283 (
      {stage1_3[243]},
      {stage2_3[175]}
   );
   gpc1_1 gpc7284 (
      {stage1_3[244]},
      {stage2_3[176]}
   );
   gpc1_1 gpc7285 (
      {stage1_3[245]},
      {stage2_3[177]}
   );
   gpc1_1 gpc7286 (
      {stage1_3[246]},
      {stage2_3[178]}
   );
   gpc1_1 gpc7287 (
      {stage1_3[247]},
      {stage2_3[179]}
   );
   gpc1_1 gpc7288 (
      {stage1_3[248]},
      {stage2_3[180]}
   );
   gpc1_1 gpc7289 (
      {stage1_3[249]},
      {stage2_3[181]}
   );
   gpc1_1 gpc7290 (
      {stage1_3[250]},
      {stage2_3[182]}
   );
   gpc1_1 gpc7291 (
      {stage1_3[251]},
      {stage2_3[183]}
   );
   gpc1_1 gpc7292 (
      {stage1_3[252]},
      {stage2_3[184]}
   );
   gpc1_1 gpc7293 (
      {stage1_3[253]},
      {stage2_3[185]}
   );
   gpc1_1 gpc7294 (
      {stage1_3[254]},
      {stage2_3[186]}
   );
   gpc1_1 gpc7295 (
      {stage1_3[255]},
      {stage2_3[187]}
   );
   gpc1_1 gpc7296 (
      {stage1_3[256]},
      {stage2_3[188]}
   );
   gpc1_1 gpc7297 (
      {stage1_3[257]},
      {stage2_3[189]}
   );
   gpc1_1 gpc7298 (
      {stage1_3[258]},
      {stage2_3[190]}
   );
   gpc1_1 gpc7299 (
      {stage1_3[259]},
      {stage2_3[191]}
   );
   gpc1_1 gpc7300 (
      {stage1_3[260]},
      {stage2_3[192]}
   );
   gpc1_1 gpc7301 (
      {stage1_3[261]},
      {stage2_3[193]}
   );
   gpc1_1 gpc7302 (
      {stage1_3[262]},
      {stage2_3[194]}
   );
   gpc1_1 gpc7303 (
      {stage1_3[263]},
      {stage2_3[195]}
   );
   gpc1_1 gpc7304 (
      {stage1_3[264]},
      {stage2_3[196]}
   );
   gpc1_1 gpc7305 (
      {stage1_3[265]},
      {stage2_3[197]}
   );
   gpc1_1 gpc7306 (
      {stage1_3[266]},
      {stage2_3[198]}
   );
   gpc1_1 gpc7307 (
      {stage1_3[267]},
      {stage2_3[199]}
   );
   gpc1_1 gpc7308 (
      {stage1_3[268]},
      {stage2_3[200]}
   );
   gpc1_1 gpc7309 (
      {stage1_3[269]},
      {stage2_3[201]}
   );
   gpc1_1 gpc7310 (
      {stage1_3[270]},
      {stage2_3[202]}
   );
   gpc1_1 gpc7311 (
      {stage1_3[271]},
      {stage2_3[203]}
   );
   gpc1_1 gpc7312 (
      {stage1_3[272]},
      {stage2_3[204]}
   );
   gpc1_1 gpc7313 (
      {stage1_3[273]},
      {stage2_3[205]}
   );
   gpc1_1 gpc7314 (
      {stage1_3[274]},
      {stage2_3[206]}
   );
   gpc1_1 gpc7315 (
      {stage1_3[275]},
      {stage2_3[207]}
   );
   gpc1_1 gpc7316 (
      {stage1_3[276]},
      {stage2_3[208]}
   );
   gpc1_1 gpc7317 (
      {stage1_3[277]},
      {stage2_3[209]}
   );
   gpc1_1 gpc7318 (
      {stage1_3[278]},
      {stage2_3[210]}
   );
   gpc1_1 gpc7319 (
      {stage1_3[279]},
      {stage2_3[211]}
   );
   gpc1_1 gpc7320 (
      {stage1_3[280]},
      {stage2_3[212]}
   );
   gpc1_1 gpc7321 (
      {stage1_3[281]},
      {stage2_3[213]}
   );
   gpc1_1 gpc7322 (
      {stage1_3[282]},
      {stage2_3[214]}
   );
   gpc1_1 gpc7323 (
      {stage1_3[283]},
      {stage2_3[215]}
   );
   gpc1_1 gpc7324 (
      {stage1_3[284]},
      {stage2_3[216]}
   );
   gpc1_1 gpc7325 (
      {stage1_3[285]},
      {stage2_3[217]}
   );
   gpc1_1 gpc7326 (
      {stage1_3[286]},
      {stage2_3[218]}
   );
   gpc1_1 gpc7327 (
      {stage1_3[287]},
      {stage2_3[219]}
   );
   gpc1_1 gpc7328 (
      {stage1_3[288]},
      {stage2_3[220]}
   );
   gpc1_1 gpc7329 (
      {stage1_3[289]},
      {stage2_3[221]}
   );
   gpc1_1 gpc7330 (
      {stage1_3[290]},
      {stage2_3[222]}
   );
   gpc1_1 gpc7331 (
      {stage1_3[291]},
      {stage2_3[223]}
   );
   gpc1_1 gpc7332 (
      {stage1_3[292]},
      {stage2_3[224]}
   );
   gpc1_1 gpc7333 (
      {stage1_3[293]},
      {stage2_3[225]}
   );
   gpc1_1 gpc7334 (
      {stage1_3[294]},
      {stage2_3[226]}
   );
   gpc1_1 gpc7335 (
      {stage1_3[295]},
      {stage2_3[227]}
   );
   gpc1_1 gpc7336 (
      {stage1_3[296]},
      {stage2_3[228]}
   );
   gpc1_1 gpc7337 (
      {stage1_3[297]},
      {stage2_3[229]}
   );
   gpc1_1 gpc7338 (
      {stage1_3[298]},
      {stage2_3[230]}
   );
   gpc1_1 gpc7339 (
      {stage1_3[299]},
      {stage2_3[231]}
   );
   gpc1_1 gpc7340 (
      {stage1_3[300]},
      {stage2_3[232]}
   );
   gpc1_1 gpc7341 (
      {stage1_3[301]},
      {stage2_3[233]}
   );
   gpc1_1 gpc7342 (
      {stage1_3[302]},
      {stage2_3[234]}
   );
   gpc1_1 gpc7343 (
      {stage1_3[303]},
      {stage2_3[235]}
   );
   gpc1_1 gpc7344 (
      {stage1_3[304]},
      {stage2_3[236]}
   );
   gpc1_1 gpc7345 (
      {stage1_3[305]},
      {stage2_3[237]}
   );
   gpc1_1 gpc7346 (
      {stage1_3[306]},
      {stage2_3[238]}
   );
   gpc1_1 gpc7347 (
      {stage1_3[307]},
      {stage2_3[239]}
   );
   gpc1_1 gpc7348 (
      {stage1_3[308]},
      {stage2_3[240]}
   );
   gpc1_1 gpc7349 (
      {stage1_3[309]},
      {stage2_3[241]}
   );
   gpc1_1 gpc7350 (
      {stage1_3[310]},
      {stage2_3[242]}
   );
   gpc1_1 gpc7351 (
      {stage1_3[311]},
      {stage2_3[243]}
   );
   gpc1_1 gpc7352 (
      {stage1_3[312]},
      {stage2_3[244]}
   );
   gpc1_1 gpc7353 (
      {stage1_3[313]},
      {stage2_3[245]}
   );
   gpc1_1 gpc7354 (
      {stage1_3[314]},
      {stage2_3[246]}
   );
   gpc1_1 gpc7355 (
      {stage1_3[315]},
      {stage2_3[247]}
   );
   gpc1_1 gpc7356 (
      {stage1_3[316]},
      {stage2_3[248]}
   );
   gpc1_1 gpc7357 (
      {stage1_3[317]},
      {stage2_3[249]}
   );
   gpc1_1 gpc7358 (
      {stage1_3[318]},
      {stage2_3[250]}
   );
   gpc1_1 gpc7359 (
      {stage1_3[319]},
      {stage2_3[251]}
   );
   gpc1_1 gpc7360 (
      {stage1_3[320]},
      {stage2_3[252]}
   );
   gpc1_1 gpc7361 (
      {stage1_3[321]},
      {stage2_3[253]}
   );
   gpc1_1 gpc7362 (
      {stage1_4[247]},
      {stage2_4[89]}
   );
   gpc1_1 gpc7363 (
      {stage1_4[248]},
      {stage2_4[90]}
   );
   gpc1_1 gpc7364 (
      {stage1_4[249]},
      {stage2_4[91]}
   );
   gpc1_1 gpc7365 (
      {stage1_4[250]},
      {stage2_4[92]}
   );
   gpc1_1 gpc7366 (
      {stage1_5[188]},
      {stage2_5[83]}
   );
   gpc1_1 gpc7367 (
      {stage1_5[189]},
      {stage2_5[84]}
   );
   gpc1_1 gpc7368 (
      {stage1_5[190]},
      {stage2_5[85]}
   );
   gpc1_1 gpc7369 (
      {stage1_5[191]},
      {stage2_5[86]}
   );
   gpc1_1 gpc7370 (
      {stage1_5[192]},
      {stage2_5[87]}
   );
   gpc1_1 gpc7371 (
      {stage1_5[193]},
      {stage2_5[88]}
   );
   gpc1_1 gpc7372 (
      {stage1_5[194]},
      {stage2_5[89]}
   );
   gpc1_1 gpc7373 (
      {stage1_5[195]},
      {stage2_5[90]}
   );
   gpc1_1 gpc7374 (
      {stage1_5[196]},
      {stage2_5[91]}
   );
   gpc1_1 gpc7375 (
      {stage1_5[197]},
      {stage2_5[92]}
   );
   gpc1_1 gpc7376 (
      {stage1_5[198]},
      {stage2_5[93]}
   );
   gpc1_1 gpc7377 (
      {stage1_5[199]},
      {stage2_5[94]}
   );
   gpc1_1 gpc7378 (
      {stage1_5[200]},
      {stage2_5[95]}
   );
   gpc1_1 gpc7379 (
      {stage1_5[201]},
      {stage2_5[96]}
   );
   gpc1_1 gpc7380 (
      {stage1_5[202]},
      {stage2_5[97]}
   );
   gpc1_1 gpc7381 (
      {stage1_5[203]},
      {stage2_5[98]}
   );
   gpc1_1 gpc7382 (
      {stage1_5[204]},
      {stage2_5[99]}
   );
   gpc1_1 gpc7383 (
      {stage1_5[205]},
      {stage2_5[100]}
   );
   gpc1_1 gpc7384 (
      {stage1_5[206]},
      {stage2_5[101]}
   );
   gpc1_1 gpc7385 (
      {stage1_5[207]},
      {stage2_5[102]}
   );
   gpc1_1 gpc7386 (
      {stage1_5[208]},
      {stage2_5[103]}
   );
   gpc1_1 gpc7387 (
      {stage1_5[209]},
      {stage2_5[104]}
   );
   gpc1_1 gpc7388 (
      {stage1_5[210]},
      {stage2_5[105]}
   );
   gpc1_1 gpc7389 (
      {stage1_5[211]},
      {stage2_5[106]}
   );
   gpc1_1 gpc7390 (
      {stage1_5[212]},
      {stage2_5[107]}
   );
   gpc1_1 gpc7391 (
      {stage1_5[213]},
      {stage2_5[108]}
   );
   gpc1_1 gpc7392 (
      {stage1_5[214]},
      {stage2_5[109]}
   );
   gpc1_1 gpc7393 (
      {stage1_5[215]},
      {stage2_5[110]}
   );
   gpc1_1 gpc7394 (
      {stage1_5[216]},
      {stage2_5[111]}
   );
   gpc1_1 gpc7395 (
      {stage1_6[135]},
      {stage2_6[76]}
   );
   gpc1_1 gpc7396 (
      {stage1_6[136]},
      {stage2_6[77]}
   );
   gpc1_1 gpc7397 (
      {stage1_6[137]},
      {stage2_6[78]}
   );
   gpc1_1 gpc7398 (
      {stage1_6[138]},
      {stage2_6[79]}
   );
   gpc1_1 gpc7399 (
      {stage1_6[139]},
      {stage2_6[80]}
   );
   gpc1_1 gpc7400 (
      {stage1_6[140]},
      {stage2_6[81]}
   );
   gpc1_1 gpc7401 (
      {stage1_6[141]},
      {stage2_6[82]}
   );
   gpc1_1 gpc7402 (
      {stage1_6[142]},
      {stage2_6[83]}
   );
   gpc1_1 gpc7403 (
      {stage1_6[143]},
      {stage2_6[84]}
   );
   gpc1_1 gpc7404 (
      {stage1_6[144]},
      {stage2_6[85]}
   );
   gpc1_1 gpc7405 (
      {stage1_6[145]},
      {stage2_6[86]}
   );
   gpc1_1 gpc7406 (
      {stage1_6[146]},
      {stage2_6[87]}
   );
   gpc1_1 gpc7407 (
      {stage1_6[147]},
      {stage2_6[88]}
   );
   gpc1_1 gpc7408 (
      {stage1_6[148]},
      {stage2_6[89]}
   );
   gpc1_1 gpc7409 (
      {stage1_6[149]},
      {stage2_6[90]}
   );
   gpc1_1 gpc7410 (
      {stage1_6[150]},
      {stage2_6[91]}
   );
   gpc1_1 gpc7411 (
      {stage1_6[151]},
      {stage2_6[92]}
   );
   gpc1_1 gpc7412 (
      {stage1_6[152]},
      {stage2_6[93]}
   );
   gpc1_1 gpc7413 (
      {stage1_6[153]},
      {stage2_6[94]}
   );
   gpc1_1 gpc7414 (
      {stage1_6[154]},
      {stage2_6[95]}
   );
   gpc1_1 gpc7415 (
      {stage1_6[155]},
      {stage2_6[96]}
   );
   gpc1_1 gpc7416 (
      {stage1_6[156]},
      {stage2_6[97]}
   );
   gpc1_1 gpc7417 (
      {stage1_6[157]},
      {stage2_6[98]}
   );
   gpc1_1 gpc7418 (
      {stage1_6[158]},
      {stage2_6[99]}
   );
   gpc1_1 gpc7419 (
      {stage1_6[159]},
      {stage2_6[100]}
   );
   gpc1_1 gpc7420 (
      {stage1_6[160]},
      {stage2_6[101]}
   );
   gpc1_1 gpc7421 (
      {stage1_6[161]},
      {stage2_6[102]}
   );
   gpc1_1 gpc7422 (
      {stage1_6[162]},
      {stage2_6[103]}
   );
   gpc1_1 gpc7423 (
      {stage1_6[163]},
      {stage2_6[104]}
   );
   gpc1_1 gpc7424 (
      {stage1_6[164]},
      {stage2_6[105]}
   );
   gpc1_1 gpc7425 (
      {stage1_6[165]},
      {stage2_6[106]}
   );
   gpc1_1 gpc7426 (
      {stage1_6[166]},
      {stage2_6[107]}
   );
   gpc1_1 gpc7427 (
      {stage1_6[167]},
      {stage2_6[108]}
   );
   gpc1_1 gpc7428 (
      {stage1_6[168]},
      {stage2_6[109]}
   );
   gpc1_1 gpc7429 (
      {stage1_6[169]},
      {stage2_6[110]}
   );
   gpc1_1 gpc7430 (
      {stage1_6[170]},
      {stage2_6[111]}
   );
   gpc1_1 gpc7431 (
      {stage1_6[171]},
      {stage2_6[112]}
   );
   gpc1_1 gpc7432 (
      {stage1_6[172]},
      {stage2_6[113]}
   );
   gpc1_1 gpc7433 (
      {stage1_6[173]},
      {stage2_6[114]}
   );
   gpc1_1 gpc7434 (
      {stage1_6[174]},
      {stage2_6[115]}
   );
   gpc1_1 gpc7435 (
      {stage1_6[175]},
      {stage2_6[116]}
   );
   gpc1_1 gpc7436 (
      {stage1_6[176]},
      {stage2_6[117]}
   );
   gpc1_1 gpc7437 (
      {stage1_6[177]},
      {stage2_6[118]}
   );
   gpc1_1 gpc7438 (
      {stage1_6[178]},
      {stage2_6[119]}
   );
   gpc1_1 gpc7439 (
      {stage1_6[179]},
      {stage2_6[120]}
   );
   gpc1_1 gpc7440 (
      {stage1_8[168]},
      {stage2_8[102]}
   );
   gpc1_1 gpc7441 (
      {stage1_8[169]},
      {stage2_8[103]}
   );
   gpc1_1 gpc7442 (
      {stage1_8[170]},
      {stage2_8[104]}
   );
   gpc1_1 gpc7443 (
      {stage1_8[171]},
      {stage2_8[105]}
   );
   gpc1_1 gpc7444 (
      {stage1_8[172]},
      {stage2_8[106]}
   );
   gpc1_1 gpc7445 (
      {stage1_8[173]},
      {stage2_8[107]}
   );
   gpc1_1 gpc7446 (
      {stage1_8[174]},
      {stage2_8[108]}
   );
   gpc1_1 gpc7447 (
      {stage1_8[175]},
      {stage2_8[109]}
   );
   gpc1_1 gpc7448 (
      {stage1_8[176]},
      {stage2_8[110]}
   );
   gpc1_1 gpc7449 (
      {stage1_8[177]},
      {stage2_8[111]}
   );
   gpc1_1 gpc7450 (
      {stage1_8[178]},
      {stage2_8[112]}
   );
   gpc1_1 gpc7451 (
      {stage1_8[179]},
      {stage2_8[113]}
   );
   gpc1_1 gpc7452 (
      {stage1_8[180]},
      {stage2_8[114]}
   );
   gpc1_1 gpc7453 (
      {stage1_8[181]},
      {stage2_8[115]}
   );
   gpc1_1 gpc7454 (
      {stage1_8[182]},
      {stage2_8[116]}
   );
   gpc1_1 gpc7455 (
      {stage1_8[183]},
      {stage2_8[117]}
   );
   gpc1_1 gpc7456 (
      {stage1_8[184]},
      {stage2_8[118]}
   );
   gpc1_1 gpc7457 (
      {stage1_8[185]},
      {stage2_8[119]}
   );
   gpc1_1 gpc7458 (
      {stage1_8[186]},
      {stage2_8[120]}
   );
   gpc1_1 gpc7459 (
      {stage1_8[187]},
      {stage2_8[121]}
   );
   gpc1_1 gpc7460 (
      {stage1_8[188]},
      {stage2_8[122]}
   );
   gpc1_1 gpc7461 (
      {stage1_8[189]},
      {stage2_8[123]}
   );
   gpc1_1 gpc7462 (
      {stage1_8[190]},
      {stage2_8[124]}
   );
   gpc1_1 gpc7463 (
      {stage1_8[191]},
      {stage2_8[125]}
   );
   gpc1_1 gpc7464 (
      {stage1_8[192]},
      {stage2_8[126]}
   );
   gpc1_1 gpc7465 (
      {stage1_8[193]},
      {stage2_8[127]}
   );
   gpc1_1 gpc7466 (
      {stage1_8[194]},
      {stage2_8[128]}
   );
   gpc1_1 gpc7467 (
      {stage1_8[195]},
      {stage2_8[129]}
   );
   gpc1_1 gpc7468 (
      {stage1_8[196]},
      {stage2_8[130]}
   );
   gpc1_1 gpc7469 (
      {stage1_8[197]},
      {stage2_8[131]}
   );
   gpc1_1 gpc7470 (
      {stage1_8[198]},
      {stage2_8[132]}
   );
   gpc1_1 gpc7471 (
      {stage1_8[199]},
      {stage2_8[133]}
   );
   gpc1_1 gpc7472 (
      {stage1_8[200]},
      {stage2_8[134]}
   );
   gpc1_1 gpc7473 (
      {stage1_8[201]},
      {stage2_8[135]}
   );
   gpc1_1 gpc7474 (
      {stage1_8[202]},
      {stage2_8[136]}
   );
   gpc1_1 gpc7475 (
      {stage1_8[203]},
      {stage2_8[137]}
   );
   gpc1_1 gpc7476 (
      {stage1_8[204]},
      {stage2_8[138]}
   );
   gpc1_1 gpc7477 (
      {stage1_8[205]},
      {stage2_8[139]}
   );
   gpc1_1 gpc7478 (
      {stage1_8[206]},
      {stage2_8[140]}
   );
   gpc1_1 gpc7479 (
      {stage1_8[207]},
      {stage2_8[141]}
   );
   gpc1_1 gpc7480 (
      {stage1_8[208]},
      {stage2_8[142]}
   );
   gpc1_1 gpc7481 (
      {stage1_8[209]},
      {stage2_8[143]}
   );
   gpc1_1 gpc7482 (
      {stage1_8[210]},
      {stage2_8[144]}
   );
   gpc1_1 gpc7483 (
      {stage1_8[211]},
      {stage2_8[145]}
   );
   gpc1_1 gpc7484 (
      {stage1_8[212]},
      {stage2_8[146]}
   );
   gpc1_1 gpc7485 (
      {stage1_8[213]},
      {stage2_8[147]}
   );
   gpc1_1 gpc7486 (
      {stage1_8[214]},
      {stage2_8[148]}
   );
   gpc1_1 gpc7487 (
      {stage1_8[215]},
      {stage2_8[149]}
   );
   gpc1_1 gpc7488 (
      {stage1_8[216]},
      {stage2_8[150]}
   );
   gpc1_1 gpc7489 (
      {stage1_8[217]},
      {stage2_8[151]}
   );
   gpc1_1 gpc7490 (
      {stage1_8[218]},
      {stage2_8[152]}
   );
   gpc1_1 gpc7491 (
      {stage1_8[219]},
      {stage2_8[153]}
   );
   gpc1_1 gpc7492 (
      {stage1_8[220]},
      {stage2_8[154]}
   );
   gpc1_1 gpc7493 (
      {stage1_8[221]},
      {stage2_8[155]}
   );
   gpc1_1 gpc7494 (
      {stage1_8[222]},
      {stage2_8[156]}
   );
   gpc1_1 gpc7495 (
      {stage1_8[223]},
      {stage2_8[157]}
   );
   gpc1_1 gpc7496 (
      {stage1_8[224]},
      {stage2_8[158]}
   );
   gpc1_1 gpc7497 (
      {stage1_8[225]},
      {stage2_8[159]}
   );
   gpc1_1 gpc7498 (
      {stage1_8[226]},
      {stage2_8[160]}
   );
   gpc1_1 gpc7499 (
      {stage1_8[227]},
      {stage2_8[161]}
   );
   gpc1_1 gpc7500 (
      {stage1_8[228]},
      {stage2_8[162]}
   );
   gpc1_1 gpc7501 (
      {stage1_8[229]},
      {stage2_8[163]}
   );
   gpc1_1 gpc7502 (
      {stage1_8[230]},
      {stage2_8[164]}
   );
   gpc1_1 gpc7503 (
      {stage1_8[231]},
      {stage2_8[165]}
   );
   gpc1_1 gpc7504 (
      {stage1_8[232]},
      {stage2_8[166]}
   );
   gpc1_1 gpc7505 (
      {stage1_8[233]},
      {stage2_8[167]}
   );
   gpc1_1 gpc7506 (
      {stage1_8[234]},
      {stage2_8[168]}
   );
   gpc1_1 gpc7507 (
      {stage1_8[235]},
      {stage2_8[169]}
   );
   gpc1_1 gpc7508 (
      {stage1_8[236]},
      {stage2_8[170]}
   );
   gpc1_1 gpc7509 (
      {stage1_8[237]},
      {stage2_8[171]}
   );
   gpc1_1 gpc7510 (
      {stage1_8[238]},
      {stage2_8[172]}
   );
   gpc1_1 gpc7511 (
      {stage1_9[360]},
      {stage2_9[102]}
   );
   gpc1_1 gpc7512 (
      {stage1_9[361]},
      {stage2_9[103]}
   );
   gpc1_1 gpc7513 (
      {stage1_9[362]},
      {stage2_9[104]}
   );
   gpc1_1 gpc7514 (
      {stage1_10[101]},
      {stage2_10[82]}
   );
   gpc1_1 gpc7515 (
      {stage1_10[102]},
      {stage2_10[83]}
   );
   gpc1_1 gpc7516 (
      {stage1_10[103]},
      {stage2_10[84]}
   );
   gpc1_1 gpc7517 (
      {stage1_10[104]},
      {stage2_10[85]}
   );
   gpc1_1 gpc7518 (
      {stage1_10[105]},
      {stage2_10[86]}
   );
   gpc1_1 gpc7519 (
      {stage1_10[106]},
      {stage2_10[87]}
   );
   gpc1_1 gpc7520 (
      {stage1_10[107]},
      {stage2_10[88]}
   );
   gpc1_1 gpc7521 (
      {stage1_10[108]},
      {stage2_10[89]}
   );
   gpc1_1 gpc7522 (
      {stage1_10[109]},
      {stage2_10[90]}
   );
   gpc1_1 gpc7523 (
      {stage1_10[110]},
      {stage2_10[91]}
   );
   gpc1_1 gpc7524 (
      {stage1_10[111]},
      {stage2_10[92]}
   );
   gpc1_1 gpc7525 (
      {stage1_10[112]},
      {stage2_10[93]}
   );
   gpc1_1 gpc7526 (
      {stage1_10[113]},
      {stage2_10[94]}
   );
   gpc1_1 gpc7527 (
      {stage1_10[114]},
      {stage2_10[95]}
   );
   gpc1_1 gpc7528 (
      {stage1_10[115]},
      {stage2_10[96]}
   );
   gpc1_1 gpc7529 (
      {stage1_10[116]},
      {stage2_10[97]}
   );
   gpc1_1 gpc7530 (
      {stage1_10[117]},
      {stage2_10[98]}
   );
   gpc1_1 gpc7531 (
      {stage1_10[118]},
      {stage2_10[99]}
   );
   gpc1_1 gpc7532 (
      {stage1_10[119]},
      {stage2_10[100]}
   );
   gpc1_1 gpc7533 (
      {stage1_10[120]},
      {stage2_10[101]}
   );
   gpc1_1 gpc7534 (
      {stage1_10[121]},
      {stage2_10[102]}
   );
   gpc1_1 gpc7535 (
      {stage1_10[122]},
      {stage2_10[103]}
   );
   gpc1_1 gpc7536 (
      {stage1_10[123]},
      {stage2_10[104]}
   );
   gpc1_1 gpc7537 (
      {stage1_10[124]},
      {stage2_10[105]}
   );
   gpc1_1 gpc7538 (
      {stage1_10[125]},
      {stage2_10[106]}
   );
   gpc1_1 gpc7539 (
      {stage1_10[126]},
      {stage2_10[107]}
   );
   gpc1_1 gpc7540 (
      {stage1_10[127]},
      {stage2_10[108]}
   );
   gpc1_1 gpc7541 (
      {stage1_10[128]},
      {stage2_10[109]}
   );
   gpc1_1 gpc7542 (
      {stage1_10[129]},
      {stage2_10[110]}
   );
   gpc1_1 gpc7543 (
      {stage1_10[130]},
      {stage2_10[111]}
   );
   gpc1_1 gpc7544 (
      {stage1_10[131]},
      {stage2_10[112]}
   );
   gpc1_1 gpc7545 (
      {stage1_10[132]},
      {stage2_10[113]}
   );
   gpc1_1 gpc7546 (
      {stage1_10[133]},
      {stage2_10[114]}
   );
   gpc1_1 gpc7547 (
      {stage1_10[134]},
      {stage2_10[115]}
   );
   gpc1_1 gpc7548 (
      {stage1_10[135]},
      {stage2_10[116]}
   );
   gpc1_1 gpc7549 (
      {stage1_10[136]},
      {stage2_10[117]}
   );
   gpc1_1 gpc7550 (
      {stage1_10[137]},
      {stage2_10[118]}
   );
   gpc1_1 gpc7551 (
      {stage1_10[138]},
      {stage2_10[119]}
   );
   gpc1_1 gpc7552 (
      {stage1_10[139]},
      {stage2_10[120]}
   );
   gpc1_1 gpc7553 (
      {stage1_10[140]},
      {stage2_10[121]}
   );
   gpc1_1 gpc7554 (
      {stage1_10[141]},
      {stage2_10[122]}
   );
   gpc1_1 gpc7555 (
      {stage1_10[142]},
      {stage2_10[123]}
   );
   gpc1_1 gpc7556 (
      {stage1_10[143]},
      {stage2_10[124]}
   );
   gpc1_1 gpc7557 (
      {stage1_10[144]},
      {stage2_10[125]}
   );
   gpc1_1 gpc7558 (
      {stage1_10[145]},
      {stage2_10[126]}
   );
   gpc1_1 gpc7559 (
      {stage1_10[146]},
      {stage2_10[127]}
   );
   gpc1_1 gpc7560 (
      {stage1_10[147]},
      {stage2_10[128]}
   );
   gpc1_1 gpc7561 (
      {stage1_10[148]},
      {stage2_10[129]}
   );
   gpc1_1 gpc7562 (
      {stage1_10[149]},
      {stage2_10[130]}
   );
   gpc1_1 gpc7563 (
      {stage1_10[150]},
      {stage2_10[131]}
   );
   gpc1_1 gpc7564 (
      {stage1_10[151]},
      {stage2_10[132]}
   );
   gpc1_1 gpc7565 (
      {stage1_10[152]},
      {stage2_10[133]}
   );
   gpc1_1 gpc7566 (
      {stage1_11[307]},
      {stage2_11[125]}
   );
   gpc1_1 gpc7567 (
      {stage1_11[308]},
      {stage2_11[126]}
   );
   gpc1_1 gpc7568 (
      {stage1_11[309]},
      {stage2_11[127]}
   );
   gpc1_1 gpc7569 (
      {stage1_11[310]},
      {stage2_11[128]}
   );
   gpc1_1 gpc7570 (
      {stage1_11[311]},
      {stage2_11[129]}
   );
   gpc1_1 gpc7571 (
      {stage1_11[312]},
      {stage2_11[130]}
   );
   gpc1_1 gpc7572 (
      {stage1_11[313]},
      {stage2_11[131]}
   );
   gpc1_1 gpc7573 (
      {stage1_11[314]},
      {stage2_11[132]}
   );
   gpc1_1 gpc7574 (
      {stage1_11[315]},
      {stage2_11[133]}
   );
   gpc1_1 gpc7575 (
      {stage1_11[316]},
      {stage2_11[134]}
   );
   gpc1_1 gpc7576 (
      {stage1_11[317]},
      {stage2_11[135]}
   );
   gpc1_1 gpc7577 (
      {stage1_12[177]},
      {stage2_12[86]}
   );
   gpc1_1 gpc7578 (
      {stage1_12[178]},
      {stage2_12[87]}
   );
   gpc1_1 gpc7579 (
      {stage1_12[179]},
      {stage2_12[88]}
   );
   gpc1_1 gpc7580 (
      {stage1_12[180]},
      {stage2_12[89]}
   );
   gpc1_1 gpc7581 (
      {stage1_12[181]},
      {stage2_12[90]}
   );
   gpc1_1 gpc7582 (
      {stage1_12[182]},
      {stage2_12[91]}
   );
   gpc1_1 gpc7583 (
      {stage1_12[183]},
      {stage2_12[92]}
   );
   gpc1_1 gpc7584 (
      {stage1_12[184]},
      {stage2_12[93]}
   );
   gpc1_1 gpc7585 (
      {stage1_12[185]},
      {stage2_12[94]}
   );
   gpc1_1 gpc7586 (
      {stage1_12[186]},
      {stage2_12[95]}
   );
   gpc1_1 gpc7587 (
      {stage1_12[187]},
      {stage2_12[96]}
   );
   gpc1_1 gpc7588 (
      {stage1_12[188]},
      {stage2_12[97]}
   );
   gpc1_1 gpc7589 (
      {stage1_12[189]},
      {stage2_12[98]}
   );
   gpc1_1 gpc7590 (
      {stage1_12[190]},
      {stage2_12[99]}
   );
   gpc1_1 gpc7591 (
      {stage1_12[191]},
      {stage2_12[100]}
   );
   gpc1_1 gpc7592 (
      {stage1_12[192]},
      {stage2_12[101]}
   );
   gpc1_1 gpc7593 (
      {stage1_12[193]},
      {stage2_12[102]}
   );
   gpc1_1 gpc7594 (
      {stage1_12[194]},
      {stage2_12[103]}
   );
   gpc1_1 gpc7595 (
      {stage1_12[195]},
      {stage2_12[104]}
   );
   gpc1_1 gpc7596 (
      {stage1_12[196]},
      {stage2_12[105]}
   );
   gpc1_1 gpc7597 (
      {stage1_12[197]},
      {stage2_12[106]}
   );
   gpc1_1 gpc7598 (
      {stage1_12[198]},
      {stage2_12[107]}
   );
   gpc1_1 gpc7599 (
      {stage1_12[199]},
      {stage2_12[108]}
   );
   gpc1_1 gpc7600 (
      {stage1_12[200]},
      {stage2_12[109]}
   );
   gpc1_1 gpc7601 (
      {stage1_12[201]},
      {stage2_12[110]}
   );
   gpc1_1 gpc7602 (
      {stage1_12[202]},
      {stage2_12[111]}
   );
   gpc1_1 gpc7603 (
      {stage1_12[203]},
      {stage2_12[112]}
   );
   gpc1_1 gpc7604 (
      {stage1_12[204]},
      {stage2_12[113]}
   );
   gpc1_1 gpc7605 (
      {stage1_12[205]},
      {stage2_12[114]}
   );
   gpc1_1 gpc7606 (
      {stage1_12[206]},
      {stage2_12[115]}
   );
   gpc1_1 gpc7607 (
      {stage1_12[207]},
      {stage2_12[116]}
   );
   gpc1_1 gpc7608 (
      {stage1_12[208]},
      {stage2_12[117]}
   );
   gpc1_1 gpc7609 (
      {stage1_12[209]},
      {stage2_12[118]}
   );
   gpc1_1 gpc7610 (
      {stage1_12[210]},
      {stage2_12[119]}
   );
   gpc1_1 gpc7611 (
      {stage1_12[211]},
      {stage2_12[120]}
   );
   gpc1_1 gpc7612 (
      {stage1_12[212]},
      {stage2_12[121]}
   );
   gpc1_1 gpc7613 (
      {stage1_12[213]},
      {stage2_12[122]}
   );
   gpc1_1 gpc7614 (
      {stage1_12[214]},
      {stage2_12[123]}
   );
   gpc1_1 gpc7615 (
      {stage1_12[215]},
      {stage2_12[124]}
   );
   gpc1_1 gpc7616 (
      {stage1_12[216]},
      {stage2_12[125]}
   );
   gpc1_1 gpc7617 (
      {stage1_12[217]},
      {stage2_12[126]}
   );
   gpc1_1 gpc7618 (
      {stage1_12[218]},
      {stage2_12[127]}
   );
   gpc1_1 gpc7619 (
      {stage1_13[183]},
      {stage2_13[70]}
   );
   gpc1_1 gpc7620 (
      {stage1_13[184]},
      {stage2_13[71]}
   );
   gpc1_1 gpc7621 (
      {stage1_14[246]},
      {stage2_14[105]}
   );
   gpc1_1 gpc7622 (
      {stage1_14[247]},
      {stage2_14[106]}
   );
   gpc1_1 gpc7623 (
      {stage1_14[248]},
      {stage2_14[107]}
   );
   gpc1_1 gpc7624 (
      {stage1_14[249]},
      {stage2_14[108]}
   );
   gpc1_1 gpc7625 (
      {stage1_14[250]},
      {stage2_14[109]}
   );
   gpc1_1 gpc7626 (
      {stage1_14[251]},
      {stage2_14[110]}
   );
   gpc1_1 gpc7627 (
      {stage1_14[252]},
      {stage2_14[111]}
   );
   gpc1_1 gpc7628 (
      {stage1_14[253]},
      {stage2_14[112]}
   );
   gpc1_1 gpc7629 (
      {stage1_14[254]},
      {stage2_14[113]}
   );
   gpc1_1 gpc7630 (
      {stage1_14[255]},
      {stage2_14[114]}
   );
   gpc1_1 gpc7631 (
      {stage1_15[255]},
      {stage2_15[112]}
   );
   gpc1_1 gpc7632 (
      {stage1_15[256]},
      {stage2_15[113]}
   );
   gpc1_1 gpc7633 (
      {stage1_15[257]},
      {stage2_15[114]}
   );
   gpc1_1 gpc7634 (
      {stage1_16[182]},
      {stage2_16[68]}
   );
   gpc1_1 gpc7635 (
      {stage1_16[183]},
      {stage2_16[69]}
   );
   gpc1_1 gpc7636 (
      {stage1_16[184]},
      {stage2_16[70]}
   );
   gpc1_1 gpc7637 (
      {stage1_16[185]},
      {stage2_16[71]}
   );
   gpc1_1 gpc7638 (
      {stage1_16[186]},
      {stage2_16[72]}
   );
   gpc1_1 gpc7639 (
      {stage1_16[187]},
      {stage2_16[73]}
   );
   gpc1_1 gpc7640 (
      {stage1_16[188]},
      {stage2_16[74]}
   );
   gpc1_1 gpc7641 (
      {stage1_16[189]},
      {stage2_16[75]}
   );
   gpc1_1 gpc7642 (
      {stage1_16[190]},
      {stage2_16[76]}
   );
   gpc1_1 gpc7643 (
      {stage1_16[191]},
      {stage2_16[77]}
   );
   gpc1_1 gpc7644 (
      {stage1_16[192]},
      {stage2_16[78]}
   );
   gpc1_1 gpc7645 (
      {stage1_16[193]},
      {stage2_16[79]}
   );
   gpc1_1 gpc7646 (
      {stage1_16[194]},
      {stage2_16[80]}
   );
   gpc1_1 gpc7647 (
      {stage1_16[195]},
      {stage2_16[81]}
   );
   gpc1_1 gpc7648 (
      {stage1_16[196]},
      {stage2_16[82]}
   );
   gpc1_1 gpc7649 (
      {stage1_16[197]},
      {stage2_16[83]}
   );
   gpc1_1 gpc7650 (
      {stage1_16[198]},
      {stage2_16[84]}
   );
   gpc1_1 gpc7651 (
      {stage1_16[199]},
      {stage2_16[85]}
   );
   gpc1_1 gpc7652 (
      {stage1_16[200]},
      {stage2_16[86]}
   );
   gpc1_1 gpc7653 (
      {stage1_16[201]},
      {stage2_16[87]}
   );
   gpc1_1 gpc7654 (
      {stage1_16[202]},
      {stage2_16[88]}
   );
   gpc1_1 gpc7655 (
      {stage1_16[203]},
      {stage2_16[89]}
   );
   gpc1_1 gpc7656 (
      {stage1_16[204]},
      {stage2_16[90]}
   );
   gpc1_1 gpc7657 (
      {stage1_16[205]},
      {stage2_16[91]}
   );
   gpc1_1 gpc7658 (
      {stage1_16[206]},
      {stage2_16[92]}
   );
   gpc1_1 gpc7659 (
      {stage1_16[207]},
      {stage2_16[93]}
   );
   gpc1_1 gpc7660 (
      {stage1_16[208]},
      {stage2_16[94]}
   );
   gpc1_1 gpc7661 (
      {stage1_16[209]},
      {stage2_16[95]}
   );
   gpc1_1 gpc7662 (
      {stage1_16[210]},
      {stage2_16[96]}
   );
   gpc1_1 gpc7663 (
      {stage1_16[211]},
      {stage2_16[97]}
   );
   gpc1_1 gpc7664 (
      {stage1_16[212]},
      {stage2_16[98]}
   );
   gpc1_1 gpc7665 (
      {stage1_16[213]},
      {stage2_16[99]}
   );
   gpc1_1 gpc7666 (
      {stage1_16[214]},
      {stage2_16[100]}
   );
   gpc1_1 gpc7667 (
      {stage1_16[215]},
      {stage2_16[101]}
   );
   gpc1_1 gpc7668 (
      {stage1_16[216]},
      {stage2_16[102]}
   );
   gpc1_1 gpc7669 (
      {stage1_16[217]},
      {stage2_16[103]}
   );
   gpc1_1 gpc7670 (
      {stage1_16[218]},
      {stage2_16[104]}
   );
   gpc1_1 gpc7671 (
      {stage1_16[219]},
      {stage2_16[105]}
   );
   gpc1_1 gpc7672 (
      {stage1_16[220]},
      {stage2_16[106]}
   );
   gpc1_1 gpc7673 (
      {stage1_16[221]},
      {stage2_16[107]}
   );
   gpc1_1 gpc7674 (
      {stage1_16[222]},
      {stage2_16[108]}
   );
   gpc1_1 gpc7675 (
      {stage1_16[223]},
      {stage2_16[109]}
   );
   gpc1_1 gpc7676 (
      {stage1_18[204]},
      {stage2_18[124]}
   );
   gpc1_1 gpc7677 (
      {stage1_18[205]},
      {stage2_18[125]}
   );
   gpc1_1 gpc7678 (
      {stage1_18[206]},
      {stage2_18[126]}
   );
   gpc1_1 gpc7679 (
      {stage1_18[207]},
      {stage2_18[127]}
   );
   gpc1_1 gpc7680 (
      {stage1_18[208]},
      {stage2_18[128]}
   );
   gpc1_1 gpc7681 (
      {stage1_18[209]},
      {stage2_18[129]}
   );
   gpc1_1 gpc7682 (
      {stage1_18[210]},
      {stage2_18[130]}
   );
   gpc1_1 gpc7683 (
      {stage1_18[211]},
      {stage2_18[131]}
   );
   gpc1_1 gpc7684 (
      {stage1_18[212]},
      {stage2_18[132]}
   );
   gpc1_1 gpc7685 (
      {stage1_18[213]},
      {stage2_18[133]}
   );
   gpc1_1 gpc7686 (
      {stage1_18[214]},
      {stage2_18[134]}
   );
   gpc1_1 gpc7687 (
      {stage1_18[215]},
      {stage2_18[135]}
   );
   gpc1_1 gpc7688 (
      {stage1_18[216]},
      {stage2_18[136]}
   );
   gpc1_1 gpc7689 (
      {stage1_18[217]},
      {stage2_18[137]}
   );
   gpc1_1 gpc7690 (
      {stage1_18[218]},
      {stage2_18[138]}
   );
   gpc1_1 gpc7691 (
      {stage1_18[219]},
      {stage2_18[139]}
   );
   gpc1_1 gpc7692 (
      {stage1_18[220]},
      {stage2_18[140]}
   );
   gpc1_1 gpc7693 (
      {stage1_18[221]},
      {stage2_18[141]}
   );
   gpc1_1 gpc7694 (
      {stage1_18[222]},
      {stage2_18[142]}
   );
   gpc1_1 gpc7695 (
      {stage1_18[223]},
      {stage2_18[143]}
   );
   gpc1_1 gpc7696 (
      {stage1_18[224]},
      {stage2_18[144]}
   );
   gpc1_1 gpc7697 (
      {stage1_18[225]},
      {stage2_18[145]}
   );
   gpc1_1 gpc7698 (
      {stage1_18[226]},
      {stage2_18[146]}
   );
   gpc1_1 gpc7699 (
      {stage1_18[227]},
      {stage2_18[147]}
   );
   gpc1_1 gpc7700 (
      {stage1_18[228]},
      {stage2_18[148]}
   );
   gpc1_1 gpc7701 (
      {stage1_18[229]},
      {stage2_18[149]}
   );
   gpc1_1 gpc7702 (
      {stage1_18[230]},
      {stage2_18[150]}
   );
   gpc1_1 gpc7703 (
      {stage1_18[231]},
      {stage2_18[151]}
   );
   gpc1_1 gpc7704 (
      {stage1_18[232]},
      {stage2_18[152]}
   );
   gpc1_1 gpc7705 (
      {stage1_18[233]},
      {stage2_18[153]}
   );
   gpc1_1 gpc7706 (
      {stage1_18[234]},
      {stage2_18[154]}
   );
   gpc1_1 gpc7707 (
      {stage1_18[235]},
      {stage2_18[155]}
   );
   gpc1_1 gpc7708 (
      {stage1_18[236]},
      {stage2_18[156]}
   );
   gpc1_1 gpc7709 (
      {stage1_18[237]},
      {stage2_18[157]}
   );
   gpc1_1 gpc7710 (
      {stage1_18[238]},
      {stage2_18[158]}
   );
   gpc1_1 gpc7711 (
      {stage1_18[239]},
      {stage2_18[159]}
   );
   gpc1_1 gpc7712 (
      {stage1_18[240]},
      {stage2_18[160]}
   );
   gpc1_1 gpc7713 (
      {stage1_18[241]},
      {stage2_18[161]}
   );
   gpc1_1 gpc7714 (
      {stage1_19[201]},
      {stage2_19[76]}
   );
   gpc1_1 gpc7715 (
      {stage1_19[202]},
      {stage2_19[77]}
   );
   gpc1_1 gpc7716 (
      {stage1_19[203]},
      {stage2_19[78]}
   );
   gpc1_1 gpc7717 (
      {stage1_19[204]},
      {stage2_19[79]}
   );
   gpc1_1 gpc7718 (
      {stage1_19[205]},
      {stage2_19[80]}
   );
   gpc1_1 gpc7719 (
      {stage1_19[206]},
      {stage2_19[81]}
   );
   gpc1_1 gpc7720 (
      {stage1_19[207]},
      {stage2_19[82]}
   );
   gpc1_1 gpc7721 (
      {stage1_19[208]},
      {stage2_19[83]}
   );
   gpc1_1 gpc7722 (
      {stage1_19[209]},
      {stage2_19[84]}
   );
   gpc1_1 gpc7723 (
      {stage1_19[210]},
      {stage2_19[85]}
   );
   gpc1_1 gpc7724 (
      {stage1_19[211]},
      {stage2_19[86]}
   );
   gpc1_1 gpc7725 (
      {stage1_19[212]},
      {stage2_19[87]}
   );
   gpc1_1 gpc7726 (
      {stage1_19[213]},
      {stage2_19[88]}
   );
   gpc1_1 gpc7727 (
      {stage1_19[214]},
      {stage2_19[89]}
   );
   gpc1_1 gpc7728 (
      {stage1_19[215]},
      {stage2_19[90]}
   );
   gpc1_1 gpc7729 (
      {stage1_19[216]},
      {stage2_19[91]}
   );
   gpc1_1 gpc7730 (
      {stage1_19[217]},
      {stage2_19[92]}
   );
   gpc1_1 gpc7731 (
      {stage1_19[218]},
      {stage2_19[93]}
   );
   gpc1_1 gpc7732 (
      {stage1_20[227]},
      {stage2_20[71]}
   );
   gpc1_1 gpc7733 (
      {stage1_20[228]},
      {stage2_20[72]}
   );
   gpc1_1 gpc7734 (
      {stage1_20[229]},
      {stage2_20[73]}
   );
   gpc1_1 gpc7735 (
      {stage1_20[230]},
      {stage2_20[74]}
   );
   gpc1_1 gpc7736 (
      {stage1_20[231]},
      {stage2_20[75]}
   );
   gpc1_1 gpc7737 (
      {stage1_20[232]},
      {stage2_20[76]}
   );
   gpc1_1 gpc7738 (
      {stage1_20[233]},
      {stage2_20[77]}
   );
   gpc1_1 gpc7739 (
      {stage1_20[234]},
      {stage2_20[78]}
   );
   gpc1_1 gpc7740 (
      {stage1_20[235]},
      {stage2_20[79]}
   );
   gpc1_1 gpc7741 (
      {stage1_20[236]},
      {stage2_20[80]}
   );
   gpc1_1 gpc7742 (
      {stage1_20[237]},
      {stage2_20[81]}
   );
   gpc1_1 gpc7743 (
      {stage1_20[238]},
      {stage2_20[82]}
   );
   gpc1_1 gpc7744 (
      {stage1_20[239]},
      {stage2_20[83]}
   );
   gpc1_1 gpc7745 (
      {stage1_20[240]},
      {stage2_20[84]}
   );
   gpc1_1 gpc7746 (
      {stage1_20[241]},
      {stage2_20[85]}
   );
   gpc1_1 gpc7747 (
      {stage1_20[242]},
      {stage2_20[86]}
   );
   gpc1_1 gpc7748 (
      {stage1_20[243]},
      {stage2_20[87]}
   );
   gpc1_1 gpc7749 (
      {stage1_21[186]},
      {stage2_21[93]}
   );
   gpc1_1 gpc7750 (
      {stage1_21[187]},
      {stage2_21[94]}
   );
   gpc1_1 gpc7751 (
      {stage1_21[188]},
      {stage2_21[95]}
   );
   gpc1_1 gpc7752 (
      {stage1_21[189]},
      {stage2_21[96]}
   );
   gpc1_1 gpc7753 (
      {stage1_21[190]},
      {stage2_21[97]}
   );
   gpc1_1 gpc7754 (
      {stage1_21[191]},
      {stage2_21[98]}
   );
   gpc1_1 gpc7755 (
      {stage1_21[192]},
      {stage2_21[99]}
   );
   gpc1_1 gpc7756 (
      {stage1_21[193]},
      {stage2_21[100]}
   );
   gpc1_1 gpc7757 (
      {stage1_21[194]},
      {stage2_21[101]}
   );
   gpc1_1 gpc7758 (
      {stage1_21[195]},
      {stage2_21[102]}
   );
   gpc1_1 gpc7759 (
      {stage1_21[196]},
      {stage2_21[103]}
   );
   gpc1_1 gpc7760 (
      {stage1_21[197]},
      {stage2_21[104]}
   );
   gpc1_1 gpc7761 (
      {stage1_21[198]},
      {stage2_21[105]}
   );
   gpc1_1 gpc7762 (
      {stage1_21[199]},
      {stage2_21[106]}
   );
   gpc1_1 gpc7763 (
      {stage1_21[200]},
      {stage2_21[107]}
   );
   gpc1_1 gpc7764 (
      {stage1_21[201]},
      {stage2_21[108]}
   );
   gpc1_1 gpc7765 (
      {stage1_21[202]},
      {stage2_21[109]}
   );
   gpc1_1 gpc7766 (
      {stage1_21[203]},
      {stage2_21[110]}
   );
   gpc1_1 gpc7767 (
      {stage1_21[204]},
      {stage2_21[111]}
   );
   gpc1_1 gpc7768 (
      {stage1_22[194]},
      {stage2_22[103]}
   );
   gpc1_1 gpc7769 (
      {stage1_22[195]},
      {stage2_22[104]}
   );
   gpc1_1 gpc7770 (
      {stage1_22[196]},
      {stage2_22[105]}
   );
   gpc1_1 gpc7771 (
      {stage1_22[197]},
      {stage2_22[106]}
   );
   gpc1_1 gpc7772 (
      {stage1_22[198]},
      {stage2_22[107]}
   );
   gpc1_1 gpc7773 (
      {stage1_22[199]},
      {stage2_22[108]}
   );
   gpc1_1 gpc7774 (
      {stage1_22[200]},
      {stage2_22[109]}
   );
   gpc1_1 gpc7775 (
      {stage1_23[290]},
      {stage2_23[89]}
   );
   gpc1_1 gpc7776 (
      {stage1_23[291]},
      {stage2_23[90]}
   );
   gpc1_1 gpc7777 (
      {stage1_23[292]},
      {stage2_23[91]}
   );
   gpc1_1 gpc7778 (
      {stage1_23[293]},
      {stage2_23[92]}
   );
   gpc1_1 gpc7779 (
      {stage1_23[294]},
      {stage2_23[93]}
   );
   gpc1_1 gpc7780 (
      {stage1_23[295]},
      {stage2_23[94]}
   );
   gpc1_1 gpc7781 (
      {stage1_23[296]},
      {stage2_23[95]}
   );
   gpc1_1 gpc7782 (
      {stage1_23[297]},
      {stage2_23[96]}
   );
   gpc1_1 gpc7783 (
      {stage1_23[298]},
      {stage2_23[97]}
   );
   gpc1_1 gpc7784 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc7785 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc7786 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc7787 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc7788 (
      {stage1_25[184]},
      {stage2_25[96]}
   );
   gpc1_1 gpc7789 (
      {stage1_25[185]},
      {stage2_25[97]}
   );
   gpc1_1 gpc7790 (
      {stage1_25[186]},
      {stage2_25[98]}
   );
   gpc1_1 gpc7791 (
      {stage1_25[187]},
      {stage2_25[99]}
   );
   gpc1_1 gpc7792 (
      {stage1_25[188]},
      {stage2_25[100]}
   );
   gpc1_1 gpc7793 (
      {stage1_25[189]},
      {stage2_25[101]}
   );
   gpc1_1 gpc7794 (
      {stage1_25[190]},
      {stage2_25[102]}
   );
   gpc1_1 gpc7795 (
      {stage1_25[191]},
      {stage2_25[103]}
   );
   gpc1_1 gpc7796 (
      {stage1_25[192]},
      {stage2_25[104]}
   );
   gpc1_1 gpc7797 (
      {stage1_25[193]},
      {stage2_25[105]}
   );
   gpc1_1 gpc7798 (
      {stage1_25[194]},
      {stage2_25[106]}
   );
   gpc1_1 gpc7799 (
      {stage1_25[195]},
      {stage2_25[107]}
   );
   gpc1_1 gpc7800 (
      {stage1_25[196]},
      {stage2_25[108]}
   );
   gpc1_1 gpc7801 (
      {stage1_25[197]},
      {stage2_25[109]}
   );
   gpc1_1 gpc7802 (
      {stage1_25[198]},
      {stage2_25[110]}
   );
   gpc1_1 gpc7803 (
      {stage1_25[199]},
      {stage2_25[111]}
   );
   gpc1_1 gpc7804 (
      {stage1_25[200]},
      {stage2_25[112]}
   );
   gpc1_1 gpc7805 (
      {stage1_25[201]},
      {stage2_25[113]}
   );
   gpc1_1 gpc7806 (
      {stage1_25[202]},
      {stage2_25[114]}
   );
   gpc1_1 gpc7807 (
      {stage1_25[203]},
      {stage2_25[115]}
   );
   gpc1_1 gpc7808 (
      {stage1_25[204]},
      {stage2_25[116]}
   );
   gpc1_1 gpc7809 (
      {stage1_25[205]},
      {stage2_25[117]}
   );
   gpc1_1 gpc7810 (
      {stage1_25[206]},
      {stage2_25[118]}
   );
   gpc1_1 gpc7811 (
      {stage1_25[207]},
      {stage2_25[119]}
   );
   gpc1_1 gpc7812 (
      {stage1_25[208]},
      {stage2_25[120]}
   );
   gpc1_1 gpc7813 (
      {stage1_25[209]},
      {stage2_25[121]}
   );
   gpc1_1 gpc7814 (
      {stage1_25[210]},
      {stage2_25[122]}
   );
   gpc1_1 gpc7815 (
      {stage1_26[154]},
      {stage2_26[96]}
   );
   gpc1_1 gpc7816 (
      {stage1_26[155]},
      {stage2_26[97]}
   );
   gpc1_1 gpc7817 (
      {stage1_26[156]},
      {stage2_26[98]}
   );
   gpc1_1 gpc7818 (
      {stage1_26[157]},
      {stage2_26[99]}
   );
   gpc1_1 gpc7819 (
      {stage1_26[158]},
      {stage2_26[100]}
   );
   gpc1_1 gpc7820 (
      {stage1_26[159]},
      {stage2_26[101]}
   );
   gpc1_1 gpc7821 (
      {stage1_26[160]},
      {stage2_26[102]}
   );
   gpc1_1 gpc7822 (
      {stage1_26[161]},
      {stage2_26[103]}
   );
   gpc1_1 gpc7823 (
      {stage1_26[162]},
      {stage2_26[104]}
   );
   gpc1_1 gpc7824 (
      {stage1_26[163]},
      {stage2_26[105]}
   );
   gpc1_1 gpc7825 (
      {stage1_26[164]},
      {stage2_26[106]}
   );
   gpc1_1 gpc7826 (
      {stage1_26[165]},
      {stage2_26[107]}
   );
   gpc1_1 gpc7827 (
      {stage1_26[166]},
      {stage2_26[108]}
   );
   gpc1_1 gpc7828 (
      {stage1_26[167]},
      {stage2_26[109]}
   );
   gpc1_1 gpc7829 (
      {stage1_26[168]},
      {stage2_26[110]}
   );
   gpc1_1 gpc7830 (
      {stage1_26[169]},
      {stage2_26[111]}
   );
   gpc1_1 gpc7831 (
      {stage1_26[170]},
      {stage2_26[112]}
   );
   gpc1_1 gpc7832 (
      {stage1_26[171]},
      {stage2_26[113]}
   );
   gpc1_1 gpc7833 (
      {stage1_26[172]},
      {stage2_26[114]}
   );
   gpc1_1 gpc7834 (
      {stage1_26[173]},
      {stage2_26[115]}
   );
   gpc1_1 gpc7835 (
      {stage1_26[174]},
      {stage2_26[116]}
   );
   gpc1_1 gpc7836 (
      {stage1_26[175]},
      {stage2_26[117]}
   );
   gpc1_1 gpc7837 (
      {stage1_26[176]},
      {stage2_26[118]}
   );
   gpc1_1 gpc7838 (
      {stage1_26[177]},
      {stage2_26[119]}
   );
   gpc1_1 gpc7839 (
      {stage1_26[178]},
      {stage2_26[120]}
   );
   gpc1_1 gpc7840 (
      {stage1_26[179]},
      {stage2_26[121]}
   );
   gpc1_1 gpc7841 (
      {stage1_26[180]},
      {stage2_26[122]}
   );
   gpc1_1 gpc7842 (
      {stage1_26[181]},
      {stage2_26[123]}
   );
   gpc1_1 gpc7843 (
      {stage1_26[182]},
      {stage2_26[124]}
   );
   gpc1_1 gpc7844 (
      {stage1_26[183]},
      {stage2_26[125]}
   );
   gpc1_1 gpc7845 (
      {stage1_26[184]},
      {stage2_26[126]}
   );
   gpc1_1 gpc7846 (
      {stage1_26[185]},
      {stage2_26[127]}
   );
   gpc1_1 gpc7847 (
      {stage1_26[186]},
      {stage2_26[128]}
   );
   gpc1_1 gpc7848 (
      {stage1_26[187]},
      {stage2_26[129]}
   );
   gpc1_1 gpc7849 (
      {stage1_26[188]},
      {stage2_26[130]}
   );
   gpc1_1 gpc7850 (
      {stage1_27[211]},
      {stage2_27[85]}
   );
   gpc1_1 gpc7851 (
      {stage1_28[240]},
      {stage2_28[71]}
   );
   gpc1_1 gpc7852 (
      {stage1_28[241]},
      {stage2_28[72]}
   );
   gpc1_1 gpc7853 (
      {stage1_28[242]},
      {stage2_28[73]}
   );
   gpc1_1 gpc7854 (
      {stage1_28[243]},
      {stage2_28[74]}
   );
   gpc1_1 gpc7855 (
      {stage1_28[244]},
      {stage2_28[75]}
   );
   gpc1_1 gpc7856 (
      {stage1_28[245]},
      {stage2_28[76]}
   );
   gpc1_1 gpc7857 (
      {stage1_28[246]},
      {stage2_28[77]}
   );
   gpc1_1 gpc7858 (
      {stage1_28[247]},
      {stage2_28[78]}
   );
   gpc1_1 gpc7859 (
      {stage1_28[248]},
      {stage2_28[79]}
   );
   gpc1_1 gpc7860 (
      {stage1_29[186]},
      {stage2_29[77]}
   );
   gpc1_1 gpc7861 (
      {stage1_29[187]},
      {stage2_29[78]}
   );
   gpc1_1 gpc7862 (
      {stage1_29[188]},
      {stage2_29[79]}
   );
   gpc1_1 gpc7863 (
      {stage1_29[189]},
      {stage2_29[80]}
   );
   gpc1_1 gpc7864 (
      {stage1_29[190]},
      {stage2_29[81]}
   );
   gpc1_1 gpc7865 (
      {stage1_29[191]},
      {stage2_29[82]}
   );
   gpc1_1 gpc7866 (
      {stage1_29[192]},
      {stage2_29[83]}
   );
   gpc1_1 gpc7867 (
      {stage1_29[193]},
      {stage2_29[84]}
   );
   gpc1_1 gpc7868 (
      {stage1_29[194]},
      {stage2_29[85]}
   );
   gpc1_1 gpc7869 (
      {stage1_29[195]},
      {stage2_29[86]}
   );
   gpc1_1 gpc7870 (
      {stage1_29[196]},
      {stage2_29[87]}
   );
   gpc1_1 gpc7871 (
      {stage1_29[197]},
      {stage2_29[88]}
   );
   gpc1_1 gpc7872 (
      {stage1_29[198]},
      {stage2_29[89]}
   );
   gpc1_1 gpc7873 (
      {stage1_29[199]},
      {stage2_29[90]}
   );
   gpc1_1 gpc7874 (
      {stage1_29[200]},
      {stage2_29[91]}
   );
   gpc1_1 gpc7875 (
      {stage1_29[201]},
      {stage2_29[92]}
   );
   gpc1_1 gpc7876 (
      {stage1_29[202]},
      {stage2_29[93]}
   );
   gpc1_1 gpc7877 (
      {stage1_29[203]},
      {stage2_29[94]}
   );
   gpc1_1 gpc7878 (
      {stage1_29[204]},
      {stage2_29[95]}
   );
   gpc1_1 gpc7879 (
      {stage1_29[205]},
      {stage2_29[96]}
   );
   gpc1_1 gpc7880 (
      {stage1_29[206]},
      {stage2_29[97]}
   );
   gpc1_1 gpc7881 (
      {stage1_29[207]},
      {stage2_29[98]}
   );
   gpc1_1 gpc7882 (
      {stage1_29[208]},
      {stage2_29[99]}
   );
   gpc1_1 gpc7883 (
      {stage1_29[209]},
      {stage2_29[100]}
   );
   gpc1_1 gpc7884 (
      {stage1_29[210]},
      {stage2_29[101]}
   );
   gpc1_1 gpc7885 (
      {stage1_29[211]},
      {stage2_29[102]}
   );
   gpc1_1 gpc7886 (
      {stage1_29[212]},
      {stage2_29[103]}
   );
   gpc1_1 gpc7887 (
      {stage1_29[213]},
      {stage2_29[104]}
   );
   gpc1_1 gpc7888 (
      {stage1_29[214]},
      {stage2_29[105]}
   );
   gpc1_1 gpc7889 (
      {stage1_29[215]},
      {stage2_29[106]}
   );
   gpc1_1 gpc7890 (
      {stage1_29[216]},
      {stage2_29[107]}
   );
   gpc1_1 gpc7891 (
      {stage1_29[217]},
      {stage2_29[108]}
   );
   gpc1_1 gpc7892 (
      {stage1_29[218]},
      {stage2_29[109]}
   );
   gpc1_1 gpc7893 (
      {stage1_29[219]},
      {stage2_29[110]}
   );
   gpc1_1 gpc7894 (
      {stage1_29[220]},
      {stage2_29[111]}
   );
   gpc1_1 gpc7895 (
      {stage1_30[232]},
      {stage2_30[99]}
   );
   gpc1_1 gpc7896 (
      {stage1_31[180]},
      {stage2_31[96]}
   );
   gpc1_1 gpc7897 (
      {stage1_31[181]},
      {stage2_31[97]}
   );
   gpc1_1 gpc7898 (
      {stage1_31[182]},
      {stage2_31[98]}
   );
   gpc1_1 gpc7899 (
      {stage1_31[183]},
      {stage2_31[99]}
   );
   gpc1_1 gpc7900 (
      {stage1_31[184]},
      {stage2_31[100]}
   );
   gpc1_1 gpc7901 (
      {stage1_31[185]},
      {stage2_31[101]}
   );
   gpc1_1 gpc7902 (
      {stage1_31[186]},
      {stage2_31[102]}
   );
   gpc1_1 gpc7903 (
      {stage1_31[187]},
      {stage2_31[103]}
   );
   gpc1_1 gpc7904 (
      {stage1_31[188]},
      {stage2_31[104]}
   );
   gpc1_1 gpc7905 (
      {stage1_31[189]},
      {stage2_31[105]}
   );
   gpc1_1 gpc7906 (
      {stage1_31[190]},
      {stage2_31[106]}
   );
   gpc1_1 gpc7907 (
      {stage1_31[191]},
      {stage2_31[107]}
   );
   gpc1_1 gpc7908 (
      {stage1_31[192]},
      {stage2_31[108]}
   );
   gpc1_1 gpc7909 (
      {stage1_31[193]},
      {stage2_31[109]}
   );
   gpc1_1 gpc7910 (
      {stage1_31[194]},
      {stage2_31[110]}
   );
   gpc1_1 gpc7911 (
      {stage1_31[195]},
      {stage2_31[111]}
   );
   gpc1_1 gpc7912 (
      {stage1_31[196]},
      {stage2_31[112]}
   );
   gpc1_1 gpc7913 (
      {stage1_31[197]},
      {stage2_31[113]}
   );
   gpc1_1 gpc7914 (
      {stage1_31[198]},
      {stage2_31[114]}
   );
   gpc1_1 gpc7915 (
      {stage1_31[199]},
      {stage2_31[115]}
   );
   gpc1_1 gpc7916 (
      {stage1_31[200]},
      {stage2_31[116]}
   );
   gpc1_1 gpc7917 (
      {stage1_31[201]},
      {stage2_31[117]}
   );
   gpc1_1 gpc7918 (
      {stage1_31[202]},
      {stage2_31[118]}
   );
   gpc1_1 gpc7919 (
      {stage1_31[203]},
      {stage2_31[119]}
   );
   gpc1_1 gpc7920 (
      {stage1_31[204]},
      {stage2_31[120]}
   );
   gpc1_1 gpc7921 (
      {stage1_31[205]},
      {stage2_31[121]}
   );
   gpc1_1 gpc7922 (
      {stage1_31[206]},
      {stage2_31[122]}
   );
   gpc1_1 gpc7923 (
      {stage1_31[207]},
      {stage2_31[123]}
   );
   gpc1_1 gpc7924 (
      {stage1_31[208]},
      {stage2_31[124]}
   );
   gpc1_1 gpc7925 (
      {stage1_31[209]},
      {stage2_31[125]}
   );
   gpc1_1 gpc7926 (
      {stage1_31[210]},
      {stage2_31[126]}
   );
   gpc1_1 gpc7927 (
      {stage1_31[211]},
      {stage2_31[127]}
   );
   gpc1_1 gpc7928 (
      {stage1_32[404]},
      {stage2_32[107]}
   );
   gpc1_1 gpc7929 (
      {stage1_32[405]},
      {stage2_32[108]}
   );
   gpc1_1 gpc7930 (
      {stage1_32[406]},
      {stage2_32[109]}
   );
   gpc1_1 gpc7931 (
      {stage1_32[407]},
      {stage2_32[110]}
   );
   gpc1_1 gpc7932 (
      {stage1_32[408]},
      {stage2_32[111]}
   );
   gpc1_1 gpc7933 (
      {stage1_32[409]},
      {stage2_32[112]}
   );
   gpc1_1 gpc7934 (
      {stage1_32[410]},
      {stage2_32[113]}
   );
   gpc1_1 gpc7935 (
      {stage1_32[411]},
      {stage2_32[114]}
   );
   gpc1_1 gpc7936 (
      {stage1_32[412]},
      {stage2_32[115]}
   );
   gpc1_1 gpc7937 (
      {stage1_32[413]},
      {stage2_32[116]}
   );
   gpc1_1 gpc7938 (
      {stage1_32[414]},
      {stage2_32[117]}
   );
   gpc1_1 gpc7939 (
      {stage1_34[242]},
      {stage2_34[102]}
   );
   gpc1_1 gpc7940 (
      {stage1_34[243]},
      {stage2_34[103]}
   );
   gpc1_1 gpc7941 (
      {stage1_34[244]},
      {stage2_34[104]}
   );
   gpc1_1 gpc7942 (
      {stage1_34[245]},
      {stage2_34[105]}
   );
   gpc1_1 gpc7943 (
      {stage1_34[246]},
      {stage2_34[106]}
   );
   gpc1_1 gpc7944 (
      {stage1_34[247]},
      {stage2_34[107]}
   );
   gpc1_1 gpc7945 (
      {stage1_34[248]},
      {stage2_34[108]}
   );
   gpc1_1 gpc7946 (
      {stage1_34[249]},
      {stage2_34[109]}
   );
   gpc1_1 gpc7947 (
      {stage1_34[250]},
      {stage2_34[110]}
   );
   gpc1_1 gpc7948 (
      {stage1_34[251]},
      {stage2_34[111]}
   );
   gpc1_1 gpc7949 (
      {stage1_34[252]},
      {stage2_34[112]}
   );
   gpc1_1 gpc7950 (
      {stage1_34[253]},
      {stage2_34[113]}
   );
   gpc1_1 gpc7951 (
      {stage1_34[254]},
      {stage2_34[114]}
   );
   gpc1_1 gpc7952 (
      {stage1_34[255]},
      {stage2_34[115]}
   );
   gpc1_1 gpc7953 (
      {stage1_34[256]},
      {stage2_34[116]}
   );
   gpc1_1 gpc7954 (
      {stage1_34[257]},
      {stage2_34[117]}
   );
   gpc1_1 gpc7955 (
      {stage1_34[258]},
      {stage2_34[118]}
   );
   gpc1_1 gpc7956 (
      {stage1_34[259]},
      {stage2_34[119]}
   );
   gpc1_1 gpc7957 (
      {stage1_34[260]},
      {stage2_34[120]}
   );
   gpc1_1 gpc7958 (
      {stage1_34[261]},
      {stage2_34[121]}
   );
   gpc1_1 gpc7959 (
      {stage1_34[262]},
      {stage2_34[122]}
   );
   gpc1_1 gpc7960 (
      {stage1_34[263]},
      {stage2_34[123]}
   );
   gpc1_1 gpc7961 (
      {stage1_34[264]},
      {stage2_34[124]}
   );
   gpc1_1 gpc7962 (
      {stage1_34[265]},
      {stage2_34[125]}
   );
   gpc1_1 gpc7963 (
      {stage1_34[266]},
      {stage2_34[126]}
   );
   gpc1_1 gpc7964 (
      {stage1_34[267]},
      {stage2_34[127]}
   );
   gpc1_1 gpc7965 (
      {stage1_35[173]},
      {stage2_35[100]}
   );
   gpc1_1 gpc7966 (
      {stage1_35[174]},
      {stage2_35[101]}
   );
   gpc1_1 gpc7967 (
      {stage1_35[175]},
      {stage2_35[102]}
   );
   gpc1_1 gpc7968 (
      {stage1_35[176]},
      {stage2_35[103]}
   );
   gpc1_1 gpc7969 (
      {stage1_35[177]},
      {stage2_35[104]}
   );
   gpc1_1 gpc7970 (
      {stage1_35[178]},
      {stage2_35[105]}
   );
   gpc1_1 gpc7971 (
      {stage1_35[179]},
      {stage2_35[106]}
   );
   gpc1_1 gpc7972 (
      {stage1_35[180]},
      {stage2_35[107]}
   );
   gpc1_1 gpc7973 (
      {stage1_35[181]},
      {stage2_35[108]}
   );
   gpc1_1 gpc7974 (
      {stage1_35[182]},
      {stage2_35[109]}
   );
   gpc1_1 gpc7975 (
      {stage1_35[183]},
      {stage2_35[110]}
   );
   gpc1_1 gpc7976 (
      {stage1_35[184]},
      {stage2_35[111]}
   );
   gpc1_1 gpc7977 (
      {stage1_35[185]},
      {stage2_35[112]}
   );
   gpc1_1 gpc7978 (
      {stage1_35[186]},
      {stage2_35[113]}
   );
   gpc1_1 gpc7979 (
      {stage1_35[187]},
      {stage2_35[114]}
   );
   gpc1_1 gpc7980 (
      {stage1_35[188]},
      {stage2_35[115]}
   );
   gpc1_1 gpc7981 (
      {stage1_35[189]},
      {stage2_35[116]}
   );
   gpc1_1 gpc7982 (
      {stage1_35[190]},
      {stage2_35[117]}
   );
   gpc1_1 gpc7983 (
      {stage1_37[297]},
      {stage2_37[108]}
   );
   gpc1_1 gpc7984 (
      {stage1_37[298]},
      {stage2_37[109]}
   );
   gpc1_1 gpc7985 (
      {stage1_37[299]},
      {stage2_37[110]}
   );
   gpc1_1 gpc7986 (
      {stage1_37[300]},
      {stage2_37[111]}
   );
   gpc1_1 gpc7987 (
      {stage1_37[301]},
      {stage2_37[112]}
   );
   gpc1_1 gpc7988 (
      {stage1_37[302]},
      {stage2_37[113]}
   );
   gpc1_1 gpc7989 (
      {stage1_39[194]},
      {stage2_39[105]}
   );
   gpc1_1 gpc7990 (
      {stage1_39[195]},
      {stage2_39[106]}
   );
   gpc1_1 gpc7991 (
      {stage1_39[196]},
      {stage2_39[107]}
   );
   gpc1_1 gpc7992 (
      {stage1_40[203]},
      {stage2_40[113]}
   );
   gpc1_1 gpc7993 (
      {stage1_40[204]},
      {stage2_40[114]}
   );
   gpc1_1 gpc7994 (
      {stage1_40[205]},
      {stage2_40[115]}
   );
   gpc1_1 gpc7995 (
      {stage1_40[206]},
      {stage2_40[116]}
   );
   gpc1_1 gpc7996 (
      {stage1_40[207]},
      {stage2_40[117]}
   );
   gpc1_1 gpc7997 (
      {stage1_40[208]},
      {stage2_40[118]}
   );
   gpc1_1 gpc7998 (
      {stage1_40[209]},
      {stage2_40[119]}
   );
   gpc1_1 gpc7999 (
      {stage1_40[210]},
      {stage2_40[120]}
   );
   gpc1_1 gpc8000 (
      {stage1_40[211]},
      {stage2_40[121]}
   );
   gpc1_1 gpc8001 (
      {stage1_40[212]},
      {stage2_40[122]}
   );
   gpc1_1 gpc8002 (
      {stage1_40[213]},
      {stage2_40[123]}
   );
   gpc1_1 gpc8003 (
      {stage1_40[214]},
      {stage2_40[124]}
   );
   gpc1_1 gpc8004 (
      {stage1_40[215]},
      {stage2_40[125]}
   );
   gpc1_1 gpc8005 (
      {stage1_40[216]},
      {stage2_40[126]}
   );
   gpc1_1 gpc8006 (
      {stage1_40[217]},
      {stage2_40[127]}
   );
   gpc1_1 gpc8007 (
      {stage1_40[218]},
      {stage2_40[128]}
   );
   gpc1_1 gpc8008 (
      {stage1_40[219]},
      {stage2_40[129]}
   );
   gpc1_1 gpc8009 (
      {stage1_40[220]},
      {stage2_40[130]}
   );
   gpc1_1 gpc8010 (
      {stage1_40[221]},
      {stage2_40[131]}
   );
   gpc1_1 gpc8011 (
      {stage1_40[222]},
      {stage2_40[132]}
   );
   gpc1_1 gpc8012 (
      {stage1_40[223]},
      {stage2_40[133]}
   );
   gpc1_1 gpc8013 (
      {stage1_40[224]},
      {stage2_40[134]}
   );
   gpc1_1 gpc8014 (
      {stage1_40[225]},
      {stage2_40[135]}
   );
   gpc1_1 gpc8015 (
      {stage1_40[226]},
      {stage2_40[136]}
   );
   gpc1_1 gpc8016 (
      {stage1_40[227]},
      {stage2_40[137]}
   );
   gpc1_1 gpc8017 (
      {stage1_40[228]},
      {stage2_40[138]}
   );
   gpc1_1 gpc8018 (
      {stage1_40[229]},
      {stage2_40[139]}
   );
   gpc1_1 gpc8019 (
      {stage1_41[252]},
      {stage2_41[98]}
   );
   gpc1_1 gpc8020 (
      {stage1_41[253]},
      {stage2_41[99]}
   );
   gpc1_1 gpc8021 (
      {stage1_41[254]},
      {stage2_41[100]}
   );
   gpc1_1 gpc8022 (
      {stage1_41[255]},
      {stage2_41[101]}
   );
   gpc1_1 gpc8023 (
      {stage1_41[256]},
      {stage2_41[102]}
   );
   gpc1_1 gpc8024 (
      {stage1_41[257]},
      {stage2_41[103]}
   );
   gpc1_1 gpc8025 (
      {stage1_41[258]},
      {stage2_41[104]}
   );
   gpc1_1 gpc8026 (
      {stage1_41[259]},
      {stage2_41[105]}
   );
   gpc1_1 gpc8027 (
      {stage1_41[260]},
      {stage2_41[106]}
   );
   gpc1_1 gpc8028 (
      {stage1_41[261]},
      {stage2_41[107]}
   );
   gpc1_1 gpc8029 (
      {stage1_41[262]},
      {stage2_41[108]}
   );
   gpc1_1 gpc8030 (
      {stage1_41[263]},
      {stage2_41[109]}
   );
   gpc1_1 gpc8031 (
      {stage1_41[264]},
      {stage2_41[110]}
   );
   gpc1_1 gpc8032 (
      {stage1_41[265]},
      {stage2_41[111]}
   );
   gpc1_1 gpc8033 (
      {stage1_41[266]},
      {stage2_41[112]}
   );
   gpc1_1 gpc8034 (
      {stage1_41[267]},
      {stage2_41[113]}
   );
   gpc1_1 gpc8035 (
      {stage1_41[268]},
      {stage2_41[114]}
   );
   gpc1_1 gpc8036 (
      {stage1_41[269]},
      {stage2_41[115]}
   );
   gpc1_1 gpc8037 (
      {stage1_41[270]},
      {stage2_41[116]}
   );
   gpc1_1 gpc8038 (
      {stage1_41[271]},
      {stage2_41[117]}
   );
   gpc1_1 gpc8039 (
      {stage1_41[272]},
      {stage2_41[118]}
   );
   gpc1_1 gpc8040 (
      {stage1_41[273]},
      {stage2_41[119]}
   );
   gpc1_1 gpc8041 (
      {stage1_41[274]},
      {stage2_41[120]}
   );
   gpc1_1 gpc8042 (
      {stage1_41[275]},
      {stage2_41[121]}
   );
   gpc1_1 gpc8043 (
      {stage1_41[276]},
      {stage2_41[122]}
   );
   gpc1_1 gpc8044 (
      {stage1_42[228]},
      {stage2_42[81]}
   );
   gpc1_1 gpc8045 (
      {stage1_43[218]},
      {stage2_43[85]}
   );
   gpc1_1 gpc8046 (
      {stage1_43[219]},
      {stage2_43[86]}
   );
   gpc1_1 gpc8047 (
      {stage1_43[220]},
      {stage2_43[87]}
   );
   gpc1_1 gpc8048 (
      {stage1_43[221]},
      {stage2_43[88]}
   );
   gpc1_1 gpc8049 (
      {stage1_43[222]},
      {stage2_43[89]}
   );
   gpc1_1 gpc8050 (
      {stage1_43[223]},
      {stage2_43[90]}
   );
   gpc1_1 gpc8051 (
      {stage1_43[224]},
      {stage2_43[91]}
   );
   gpc1_1 gpc8052 (
      {stage1_43[225]},
      {stage2_43[92]}
   );
   gpc1_1 gpc8053 (
      {stage1_43[226]},
      {stage2_43[93]}
   );
   gpc1_1 gpc8054 (
      {stage1_43[227]},
      {stage2_43[94]}
   );
   gpc1_1 gpc8055 (
      {stage1_43[228]},
      {stage2_43[95]}
   );
   gpc1_1 gpc8056 (
      {stage1_43[229]},
      {stage2_43[96]}
   );
   gpc1_1 gpc8057 (
      {stage1_43[230]},
      {stage2_43[97]}
   );
   gpc1_1 gpc8058 (
      {stage1_43[231]},
      {stage2_43[98]}
   );
   gpc1_1 gpc8059 (
      {stage1_43[232]},
      {stage2_43[99]}
   );
   gpc1_1 gpc8060 (
      {stage1_43[233]},
      {stage2_43[100]}
   );
   gpc1_1 gpc8061 (
      {stage1_43[234]},
      {stage2_43[101]}
   );
   gpc1_1 gpc8062 (
      {stage1_43[235]},
      {stage2_43[102]}
   );
   gpc1_1 gpc8063 (
      {stage1_43[236]},
      {stage2_43[103]}
   );
   gpc1_1 gpc8064 (
      {stage1_43[237]},
      {stage2_43[104]}
   );
   gpc1_1 gpc8065 (
      {stage1_43[238]},
      {stage2_43[105]}
   );
   gpc1_1 gpc8066 (
      {stage1_43[239]},
      {stage2_43[106]}
   );
   gpc1_1 gpc8067 (
      {stage1_43[240]},
      {stage2_43[107]}
   );
   gpc1_1 gpc8068 (
      {stage1_43[241]},
      {stage2_43[108]}
   );
   gpc1_1 gpc8069 (
      {stage1_43[242]},
      {stage2_43[109]}
   );
   gpc1_1 gpc8070 (
      {stage1_43[243]},
      {stage2_43[110]}
   );
   gpc1_1 gpc8071 (
      {stage1_44[244]},
      {stage2_44[113]}
   );
   gpc1_1 gpc8072 (
      {stage1_44[245]},
      {stage2_44[114]}
   );
   gpc1_1 gpc8073 (
      {stage1_44[246]},
      {stage2_44[115]}
   );
   gpc1_1 gpc8074 (
      {stage1_44[247]},
      {stage2_44[116]}
   );
   gpc1_1 gpc8075 (
      {stage1_44[248]},
      {stage2_44[117]}
   );
   gpc1_1 gpc8076 (
      {stage1_44[249]},
      {stage2_44[118]}
   );
   gpc1_1 gpc8077 (
      {stage1_44[250]},
      {stage2_44[119]}
   );
   gpc1_1 gpc8078 (
      {stage1_44[251]},
      {stage2_44[120]}
   );
   gpc1_1 gpc8079 (
      {stage1_44[252]},
      {stage2_44[121]}
   );
   gpc1_1 gpc8080 (
      {stage1_44[253]},
      {stage2_44[122]}
   );
   gpc1_1 gpc8081 (
      {stage1_44[254]},
      {stage2_44[123]}
   );
   gpc1_1 gpc8082 (
      {stage1_44[255]},
      {stage2_44[124]}
   );
   gpc1_1 gpc8083 (
      {stage1_44[256]},
      {stage2_44[125]}
   );
   gpc1_1 gpc8084 (
      {stage1_44[257]},
      {stage2_44[126]}
   );
   gpc1_1 gpc8085 (
      {stage1_44[258]},
      {stage2_44[127]}
   );
   gpc1_1 gpc8086 (
      {stage1_44[259]},
      {stage2_44[128]}
   );
   gpc1_1 gpc8087 (
      {stage1_44[260]},
      {stage2_44[129]}
   );
   gpc1_1 gpc8088 (
      {stage1_44[261]},
      {stage2_44[130]}
   );
   gpc1_1 gpc8089 (
      {stage1_44[262]},
      {stage2_44[131]}
   );
   gpc1_1 gpc8090 (
      {stage1_44[263]},
      {stage2_44[132]}
   );
   gpc1_1 gpc8091 (
      {stage1_44[264]},
      {stage2_44[133]}
   );
   gpc1_1 gpc8092 (
      {stage1_44[265]},
      {stage2_44[134]}
   );
   gpc1_1 gpc8093 (
      {stage1_44[266]},
      {stage2_44[135]}
   );
   gpc1_1 gpc8094 (
      {stage1_44[267]},
      {stage2_44[136]}
   );
   gpc1_1 gpc8095 (
      {stage1_44[268]},
      {stage2_44[137]}
   );
   gpc1_1 gpc8096 (
      {stage1_45[157]},
      {stage2_45[100]}
   );
   gpc1_1 gpc8097 (
      {stage1_45[158]},
      {stage2_45[101]}
   );
   gpc1_1 gpc8098 (
      {stage1_45[159]},
      {stage2_45[102]}
   );
   gpc1_1 gpc8099 (
      {stage1_45[160]},
      {stage2_45[103]}
   );
   gpc1_1 gpc8100 (
      {stage1_45[161]},
      {stage2_45[104]}
   );
   gpc1_1 gpc8101 (
      {stage1_45[162]},
      {stage2_45[105]}
   );
   gpc1_1 gpc8102 (
      {stage1_45[163]},
      {stage2_45[106]}
   );
   gpc1_1 gpc8103 (
      {stage1_45[164]},
      {stage2_45[107]}
   );
   gpc1_1 gpc8104 (
      {stage1_45[165]},
      {stage2_45[108]}
   );
   gpc1_1 gpc8105 (
      {stage1_45[166]},
      {stage2_45[109]}
   );
   gpc1_1 gpc8106 (
      {stage1_45[167]},
      {stage2_45[110]}
   );
   gpc1_1 gpc8107 (
      {stage1_45[168]},
      {stage2_45[111]}
   );
   gpc1_1 gpc8108 (
      {stage1_45[169]},
      {stage2_45[112]}
   );
   gpc1_1 gpc8109 (
      {stage1_45[170]},
      {stage2_45[113]}
   );
   gpc1_1 gpc8110 (
      {stage1_45[171]},
      {stage2_45[114]}
   );
   gpc1_1 gpc8111 (
      {stage1_45[172]},
      {stage2_45[115]}
   );
   gpc1_1 gpc8112 (
      {stage1_45[173]},
      {stage2_45[116]}
   );
   gpc1_1 gpc8113 (
      {stage1_45[174]},
      {stage2_45[117]}
   );
   gpc1_1 gpc8114 (
      {stage1_45[175]},
      {stage2_45[118]}
   );
   gpc1_1 gpc8115 (
      {stage1_45[176]},
      {stage2_45[119]}
   );
   gpc1_1 gpc8116 (
      {stage1_45[177]},
      {stage2_45[120]}
   );
   gpc1_1 gpc8117 (
      {stage1_45[178]},
      {stage2_45[121]}
   );
   gpc1_1 gpc8118 (
      {stage1_45[179]},
      {stage2_45[122]}
   );
   gpc1_1 gpc8119 (
      {stage1_45[180]},
      {stage2_45[123]}
   );
   gpc1_1 gpc8120 (
      {stage1_45[181]},
      {stage2_45[124]}
   );
   gpc1_1 gpc8121 (
      {stage1_45[182]},
      {stage2_45[125]}
   );
   gpc1_1 gpc8122 (
      {stage1_45[183]},
      {stage2_45[126]}
   );
   gpc1_1 gpc8123 (
      {stage1_45[184]},
      {stage2_45[127]}
   );
   gpc1_1 gpc8124 (
      {stage1_45[185]},
      {stage2_45[128]}
   );
   gpc1_1 gpc8125 (
      {stage1_45[186]},
      {stage2_45[129]}
   );
   gpc1_1 gpc8126 (
      {stage1_45[187]},
      {stage2_45[130]}
   );
   gpc1_1 gpc8127 (
      {stage1_45[188]},
      {stage2_45[131]}
   );
   gpc1_1 gpc8128 (
      {stage1_46[285]},
      {stage2_46[78]}
   );
   gpc1_1 gpc8129 (
      {stage1_46[286]},
      {stage2_46[79]}
   );
   gpc1_1 gpc8130 (
      {stage1_46[287]},
      {stage2_46[80]}
   );
   gpc1_1 gpc8131 (
      {stage1_46[288]},
      {stage2_46[81]}
   );
   gpc1_1 gpc8132 (
      {stage1_46[289]},
      {stage2_46[82]}
   );
   gpc1_1 gpc8133 (
      {stage1_46[290]},
      {stage2_46[83]}
   );
   gpc1_1 gpc8134 (
      {stage1_46[291]},
      {stage2_46[84]}
   );
   gpc1_1 gpc8135 (
      {stage1_46[292]},
      {stage2_46[85]}
   );
   gpc1_1 gpc8136 (
      {stage1_46[293]},
      {stage2_46[86]}
   );
   gpc1_1 gpc8137 (
      {stage1_46[294]},
      {stage2_46[87]}
   );
   gpc1_1 gpc8138 (
      {stage1_46[295]},
      {stage2_46[88]}
   );
   gpc1_1 gpc8139 (
      {stage1_46[296]},
      {stage2_46[89]}
   );
   gpc1_1 gpc8140 (
      {stage1_46[297]},
      {stage2_46[90]}
   );
   gpc1_1 gpc8141 (
      {stage1_46[298]},
      {stage2_46[91]}
   );
   gpc1_1 gpc8142 (
      {stage1_46[299]},
      {stage2_46[92]}
   );
   gpc1_1 gpc8143 (
      {stage1_47[270]},
      {stage2_47[100]}
   );
   gpc1_1 gpc8144 (
      {stage1_47[271]},
      {stage2_47[101]}
   );
   gpc1_1 gpc8145 (
      {stage1_47[272]},
      {stage2_47[102]}
   );
   gpc1_1 gpc8146 (
      {stage1_47[273]},
      {stage2_47[103]}
   );
   gpc1_1 gpc8147 (
      {stage1_47[274]},
      {stage2_47[104]}
   );
   gpc1_1 gpc8148 (
      {stage1_47[275]},
      {stage2_47[105]}
   );
   gpc1_1 gpc8149 (
      {stage1_47[276]},
      {stage2_47[106]}
   );
   gpc1_1 gpc8150 (
      {stage1_47[277]},
      {stage2_47[107]}
   );
   gpc1_1 gpc8151 (
      {stage1_48[166]},
      {stage2_48[109]}
   );
   gpc1_1 gpc8152 (
      {stage1_48[167]},
      {stage2_48[110]}
   );
   gpc1_1 gpc8153 (
      {stage1_48[168]},
      {stage2_48[111]}
   );
   gpc1_1 gpc8154 (
      {stage1_48[169]},
      {stage2_48[112]}
   );
   gpc1_1 gpc8155 (
      {stage1_48[170]},
      {stage2_48[113]}
   );
   gpc1_1 gpc8156 (
      {stage1_48[171]},
      {stage2_48[114]}
   );
   gpc1_1 gpc8157 (
      {stage1_48[172]},
      {stage2_48[115]}
   );
   gpc1_1 gpc8158 (
      {stage1_48[173]},
      {stage2_48[116]}
   );
   gpc1_1 gpc8159 (
      {stage1_48[174]},
      {stage2_48[117]}
   );
   gpc1_1 gpc8160 (
      {stage1_48[175]},
      {stage2_48[118]}
   );
   gpc1_1 gpc8161 (
      {stage1_48[176]},
      {stage2_48[119]}
   );
   gpc1_1 gpc8162 (
      {stage1_48[177]},
      {stage2_48[120]}
   );
   gpc1_1 gpc8163 (
      {stage1_48[178]},
      {stage2_48[121]}
   );
   gpc1_1 gpc8164 (
      {stage1_48[179]},
      {stage2_48[122]}
   );
   gpc1_1 gpc8165 (
      {stage1_48[180]},
      {stage2_48[123]}
   );
   gpc1_1 gpc8166 (
      {stage1_48[181]},
      {stage2_48[124]}
   );
   gpc1_1 gpc8167 (
      {stage1_48[182]},
      {stage2_48[125]}
   );
   gpc1_1 gpc8168 (
      {stage1_48[183]},
      {stage2_48[126]}
   );
   gpc1_1 gpc8169 (
      {stage1_48[184]},
      {stage2_48[127]}
   );
   gpc1_1 gpc8170 (
      {stage1_48[185]},
      {stage2_48[128]}
   );
   gpc1_1 gpc8171 (
      {stage1_48[186]},
      {stage2_48[129]}
   );
   gpc1_1 gpc8172 (
      {stage1_48[187]},
      {stage2_48[130]}
   );
   gpc1_1 gpc8173 (
      {stage1_48[188]},
      {stage2_48[131]}
   );
   gpc1_1 gpc8174 (
      {stage1_48[189]},
      {stage2_48[132]}
   );
   gpc1_1 gpc8175 (
      {stage1_48[190]},
      {stage2_48[133]}
   );
   gpc1_1 gpc8176 (
      {stage1_48[191]},
      {stage2_48[134]}
   );
   gpc1_1 gpc8177 (
      {stage1_48[192]},
      {stage2_48[135]}
   );
   gpc1_1 gpc8178 (
      {stage1_48[193]},
      {stage2_48[136]}
   );
   gpc1_1 gpc8179 (
      {stage1_48[194]},
      {stage2_48[137]}
   );
   gpc1_1 gpc8180 (
      {stage1_48[195]},
      {stage2_48[138]}
   );
   gpc1_1 gpc8181 (
      {stage1_48[196]},
      {stage2_48[139]}
   );
   gpc1_1 gpc8182 (
      {stage1_48[197]},
      {stage2_48[140]}
   );
   gpc1_1 gpc8183 (
      {stage1_48[198]},
      {stage2_48[141]}
   );
   gpc1_1 gpc8184 (
      {stage1_48[199]},
      {stage2_48[142]}
   );
   gpc1_1 gpc8185 (
      {stage1_48[200]},
      {stage2_48[143]}
   );
   gpc1_1 gpc8186 (
      {stage1_48[201]},
      {stage2_48[144]}
   );
   gpc1_1 gpc8187 (
      {stage1_48[202]},
      {stage2_48[145]}
   );
   gpc1_1 gpc8188 (
      {stage1_48[203]},
      {stage2_48[146]}
   );
   gpc1_1 gpc8189 (
      {stage1_48[204]},
      {stage2_48[147]}
   );
   gpc1_1 gpc8190 (
      {stage1_48[205]},
      {stage2_48[148]}
   );
   gpc1_1 gpc8191 (
      {stage1_48[206]},
      {stage2_48[149]}
   );
   gpc1_1 gpc8192 (
      {stage1_48[207]},
      {stage2_48[150]}
   );
   gpc1_1 gpc8193 (
      {stage1_48[208]},
      {stage2_48[151]}
   );
   gpc1_1 gpc8194 (
      {stage1_48[209]},
      {stage2_48[152]}
   );
   gpc1_1 gpc8195 (
      {stage1_48[210]},
      {stage2_48[153]}
   );
   gpc1_1 gpc8196 (
      {stage1_49[203]},
      {stage2_49[77]}
   );
   gpc1_1 gpc8197 (
      {stage1_49[204]},
      {stage2_49[78]}
   );
   gpc1_1 gpc8198 (
      {stage1_49[205]},
      {stage2_49[79]}
   );
   gpc1_1 gpc8199 (
      {stage1_49[206]},
      {stage2_49[80]}
   );
   gpc1_1 gpc8200 (
      {stage1_49[207]},
      {stage2_49[81]}
   );
   gpc1_1 gpc8201 (
      {stage1_49[208]},
      {stage2_49[82]}
   );
   gpc1_1 gpc8202 (
      {stage1_49[209]},
      {stage2_49[83]}
   );
   gpc1_1 gpc8203 (
      {stage1_49[210]},
      {stage2_49[84]}
   );
   gpc1_1 gpc8204 (
      {stage1_49[211]},
      {stage2_49[85]}
   );
   gpc1_1 gpc8205 (
      {stage1_49[212]},
      {stage2_49[86]}
   );
   gpc1_1 gpc8206 (
      {stage1_49[213]},
      {stage2_49[87]}
   );
   gpc1_1 gpc8207 (
      {stage1_49[214]},
      {stage2_49[88]}
   );
   gpc1_1 gpc8208 (
      {stage1_49[215]},
      {stage2_49[89]}
   );
   gpc1_1 gpc8209 (
      {stage1_49[216]},
      {stage2_49[90]}
   );
   gpc1_1 gpc8210 (
      {stage1_49[217]},
      {stage2_49[91]}
   );
   gpc1_1 gpc8211 (
      {stage1_49[218]},
      {stage2_49[92]}
   );
   gpc1_1 gpc8212 (
      {stage1_49[219]},
      {stage2_49[93]}
   );
   gpc1_1 gpc8213 (
      {stage1_49[220]},
      {stage2_49[94]}
   );
   gpc1_1 gpc8214 (
      {stage1_49[221]},
      {stage2_49[95]}
   );
   gpc1_1 gpc8215 (
      {stage1_49[222]},
      {stage2_49[96]}
   );
   gpc1_1 gpc8216 (
      {stage1_49[223]},
      {stage2_49[97]}
   );
   gpc1_1 gpc8217 (
      {stage1_49[224]},
      {stage2_49[98]}
   );
   gpc1_1 gpc8218 (
      {stage1_49[225]},
      {stage2_49[99]}
   );
   gpc1_1 gpc8219 (
      {stage1_49[226]},
      {stage2_49[100]}
   );
   gpc1_1 gpc8220 (
      {stage1_49[227]},
      {stage2_49[101]}
   );
   gpc1_1 gpc8221 (
      {stage1_49[228]},
      {stage2_49[102]}
   );
   gpc1_1 gpc8222 (
      {stage1_49[229]},
      {stage2_49[103]}
   );
   gpc1_1 gpc8223 (
      {stage1_49[230]},
      {stage2_49[104]}
   );
   gpc1_1 gpc8224 (
      {stage1_49[231]},
      {stage2_49[105]}
   );
   gpc1_1 gpc8225 (
      {stage1_49[232]},
      {stage2_49[106]}
   );
   gpc1_1 gpc8226 (
      {stage1_49[233]},
      {stage2_49[107]}
   );
   gpc1_1 gpc8227 (
      {stage1_49[234]},
      {stage2_49[108]}
   );
   gpc1_1 gpc8228 (
      {stage1_49[235]},
      {stage2_49[109]}
   );
   gpc1_1 gpc8229 (
      {stage1_49[236]},
      {stage2_49[110]}
   );
   gpc1_1 gpc8230 (
      {stage1_49[237]},
      {stage2_49[111]}
   );
   gpc1_1 gpc8231 (
      {stage1_49[238]},
      {stage2_49[112]}
   );
   gpc1_1 gpc8232 (
      {stage1_49[239]},
      {stage2_49[113]}
   );
   gpc1_1 gpc8233 (
      {stage1_49[240]},
      {stage2_49[114]}
   );
   gpc1_1 gpc8234 (
      {stage1_49[241]},
      {stage2_49[115]}
   );
   gpc1_1 gpc8235 (
      {stage1_50[134]},
      {stage2_50[70]}
   );
   gpc1_1 gpc8236 (
      {stage1_50[135]},
      {stage2_50[71]}
   );
   gpc1_1 gpc8237 (
      {stage1_50[136]},
      {stage2_50[72]}
   );
   gpc1_1 gpc8238 (
      {stage1_50[137]},
      {stage2_50[73]}
   );
   gpc1_1 gpc8239 (
      {stage1_50[138]},
      {stage2_50[74]}
   );
   gpc1_1 gpc8240 (
      {stage1_50[139]},
      {stage2_50[75]}
   );
   gpc1_1 gpc8241 (
      {stage1_50[140]},
      {stage2_50[76]}
   );
   gpc1_1 gpc8242 (
      {stage1_50[141]},
      {stage2_50[77]}
   );
   gpc1_1 gpc8243 (
      {stage1_50[142]},
      {stage2_50[78]}
   );
   gpc1_1 gpc8244 (
      {stage1_50[143]},
      {stage2_50[79]}
   );
   gpc1_1 gpc8245 (
      {stage1_50[144]},
      {stage2_50[80]}
   );
   gpc1_1 gpc8246 (
      {stage1_50[145]},
      {stage2_50[81]}
   );
   gpc1_1 gpc8247 (
      {stage1_50[146]},
      {stage2_50[82]}
   );
   gpc1_1 gpc8248 (
      {stage1_50[147]},
      {stage2_50[83]}
   );
   gpc1_1 gpc8249 (
      {stage1_50[148]},
      {stage2_50[84]}
   );
   gpc1_1 gpc8250 (
      {stage1_50[149]},
      {stage2_50[85]}
   );
   gpc1_1 gpc8251 (
      {stage1_50[150]},
      {stage2_50[86]}
   );
   gpc1_1 gpc8252 (
      {stage1_50[151]},
      {stage2_50[87]}
   );
   gpc1_1 gpc8253 (
      {stage1_50[152]},
      {stage2_50[88]}
   );
   gpc1_1 gpc8254 (
      {stage1_50[153]},
      {stage2_50[89]}
   );
   gpc1_1 gpc8255 (
      {stage1_50[154]},
      {stage2_50[90]}
   );
   gpc1_1 gpc8256 (
      {stage1_50[155]},
      {stage2_50[91]}
   );
   gpc1_1 gpc8257 (
      {stage1_50[156]},
      {stage2_50[92]}
   );
   gpc1_1 gpc8258 (
      {stage1_50[157]},
      {stage2_50[93]}
   );
   gpc1_1 gpc8259 (
      {stage1_50[158]},
      {stage2_50[94]}
   );
   gpc1_1 gpc8260 (
      {stage1_50[159]},
      {stage2_50[95]}
   );
   gpc1_1 gpc8261 (
      {stage1_50[160]},
      {stage2_50[96]}
   );
   gpc1_1 gpc8262 (
      {stage1_50[161]},
      {stage2_50[97]}
   );
   gpc1_1 gpc8263 (
      {stage1_50[162]},
      {stage2_50[98]}
   );
   gpc1_1 gpc8264 (
      {stage1_50[163]},
      {stage2_50[99]}
   );
   gpc1_1 gpc8265 (
      {stage1_50[164]},
      {stage2_50[100]}
   );
   gpc1_1 gpc8266 (
      {stage1_50[165]},
      {stage2_50[101]}
   );
   gpc1_1 gpc8267 (
      {stage1_50[166]},
      {stage2_50[102]}
   );
   gpc1_1 gpc8268 (
      {stage1_50[167]},
      {stage2_50[103]}
   );
   gpc1_1 gpc8269 (
      {stage1_50[168]},
      {stage2_50[104]}
   );
   gpc1_1 gpc8270 (
      {stage1_50[169]},
      {stage2_50[105]}
   );
   gpc1_1 gpc8271 (
      {stage1_50[170]},
      {stage2_50[106]}
   );
   gpc1_1 gpc8272 (
      {stage1_50[171]},
      {stage2_50[107]}
   );
   gpc1_1 gpc8273 (
      {stage1_50[172]},
      {stage2_50[108]}
   );
   gpc1_1 gpc8274 (
      {stage1_50[173]},
      {stage2_50[109]}
   );
   gpc1_1 gpc8275 (
      {stage1_50[174]},
      {stage2_50[110]}
   );
   gpc1_1 gpc8276 (
      {stage1_50[175]},
      {stage2_50[111]}
   );
   gpc1_1 gpc8277 (
      {stage1_50[176]},
      {stage2_50[112]}
   );
   gpc1_1 gpc8278 (
      {stage1_50[177]},
      {stage2_50[113]}
   );
   gpc1_1 gpc8279 (
      {stage1_50[178]},
      {stage2_50[114]}
   );
   gpc1_1 gpc8280 (
      {stage1_50[179]},
      {stage2_50[115]}
   );
   gpc1_1 gpc8281 (
      {stage1_50[180]},
      {stage2_50[116]}
   );
   gpc1_1 gpc8282 (
      {stage1_50[181]},
      {stage2_50[117]}
   );
   gpc1_1 gpc8283 (
      {stage1_50[182]},
      {stage2_50[118]}
   );
   gpc1_1 gpc8284 (
      {stage1_50[183]},
      {stage2_50[119]}
   );
   gpc1_1 gpc8285 (
      {stage1_50[184]},
      {stage2_50[120]}
   );
   gpc1_1 gpc8286 (
      {stage1_50[185]},
      {stage2_50[121]}
   );
   gpc1_1 gpc8287 (
      {stage1_50[186]},
      {stage2_50[122]}
   );
   gpc1_1 gpc8288 (
      {stage1_50[187]},
      {stage2_50[123]}
   );
   gpc1_1 gpc8289 (
      {stage1_50[188]},
      {stage2_50[124]}
   );
   gpc1_1 gpc8290 (
      {stage1_50[189]},
      {stage2_50[125]}
   );
   gpc1_1 gpc8291 (
      {stage1_50[190]},
      {stage2_50[126]}
   );
   gpc1_1 gpc8292 (
      {stage1_50[191]},
      {stage2_50[127]}
   );
   gpc1_1 gpc8293 (
      {stage1_50[192]},
      {stage2_50[128]}
   );
   gpc1_1 gpc8294 (
      {stage1_50[193]},
      {stage2_50[129]}
   );
   gpc1_1 gpc8295 (
      {stage1_50[194]},
      {stage2_50[130]}
   );
   gpc1_1 gpc8296 (
      {stage1_50[195]},
      {stage2_50[131]}
   );
   gpc1_1 gpc8297 (
      {stage1_50[196]},
      {stage2_50[132]}
   );
   gpc1_1 gpc8298 (
      {stage1_50[197]},
      {stage2_50[133]}
   );
   gpc1_1 gpc8299 (
      {stage1_50[198]},
      {stage2_50[134]}
   );
   gpc1_1 gpc8300 (
      {stage1_50[199]},
      {stage2_50[135]}
   );
   gpc1_1 gpc8301 (
      {stage1_50[200]},
      {stage2_50[136]}
   );
   gpc1_1 gpc8302 (
      {stage1_50[201]},
      {stage2_50[137]}
   );
   gpc1_1 gpc8303 (
      {stage1_50[202]},
      {stage2_50[138]}
   );
   gpc1_1 gpc8304 (
      {stage1_50[203]},
      {stage2_50[139]}
   );
   gpc1_1 gpc8305 (
      {stage1_50[204]},
      {stage2_50[140]}
   );
   gpc1_1 gpc8306 (
      {stage1_50[205]},
      {stage2_50[141]}
   );
   gpc1_1 gpc8307 (
      {stage1_50[206]},
      {stage2_50[142]}
   );
   gpc1_1 gpc8308 (
      {stage1_50[207]},
      {stage2_50[143]}
   );
   gpc1_1 gpc8309 (
      {stage1_50[208]},
      {stage2_50[144]}
   );
   gpc1_1 gpc8310 (
      {stage1_50[209]},
      {stage2_50[145]}
   );
   gpc1_1 gpc8311 (
      {stage1_50[210]},
      {stage2_50[146]}
   );
   gpc1_1 gpc8312 (
      {stage1_50[211]},
      {stage2_50[147]}
   );
   gpc1_1 gpc8313 (
      {stage1_50[212]},
      {stage2_50[148]}
   );
   gpc1_1 gpc8314 (
      {stage1_50[213]},
      {stage2_50[149]}
   );
   gpc1_1 gpc8315 (
      {stage1_50[214]},
      {stage2_50[150]}
   );
   gpc1_1 gpc8316 (
      {stage1_50[215]},
      {stage2_50[151]}
   );
   gpc1_1 gpc8317 (
      {stage1_50[216]},
      {stage2_50[152]}
   );
   gpc1_1 gpc8318 (
      {stage1_51[224]},
      {stage2_51[85]}
   );
   gpc1_1 gpc8319 (
      {stage1_51[225]},
      {stage2_51[86]}
   );
   gpc1_1 gpc8320 (
      {stage1_51[226]},
      {stage2_51[87]}
   );
   gpc1_1 gpc8321 (
      {stage1_52[269]},
      {stage2_52[93]}
   );
   gpc1_1 gpc8322 (
      {stage1_52[270]},
      {stage2_52[94]}
   );
   gpc1_1 gpc8323 (
      {stage1_52[271]},
      {stage2_52[95]}
   );
   gpc1_1 gpc8324 (
      {stage1_52[272]},
      {stage2_52[96]}
   );
   gpc1_1 gpc8325 (
      {stage1_52[273]},
      {stage2_52[97]}
   );
   gpc1_1 gpc8326 (
      {stage1_52[274]},
      {stage2_52[98]}
   );
   gpc1_1 gpc8327 (
      {stage1_52[275]},
      {stage2_52[99]}
   );
   gpc1_1 gpc8328 (
      {stage1_52[276]},
      {stage2_52[100]}
   );
   gpc1_1 gpc8329 (
      {stage1_52[277]},
      {stage2_52[101]}
   );
   gpc1_1 gpc8330 (
      {stage1_52[278]},
      {stage2_52[102]}
   );
   gpc1_1 gpc8331 (
      {stage1_52[279]},
      {stage2_52[103]}
   );
   gpc1_1 gpc8332 (
      {stage1_52[280]},
      {stage2_52[104]}
   );
   gpc1_1 gpc8333 (
      {stage1_52[281]},
      {stage2_52[105]}
   );
   gpc1_1 gpc8334 (
      {stage1_52[282]},
      {stage2_52[106]}
   );
   gpc1_1 gpc8335 (
      {stage1_52[283]},
      {stage2_52[107]}
   );
   gpc1_1 gpc8336 (
      {stage1_52[284]},
      {stage2_52[108]}
   );
   gpc1_1 gpc8337 (
      {stage1_52[285]},
      {stage2_52[109]}
   );
   gpc1_1 gpc8338 (
      {stage1_52[286]},
      {stage2_52[110]}
   );
   gpc1_1 gpc8339 (
      {stage1_52[287]},
      {stage2_52[111]}
   );
   gpc1_1 gpc8340 (
      {stage1_52[288]},
      {stage2_52[112]}
   );
   gpc1_1 gpc8341 (
      {stage1_52[289]},
      {stage2_52[113]}
   );
   gpc1_1 gpc8342 (
      {stage1_52[290]},
      {stage2_52[114]}
   );
   gpc1_1 gpc8343 (
      {stage1_52[291]},
      {stage2_52[115]}
   );
   gpc1_1 gpc8344 (
      {stage1_52[292]},
      {stage2_52[116]}
   );
   gpc1_1 gpc8345 (
      {stage1_52[293]},
      {stage2_52[117]}
   );
   gpc1_1 gpc8346 (
      {stage1_52[294]},
      {stage2_52[118]}
   );
   gpc1_1 gpc8347 (
      {stage1_52[295]},
      {stage2_52[119]}
   );
   gpc1_1 gpc8348 (
      {stage1_52[296]},
      {stage2_52[120]}
   );
   gpc1_1 gpc8349 (
      {stage1_52[297]},
      {stage2_52[121]}
   );
   gpc1_1 gpc8350 (
      {stage1_52[298]},
      {stage2_52[122]}
   );
   gpc1_1 gpc8351 (
      {stage1_52[299]},
      {stage2_52[123]}
   );
   gpc1_1 gpc8352 (
      {stage1_52[300]},
      {stage2_52[124]}
   );
   gpc1_1 gpc8353 (
      {stage1_52[301]},
      {stage2_52[125]}
   );
   gpc1_1 gpc8354 (
      {stage1_52[302]},
      {stage2_52[126]}
   );
   gpc1_1 gpc8355 (
      {stage1_52[303]},
      {stage2_52[127]}
   );
   gpc1_1 gpc8356 (
      {stage1_53[173]},
      {stage2_53[83]}
   );
   gpc1_1 gpc8357 (
      {stage1_53[174]},
      {stage2_53[84]}
   );
   gpc1_1 gpc8358 (
      {stage1_53[175]},
      {stage2_53[85]}
   );
   gpc1_1 gpc8359 (
      {stage1_53[176]},
      {stage2_53[86]}
   );
   gpc1_1 gpc8360 (
      {stage1_53[177]},
      {stage2_53[87]}
   );
   gpc1_1 gpc8361 (
      {stage1_53[178]},
      {stage2_53[88]}
   );
   gpc1_1 gpc8362 (
      {stage1_53[179]},
      {stage2_53[89]}
   );
   gpc1_1 gpc8363 (
      {stage1_53[180]},
      {stage2_53[90]}
   );
   gpc1_1 gpc8364 (
      {stage1_53[181]},
      {stage2_53[91]}
   );
   gpc1_1 gpc8365 (
      {stage1_53[182]},
      {stage2_53[92]}
   );
   gpc1_1 gpc8366 (
      {stage1_53[183]},
      {stage2_53[93]}
   );
   gpc1_1 gpc8367 (
      {stage1_53[184]},
      {stage2_53[94]}
   );
   gpc1_1 gpc8368 (
      {stage1_53[185]},
      {stage2_53[95]}
   );
   gpc1_1 gpc8369 (
      {stage1_53[186]},
      {stage2_53[96]}
   );
   gpc1_1 gpc8370 (
      {stage1_54[216]},
      {stage2_54[77]}
   );
   gpc1_1 gpc8371 (
      {stage1_54[217]},
      {stage2_54[78]}
   );
   gpc1_1 gpc8372 (
      {stage1_54[218]},
      {stage2_54[79]}
   );
   gpc1_1 gpc8373 (
      {stage1_54[219]},
      {stage2_54[80]}
   );
   gpc1_1 gpc8374 (
      {stage1_54[220]},
      {stage2_54[81]}
   );
   gpc1_1 gpc8375 (
      {stage1_54[221]},
      {stage2_54[82]}
   );
   gpc1_1 gpc8376 (
      {stage1_54[222]},
      {stage2_54[83]}
   );
   gpc1_1 gpc8377 (
      {stage1_54[223]},
      {stage2_54[84]}
   );
   gpc1_1 gpc8378 (
      {stage1_54[224]},
      {stage2_54[85]}
   );
   gpc1_1 gpc8379 (
      {stage1_54[225]},
      {stage2_54[86]}
   );
   gpc1_1 gpc8380 (
      {stage1_54[226]},
      {stage2_54[87]}
   );
   gpc1_1 gpc8381 (
      {stage1_54[227]},
      {stage2_54[88]}
   );
   gpc1_1 gpc8382 (
      {stage1_54[228]},
      {stage2_54[89]}
   );
   gpc1_1 gpc8383 (
      {stage1_54[229]},
      {stage2_54[90]}
   );
   gpc1_1 gpc8384 (
      {stage1_54[230]},
      {stage2_54[91]}
   );
   gpc1_1 gpc8385 (
      {stage1_54[231]},
      {stage2_54[92]}
   );
   gpc1_1 gpc8386 (
      {stage1_54[232]},
      {stage2_54[93]}
   );
   gpc1_1 gpc8387 (
      {stage1_54[233]},
      {stage2_54[94]}
   );
   gpc1_1 gpc8388 (
      {stage1_54[234]},
      {stage2_54[95]}
   );
   gpc1_1 gpc8389 (
      {stage1_54[235]},
      {stage2_54[96]}
   );
   gpc1_1 gpc8390 (
      {stage1_54[236]},
      {stage2_54[97]}
   );
   gpc1_1 gpc8391 (
      {stage1_54[237]},
      {stage2_54[98]}
   );
   gpc1_1 gpc8392 (
      {stage1_54[238]},
      {stage2_54[99]}
   );
   gpc1_1 gpc8393 (
      {stage1_54[239]},
      {stage2_54[100]}
   );
   gpc1_1 gpc8394 (
      {stage1_54[240]},
      {stage2_54[101]}
   );
   gpc1_1 gpc8395 (
      {stage1_54[241]},
      {stage2_54[102]}
   );
   gpc1_1 gpc8396 (
      {stage1_54[242]},
      {stage2_54[103]}
   );
   gpc1_1 gpc8397 (
      {stage1_54[243]},
      {stage2_54[104]}
   );
   gpc1_1 gpc8398 (
      {stage1_54[244]},
      {stage2_54[105]}
   );
   gpc1_1 gpc8399 (
      {stage1_54[245]},
      {stage2_54[106]}
   );
   gpc1_1 gpc8400 (
      {stage1_54[246]},
      {stage2_54[107]}
   );
   gpc1_1 gpc8401 (
      {stage1_54[247]},
      {stage2_54[108]}
   );
   gpc1_1 gpc8402 (
      {stage1_54[248]},
      {stage2_54[109]}
   );
   gpc1_1 gpc8403 (
      {stage1_54[249]},
      {stage2_54[110]}
   );
   gpc1_1 gpc8404 (
      {stage1_54[250]},
      {stage2_54[111]}
   );
   gpc1_1 gpc8405 (
      {stage1_54[251]},
      {stage2_54[112]}
   );
   gpc1_1 gpc8406 (
      {stage1_54[252]},
      {stage2_54[113]}
   );
   gpc1_1 gpc8407 (
      {stage1_54[253]},
      {stage2_54[114]}
   );
   gpc1_1 gpc8408 (
      {stage1_54[254]},
      {stage2_54[115]}
   );
   gpc1_1 gpc8409 (
      {stage1_54[255]},
      {stage2_54[116]}
   );
   gpc1_1 gpc8410 (
      {stage1_54[256]},
      {stage2_54[117]}
   );
   gpc1_1 gpc8411 (
      {stage1_54[257]},
      {stage2_54[118]}
   );
   gpc1_1 gpc8412 (
      {stage1_54[258]},
      {stage2_54[119]}
   );
   gpc1_1 gpc8413 (
      {stage1_54[259]},
      {stage2_54[120]}
   );
   gpc1_1 gpc8414 (
      {stage1_54[260]},
      {stage2_54[121]}
   );
   gpc1_1 gpc8415 (
      {stage1_54[261]},
      {stage2_54[122]}
   );
   gpc1_1 gpc8416 (
      {stage1_54[262]},
      {stage2_54[123]}
   );
   gpc1_1 gpc8417 (
      {stage1_55[219]},
      {stage2_55[104]}
   );
   gpc1_1 gpc8418 (
      {stage1_55[220]},
      {stage2_55[105]}
   );
   gpc1_1 gpc8419 (
      {stage1_55[221]},
      {stage2_55[106]}
   );
   gpc1_1 gpc8420 (
      {stage1_55[222]},
      {stage2_55[107]}
   );
   gpc1_1 gpc8421 (
      {stage1_55[223]},
      {stage2_55[108]}
   );
   gpc1_1 gpc8422 (
      {stage1_55[224]},
      {stage2_55[109]}
   );
   gpc1_1 gpc8423 (
      {stage1_55[225]},
      {stage2_55[110]}
   );
   gpc1_1 gpc8424 (
      {stage1_56[225]},
      {stage2_56[100]}
   );
   gpc1_1 gpc8425 (
      {stage1_56[226]},
      {stage2_56[101]}
   );
   gpc1_1 gpc8426 (
      {stage1_56[227]},
      {stage2_56[102]}
   );
   gpc1_1 gpc8427 (
      {stage1_56[228]},
      {stage2_56[103]}
   );
   gpc1_1 gpc8428 (
      {stage1_56[229]},
      {stage2_56[104]}
   );
   gpc1_1 gpc8429 (
      {stage1_56[230]},
      {stage2_56[105]}
   );
   gpc1_1 gpc8430 (
      {stage1_56[231]},
      {stage2_56[106]}
   );
   gpc1_1 gpc8431 (
      {stage1_56[232]},
      {stage2_56[107]}
   );
   gpc1_1 gpc8432 (
      {stage1_56[233]},
      {stage2_56[108]}
   );
   gpc1_1 gpc8433 (
      {stage1_56[234]},
      {stage2_56[109]}
   );
   gpc1_1 gpc8434 (
      {stage1_56[235]},
      {stage2_56[110]}
   );
   gpc1_1 gpc8435 (
      {stage1_56[236]},
      {stage2_56[111]}
   );
   gpc1_1 gpc8436 (
      {stage1_56[237]},
      {stage2_56[112]}
   );
   gpc1_1 gpc8437 (
      {stage1_56[238]},
      {stage2_56[113]}
   );
   gpc1_1 gpc8438 (
      {stage1_56[239]},
      {stage2_56[114]}
   );
   gpc1_1 gpc8439 (
      {stage1_56[240]},
      {stage2_56[115]}
   );
   gpc1_1 gpc8440 (
      {stage1_56[241]},
      {stage2_56[116]}
   );
   gpc1_1 gpc8441 (
      {stage1_56[242]},
      {stage2_56[117]}
   );
   gpc1_1 gpc8442 (
      {stage1_56[243]},
      {stage2_56[118]}
   );
   gpc1_1 gpc8443 (
      {stage1_56[244]},
      {stage2_56[119]}
   );
   gpc1_1 gpc8444 (
      {stage1_56[245]},
      {stage2_56[120]}
   );
   gpc1_1 gpc8445 (
      {stage1_56[246]},
      {stage2_56[121]}
   );
   gpc1_1 gpc8446 (
      {stage1_56[247]},
      {stage2_56[122]}
   );
   gpc1_1 gpc8447 (
      {stage1_56[248]},
      {stage2_56[123]}
   );
   gpc1_1 gpc8448 (
      {stage1_56[249]},
      {stage2_56[124]}
   );
   gpc1_1 gpc8449 (
      {stage1_56[250]},
      {stage2_56[125]}
   );
   gpc1_1 gpc8450 (
      {stage1_56[251]},
      {stage2_56[126]}
   );
   gpc1_1 gpc8451 (
      {stage1_56[252]},
      {stage2_56[127]}
   );
   gpc1_1 gpc8452 (
      {stage1_56[253]},
      {stage2_56[128]}
   );
   gpc1_1 gpc8453 (
      {stage1_56[254]},
      {stage2_56[129]}
   );
   gpc1_1 gpc8454 (
      {stage1_56[255]},
      {stage2_56[130]}
   );
   gpc1_1 gpc8455 (
      {stage1_56[256]},
      {stage2_56[131]}
   );
   gpc1_1 gpc8456 (
      {stage1_59[268]},
      {stage2_59[114]}
   );
   gpc1_1 gpc8457 (
      {stage1_59[269]},
      {stage2_59[115]}
   );
   gpc1_1 gpc8458 (
      {stage1_59[270]},
      {stage2_59[116]}
   );
   gpc1_1 gpc8459 (
      {stage1_59[271]},
      {stage2_59[117]}
   );
   gpc1_1 gpc8460 (
      {stage1_59[272]},
      {stage2_59[118]}
   );
   gpc1_1 gpc8461 (
      {stage1_59[273]},
      {stage2_59[119]}
   );
   gpc1_1 gpc8462 (
      {stage1_59[274]},
      {stage2_59[120]}
   );
   gpc1_1 gpc8463 (
      {stage1_59[275]},
      {stage2_59[121]}
   );
   gpc1_1 gpc8464 (
      {stage1_59[276]},
      {stage2_59[122]}
   );
   gpc1_1 gpc8465 (
      {stage1_59[277]},
      {stage2_59[123]}
   );
   gpc1_1 gpc8466 (
      {stage1_59[278]},
      {stage2_59[124]}
   );
   gpc1_1 gpc8467 (
      {stage1_59[279]},
      {stage2_59[125]}
   );
   gpc1_1 gpc8468 (
      {stage1_59[280]},
      {stage2_59[126]}
   );
   gpc1_1 gpc8469 (
      {stage1_59[281]},
      {stage2_59[127]}
   );
   gpc1_1 gpc8470 (
      {stage1_59[282]},
      {stage2_59[128]}
   );
   gpc1_1 gpc8471 (
      {stage1_59[283]},
      {stage2_59[129]}
   );
   gpc1_1 gpc8472 (
      {stage1_59[284]},
      {stage2_59[130]}
   );
   gpc1_1 gpc8473 (
      {stage1_59[285]},
      {stage2_59[131]}
   );
   gpc1_1 gpc8474 (
      {stage1_59[286]},
      {stage2_59[132]}
   );
   gpc1_1 gpc8475 (
      {stage1_59[287]},
      {stage2_59[133]}
   );
   gpc1_1 gpc8476 (
      {stage1_59[288]},
      {stage2_59[134]}
   );
   gpc1_1 gpc8477 (
      {stage1_59[289]},
      {stage2_59[135]}
   );
   gpc1_1 gpc8478 (
      {stage1_59[290]},
      {stage2_59[136]}
   );
   gpc1_1 gpc8479 (
      {stage1_59[291]},
      {stage2_59[137]}
   );
   gpc1_1 gpc8480 (
      {stage1_59[292]},
      {stage2_59[138]}
   );
   gpc1_1 gpc8481 (
      {stage1_59[293]},
      {stage2_59[139]}
   );
   gpc1_1 gpc8482 (
      {stage1_60[190]},
      {stage2_60[101]}
   );
   gpc1_1 gpc8483 (
      {stage1_60[191]},
      {stage2_60[102]}
   );
   gpc1_1 gpc8484 (
      {stage1_60[192]},
      {stage2_60[103]}
   );
   gpc1_1 gpc8485 (
      {stage1_60[193]},
      {stage2_60[104]}
   );
   gpc1_1 gpc8486 (
      {stage1_60[194]},
      {stage2_60[105]}
   );
   gpc1_1 gpc8487 (
      {stage1_60[195]},
      {stage2_60[106]}
   );
   gpc1_1 gpc8488 (
      {stage1_60[196]},
      {stage2_60[107]}
   );
   gpc1_1 gpc8489 (
      {stage1_60[197]},
      {stage2_60[108]}
   );
   gpc1_1 gpc8490 (
      {stage1_60[198]},
      {stage2_60[109]}
   );
   gpc1_1 gpc8491 (
      {stage1_60[199]},
      {stage2_60[110]}
   );
   gpc1_1 gpc8492 (
      {stage1_61[198]},
      {stage2_61[83]}
   );
   gpc1_1 gpc8493 (
      {stage1_61[199]},
      {stage2_61[84]}
   );
   gpc1_1 gpc8494 (
      {stage1_61[200]},
      {stage2_61[85]}
   );
   gpc1_1 gpc8495 (
      {stage1_61[201]},
      {stage2_61[86]}
   );
   gpc1_1 gpc8496 (
      {stage1_61[202]},
      {stage2_61[87]}
   );
   gpc1_1 gpc8497 (
      {stage1_61[203]},
      {stage2_61[88]}
   );
   gpc1_1 gpc8498 (
      {stage1_61[204]},
      {stage2_61[89]}
   );
   gpc1_1 gpc8499 (
      {stage1_61[205]},
      {stage2_61[90]}
   );
   gpc1_1 gpc8500 (
      {stage1_61[206]},
      {stage2_61[91]}
   );
   gpc1_1 gpc8501 (
      {stage1_61[207]},
      {stage2_61[92]}
   );
   gpc1_1 gpc8502 (
      {stage1_61[208]},
      {stage2_61[93]}
   );
   gpc1_1 gpc8503 (
      {stage1_61[209]},
      {stage2_61[94]}
   );
   gpc1_1 gpc8504 (
      {stage1_61[210]},
      {stage2_61[95]}
   );
   gpc1_1 gpc8505 (
      {stage1_61[211]},
      {stage2_61[96]}
   );
   gpc1_1 gpc8506 (
      {stage1_61[212]},
      {stage2_61[97]}
   );
   gpc1_1 gpc8507 (
      {stage1_61[213]},
      {stage2_61[98]}
   );
   gpc1_1 gpc8508 (
      {stage1_61[214]},
      {stage2_61[99]}
   );
   gpc1_1 gpc8509 (
      {stage1_61[215]},
      {stage2_61[100]}
   );
   gpc1_1 gpc8510 (
      {stage1_61[216]},
      {stage2_61[101]}
   );
   gpc1_1 gpc8511 (
      {stage1_62[346]},
      {stage2_62[118]}
   );
   gpc1_1 gpc8512 (
      {stage1_62[347]},
      {stage2_62[119]}
   );
   gpc1_1 gpc8513 (
      {stage1_62[348]},
      {stage2_62[120]}
   );
   gpc1_1 gpc8514 (
      {stage1_62[349]},
      {stage2_62[121]}
   );
   gpc1_1 gpc8515 (
      {stage1_62[350]},
      {stage2_62[122]}
   );
   gpc1_1 gpc8516 (
      {stage1_62[351]},
      {stage2_62[123]}
   );
   gpc1_1 gpc8517 (
      {stage1_62[352]},
      {stage2_62[124]}
   );
   gpc1_1 gpc8518 (
      {stage1_62[353]},
      {stage2_62[125]}
   );
   gpc1_1 gpc8519 (
      {stage1_62[354]},
      {stage2_62[126]}
   );
   gpc1_1 gpc8520 (
      {stage1_62[355]},
      {stage2_62[127]}
   );
   gpc1_1 gpc8521 (
      {stage1_62[356]},
      {stage2_62[128]}
   );
   gpc1_1 gpc8522 (
      {stage1_62[357]},
      {stage2_62[129]}
   );
   gpc1_1 gpc8523 (
      {stage1_62[358]},
      {stage2_62[130]}
   );
   gpc1_1 gpc8524 (
      {stage1_62[359]},
      {stage2_62[131]}
   );
   gpc1_1 gpc8525 (
      {stage1_62[360]},
      {stage2_62[132]}
   );
   gpc1_1 gpc8526 (
      {stage1_62[361]},
      {stage2_62[133]}
   );
   gpc1_1 gpc8527 (
      {stage1_62[362]},
      {stage2_62[134]}
   );
   gpc1_1 gpc8528 (
      {stage1_62[363]},
      {stage2_62[135]}
   );
   gpc1_1 gpc8529 (
      {stage1_62[364]},
      {stage2_62[136]}
   );
   gpc1_1 gpc8530 (
      {stage1_62[365]},
      {stage2_62[137]}
   );
   gpc1_1 gpc8531 (
      {stage1_62[366]},
      {stage2_62[138]}
   );
   gpc1_1 gpc8532 (
      {stage1_62[367]},
      {stage2_62[139]}
   );
   gpc1_1 gpc8533 (
      {stage1_62[368]},
      {stage2_62[140]}
   );
   gpc1_1 gpc8534 (
      {stage1_62[369]},
      {stage2_62[141]}
   );
   gpc1_1 gpc8535 (
      {stage1_62[370]},
      {stage2_62[142]}
   );
   gpc1_1 gpc8536 (
      {stage1_62[371]},
      {stage2_62[143]}
   );
   gpc1_1 gpc8537 (
      {stage1_62[372]},
      {stage2_62[144]}
   );
   gpc1_1 gpc8538 (
      {stage1_64[94]},
      {stage2_64[84]}
   );
   gpc1_1 gpc8539 (
      {stage1_64[95]},
      {stage2_64[85]}
   );
   gpc1_1 gpc8540 (
      {stage1_64[96]},
      {stage2_64[86]}
   );
   gpc1_1 gpc8541 (
      {stage1_64[97]},
      {stage2_64[87]}
   );
   gpc1_1 gpc8542 (
      {stage1_64[98]},
      {stage2_64[88]}
   );
   gpc1_1 gpc8543 (
      {stage1_64[99]},
      {stage2_64[89]}
   );
   gpc1_1 gpc8544 (
      {stage1_64[100]},
      {stage2_64[90]}
   );
   gpc1_1 gpc8545 (
      {stage1_64[101]},
      {stage2_64[91]}
   );
   gpc1_1 gpc8546 (
      {stage1_64[102]},
      {stage2_64[92]}
   );
   gpc1_1 gpc8547 (
      {stage1_64[103]},
      {stage2_64[93]}
   );
   gpc1_1 gpc8548 (
      {stage1_64[104]},
      {stage2_64[94]}
   );
   gpc1_1 gpc8549 (
      {stage1_64[105]},
      {stage2_64[95]}
   );
   gpc1_1 gpc8550 (
      {stage1_64[106]},
      {stage2_64[96]}
   );
   gpc1_1 gpc8551 (
      {stage1_64[107]},
      {stage2_64[97]}
   );
   gpc1_1 gpc8552 (
      {stage1_64[108]},
      {stage2_64[98]}
   );
   gpc1_1 gpc8553 (
      {stage1_64[109]},
      {stage2_64[99]}
   );
   gpc1_1 gpc8554 (
      {stage1_64[110]},
      {stage2_64[100]}
   );
   gpc1_1 gpc8555 (
      {stage1_64[111]},
      {stage2_64[101]}
   );
   gpc1_1 gpc8556 (
      {stage1_65[46]},
      {stage2_65[57]}
   );
   gpc1_1 gpc8557 (
      {stage1_65[47]},
      {stage2_65[58]}
   );
   gpc1_1 gpc8558 (
      {stage1_65[48]},
      {stage2_65[59]}
   );
   gpc1_1 gpc8559 (
      {stage1_65[49]},
      {stage2_65[60]}
   );
   gpc1_1 gpc8560 (
      {stage1_65[50]},
      {stage2_65[61]}
   );
   gpc1_1 gpc8561 (
      {stage1_65[51]},
      {stage2_65[62]}
   );
   gpc1_1 gpc8562 (
      {stage1_65[52]},
      {stage2_65[63]}
   );
   gpc1_1 gpc8563 (
      {stage1_65[53]},
      {stage2_65[64]}
   );
   gpc1_1 gpc8564 (
      {stage1_65[54]},
      {stage2_65[65]}
   );
   gpc1_1 gpc8565 (
      {stage1_65[55]},
      {stage2_65[66]}
   );
   gpc1_1 gpc8566 (
      {stage1_65[56]},
      {stage2_65[67]}
   );
   gpc1163_5 gpc8567 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc8568 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc8569 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[6]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc8570 (
      {stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18]},
      {stage2_1[7]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc615_5 gpc8571 (
      {stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_1[8]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc615_5 gpc8572 (
      {stage2_0[24], stage2_0[25], stage2_0[26], stage2_0[27], stage2_0[28]},
      {stage2_1[9]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1343_5 gpc8573 (
      {stage2_1[10], stage2_1[11], stage2_1[12]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[1], stage2_3[2], stage2_3[3]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc1343_5 gpc8574 (
      {stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[1]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc8575 (
      {stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc8576 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage3_6[0],stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9]}
   );
   gpc606_5 gpc8577 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49], stage2_2[50]},
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage3_6[1],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc8578 (
      {stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54], stage2_2[55], stage2_2[56]},
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage3_6[2],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc606_5 gpc8579 (
      {stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60], stage2_2[61], stage2_2[62]},
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage3_6[3],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc8580 (
      {stage2_2[63], stage2_2[64], stage2_2[65], stage2_2[66], stage2_2[67], stage2_2[68]},
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage3_6[4],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc8581 (
      {stage2_2[69], stage2_2[70], stage2_2[71], stage2_2[72], 1'b0, 1'b0},
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage3_6[5],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc207_4 gpc8582 (
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_5[0], stage2_5[1]},
      {stage3_6[6],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc207_4 gpc8583 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26]},
      {stage2_5[2], stage2_5[3]},
      {stage3_6[7],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc207_4 gpc8584 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_5[4], stage2_5[5]},
      {stage3_6[8],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc207_4 gpc8585 (
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40]},
      {stage2_5[6], stage2_5[7]},
      {stage3_6[9],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc207_4 gpc8586 (
      {stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[8], stage2_5[9]},
      {stage3_6[10],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc207_4 gpc8587 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_5[10], stage2_5[11]},
      {stage3_6[11],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc207_4 gpc8588 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_5[12], stage2_5[13]},
      {stage3_6[12],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc207_4 gpc8589 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_5[14], stage2_5[15]},
      {stage3_6[13],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc207_4 gpc8590 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75]},
      {stage2_5[16], stage2_5[17]},
      {stage3_6[14],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc207_4 gpc8591 (
      {stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_5[18], stage2_5[19]},
      {stage3_6[15],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc207_4 gpc8592 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_5[20], stage2_5[21]},
      {stage3_6[16],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc207_4 gpc8593 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96]},
      {stage2_5[22], stage2_5[23]},
      {stage3_6[17],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc207_4 gpc8594 (
      {stage2_3[97], stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103]},
      {stage2_5[24], stage2_5[25]},
      {stage3_6[18],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc207_4 gpc8595 (
      {stage2_3[104], stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109], stage2_3[110]},
      {stage2_5[26], stage2_5[27]},
      {stage3_6[19],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc207_4 gpc8596 (
      {stage2_3[111], stage2_3[112], stage2_3[113], stage2_3[114], stage2_3[115], stage2_3[116], stage2_3[117]},
      {stage2_5[28], stage2_5[29]},
      {stage3_6[20],stage3_5[23],stage3_4[29],stage3_3[29]}
   );
   gpc207_4 gpc8597 (
      {stage2_3[118], stage2_3[119], stage2_3[120], stage2_3[121], stage2_3[122], stage2_3[123], stage2_3[124]},
      {stage2_5[30], stage2_5[31]},
      {stage3_6[21],stage3_5[24],stage3_4[30],stage3_3[30]}
   );
   gpc207_4 gpc8598 (
      {stage2_3[125], stage2_3[126], stage2_3[127], stage2_3[128], stage2_3[129], stage2_3[130], stage2_3[131]},
      {stage2_5[32], stage2_5[33]},
      {stage3_6[22],stage3_5[25],stage3_4[31],stage3_3[31]}
   );
   gpc207_4 gpc8599 (
      {stage2_3[132], stage2_3[133], stage2_3[134], stage2_3[135], stage2_3[136], stage2_3[137], stage2_3[138]},
      {stage2_5[34], stage2_5[35]},
      {stage3_6[23],stage3_5[26],stage3_4[32],stage3_3[32]}
   );
   gpc207_4 gpc8600 (
      {stage2_3[139], stage2_3[140], stage2_3[141], stage2_3[142], stage2_3[143], stage2_3[144], stage2_3[145]},
      {stage2_5[36], stage2_5[37]},
      {stage3_6[24],stage3_5[27],stage3_4[33],stage3_3[33]}
   );
   gpc207_4 gpc8601 (
      {stage2_3[146], stage2_3[147], stage2_3[148], stage2_3[149], stage2_3[150], stage2_3[151], stage2_3[152]},
      {stage2_5[38], stage2_5[39]},
      {stage3_6[25],stage3_5[28],stage3_4[34],stage3_3[34]}
   );
   gpc207_4 gpc8602 (
      {stage2_3[153], stage2_3[154], stage2_3[155], stage2_3[156], stage2_3[157], stage2_3[158], stage2_3[159]},
      {stage2_5[40], stage2_5[41]},
      {stage3_6[26],stage3_5[29],stage3_4[35],stage3_3[35]}
   );
   gpc207_4 gpc8603 (
      {stage2_3[160], stage2_3[161], stage2_3[162], stage2_3[163], stage2_3[164], stage2_3[165], stage2_3[166]},
      {stage2_5[42], stage2_5[43]},
      {stage3_6[27],stage3_5[30],stage3_4[36],stage3_3[36]}
   );
   gpc207_4 gpc8604 (
      {stage2_3[167], stage2_3[168], stage2_3[169], stage2_3[170], stage2_3[171], stage2_3[172], stage2_3[173]},
      {stage2_5[44], stage2_5[45]},
      {stage3_6[28],stage3_5[31],stage3_4[37],stage3_3[37]}
   );
   gpc207_4 gpc8605 (
      {stage2_3[174], stage2_3[175], stage2_3[176], stage2_3[177], stage2_3[178], stage2_3[179], stage2_3[180]},
      {stage2_5[46], stage2_5[47]},
      {stage3_6[29],stage3_5[32],stage3_4[38],stage3_3[38]}
   );
   gpc207_4 gpc8606 (
      {stage2_3[181], stage2_3[182], stage2_3[183], stage2_3[184], stage2_3[185], stage2_3[186], stage2_3[187]},
      {stage2_5[48], stage2_5[49]},
      {stage3_6[30],stage3_5[33],stage3_4[39],stage3_3[39]}
   );
   gpc207_4 gpc8607 (
      {stage2_3[188], stage2_3[189], stage2_3[190], stage2_3[191], stage2_3[192], stage2_3[193], stage2_3[194]},
      {stage2_5[50], stage2_5[51]},
      {stage3_6[31],stage3_5[34],stage3_4[40],stage3_3[40]}
   );
   gpc207_4 gpc8608 (
      {stage2_3[195], stage2_3[196], stage2_3[197], stage2_3[198], stage2_3[199], stage2_3[200], stage2_3[201]},
      {stage2_5[52], stage2_5[53]},
      {stage3_6[32],stage3_5[35],stage3_4[41],stage3_3[41]}
   );
   gpc207_4 gpc8609 (
      {stage2_3[202], stage2_3[203], stage2_3[204], stage2_3[205], stage2_3[206], stage2_3[207], stage2_3[208]},
      {stage2_5[54], stage2_5[55]},
      {stage3_6[33],stage3_5[36],stage3_4[42],stage3_3[42]}
   );
   gpc207_4 gpc8610 (
      {stage2_3[209], stage2_3[210], stage2_3[211], stage2_3[212], stage2_3[213], stage2_3[214], stage2_3[215]},
      {stage2_5[56], stage2_5[57]},
      {stage3_6[34],stage3_5[37],stage3_4[43],stage3_3[43]}
   );
   gpc615_5 gpc8611 (
      {stage2_3[216], stage2_3[217], stage2_3[218], stage2_3[219], stage2_3[220]},
      {stage2_4[38]},
      {stage2_5[58], stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63]},
      {stage3_7[0],stage3_6[35],stage3_5[38],stage3_4[44],stage3_3[44]}
   );
   gpc615_5 gpc8612 (
      {stage2_3[221], stage2_3[222], stage2_3[223], stage2_3[224], stage2_3[225]},
      {stage2_4[39]},
      {stage2_5[64], stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage3_7[1],stage3_6[36],stage3_5[39],stage3_4[45],stage3_3[45]}
   );
   gpc615_5 gpc8613 (
      {stage2_3[226], stage2_3[227], stage2_3[228], stage2_3[229], stage2_3[230]},
      {stage2_4[40]},
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75]},
      {stage3_7[2],stage3_6[37],stage3_5[40],stage3_4[46],stage3_3[46]}
   );
   gpc615_5 gpc8614 (
      {stage2_3[231], stage2_3[232], stage2_3[233], stage2_3[234], stage2_3[235]},
      {stage2_4[41]},
      {stage2_5[76], stage2_5[77], stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81]},
      {stage3_7[3],stage3_6[38],stage3_5[41],stage3_4[47],stage3_3[47]}
   );
   gpc615_5 gpc8615 (
      {stage2_3[236], stage2_3[237], stage2_3[238], stage2_3[239], stage2_3[240]},
      {stage2_4[42]},
      {stage2_5[82], stage2_5[83], stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87]},
      {stage3_7[4],stage3_6[39],stage3_5[42],stage3_4[48],stage3_3[48]}
   );
   gpc615_5 gpc8616 (
      {stage2_3[241], stage2_3[242], stage2_3[243], stage2_3[244], stage2_3[245]},
      {stage2_4[43]},
      {stage2_5[88], stage2_5[89], stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93]},
      {stage3_7[5],stage3_6[40],stage3_5[43],stage3_4[49],stage3_3[49]}
   );
   gpc615_5 gpc8617 (
      {stage2_3[246], stage2_3[247], stage2_3[248], stage2_3[249], stage2_3[250]},
      {stage2_4[44]},
      {stage2_5[94], stage2_5[95], stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99]},
      {stage3_7[6],stage3_6[41],stage3_5[44],stage3_4[50],stage3_3[50]}
   );
   gpc615_5 gpc8618 (
      {stage2_3[251], stage2_3[252], stage2_3[253], 1'b0, 1'b0},
      {stage2_4[45]},
      {stage2_5[100], stage2_5[101], stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105]},
      {stage3_7[7],stage3_6[42],stage3_5[45],stage3_4[51],stage3_3[51]}
   );
   gpc606_5 gpc8619 (
      {stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[43],stage3_5[46],stage3_4[52]}
   );
   gpc606_5 gpc8620 (
      {stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[44],stage3_5[47],stage3_4[53]}
   );
   gpc606_5 gpc8621 (
      {stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[45],stage3_5[48],stage3_4[54]}
   );
   gpc606_5 gpc8622 (
      {stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[46],stage3_5[49],stage3_4[55]}
   );
   gpc606_5 gpc8623 (
      {stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[47],stage3_5[50],stage3_4[56]}
   );
   gpc606_5 gpc8624 (
      {stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[48],stage3_5[51],stage3_4[57]}
   );
   gpc606_5 gpc8625 (
      {stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[14],stage3_6[49],stage3_5[52],stage3_4[58]}
   );
   gpc606_5 gpc8626 (
      {stage2_4[88], stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], 1'b0},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[15],stage3_6[50],stage3_5[53],stage3_4[59]}
   );
   gpc606_5 gpc8627 (
      {stage2_5[106], stage2_5[107], stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[16],stage3_6[51],stage3_5[54]}
   );
   gpc615_5 gpc8628 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[9],stage3_7[17],stage3_6[52]}
   );
   gpc615_5 gpc8629 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[7]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[10],stage3_7[18],stage3_6[53]}
   );
   gpc615_5 gpc8630 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[8]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[11],stage3_7[19],stage3_6[54]}
   );
   gpc615_5 gpc8631 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[9]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[4],stage3_8[12],stage3_7[20],stage3_6[55]}
   );
   gpc615_5 gpc8632 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[10]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[5],stage3_8[13],stage3_7[21],stage3_6[56]}
   );
   gpc615_5 gpc8633 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[11]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[6],stage3_8[14],stage3_7[22],stage3_6[57]}
   );
   gpc615_5 gpc8634 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[12]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[7],stage3_8[15],stage3_7[23],stage3_6[58]}
   );
   gpc615_5 gpc8635 (
      {stage2_6[83], stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87]},
      {stage2_7[13]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[8],stage3_8[16],stage3_7[24],stage3_6[59]}
   );
   gpc615_5 gpc8636 (
      {stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91], stage2_6[92]},
      {stage2_7[14]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[9],stage3_8[17],stage3_7[25],stage3_6[60]}
   );
   gpc615_5 gpc8637 (
      {stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_7[15]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[10],stage3_8[18],stage3_7[26],stage3_6[61]}
   );
   gpc615_5 gpc8638 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102]},
      {stage2_7[16]},
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage3_10[10],stage3_9[11],stage3_8[19],stage3_7[27],stage3_6[62]}
   );
   gpc615_5 gpc8639 (
      {stage2_6[103], stage2_6[104], stage2_6[105], stage2_6[106], stage2_6[107]},
      {stage2_7[17]},
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage3_10[11],stage3_9[12],stage3_8[20],stage3_7[28],stage3_6[63]}
   );
   gpc615_5 gpc8640 (
      {stage2_6[108], stage2_6[109], stage2_6[110], stage2_6[111], stage2_6[112]},
      {stage2_7[18]},
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage3_10[12],stage3_9[13],stage3_8[21],stage3_7[29],stage3_6[64]}
   );
   gpc615_5 gpc8641 (
      {stage2_6[113], stage2_6[114], stage2_6[115], stage2_6[116], stage2_6[117]},
      {stage2_7[19]},
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage3_10[13],stage3_9[14],stage3_8[22],stage3_7[30],stage3_6[65]}
   );
   gpc615_5 gpc8642 (
      {stage2_6[118], stage2_6[119], stage2_6[120], 1'b0, 1'b0},
      {stage2_7[20]},
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage3_10[14],stage3_9[15],stage3_8[23],stage3_7[31],stage3_6[66]}
   );
   gpc2116_5 gpc8643 (
      {stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[90]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[15],stage3_9[16],stage3_8[24],stage3_7[32]}
   );
   gpc2116_5 gpc8644 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[91]},
      {stage2_9[1]},
      {stage2_10[2], stage2_10[3]},
      {stage3_11[1],stage3_10[16],stage3_9[17],stage3_8[25],stage3_7[33]}
   );
   gpc2116_5 gpc8645 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[92]},
      {stage2_9[2]},
      {stage2_10[4], stage2_10[5]},
      {stage3_11[2],stage3_10[17],stage3_9[18],stage3_8[26],stage3_7[34]}
   );
   gpc2116_5 gpc8646 (
      {stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44]},
      {stage2_8[93]},
      {stage2_9[3]},
      {stage2_10[6], stage2_10[7]},
      {stage3_11[3],stage3_10[18],stage3_9[19],stage3_8[27],stage3_7[35]}
   );
   gpc2116_5 gpc8647 (
      {stage2_7[45], stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[94]},
      {stage2_9[4]},
      {stage2_10[8], stage2_10[9]},
      {stage3_11[4],stage3_10[19],stage3_9[20],stage3_8[28],stage3_7[36]}
   );
   gpc2116_5 gpc8648 (
      {stage2_7[51], stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[95]},
      {stage2_9[5]},
      {stage2_10[10], stage2_10[11]},
      {stage3_11[5],stage3_10[20],stage3_9[21],stage3_8[29],stage3_7[37]}
   );
   gpc2116_5 gpc8649 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62]},
      {stage2_8[96]},
      {stage2_9[6]},
      {stage2_10[12], stage2_10[13]},
      {stage3_11[6],stage3_10[21],stage3_9[22],stage3_8[30],stage3_7[38]}
   );
   gpc2116_5 gpc8650 (
      {stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[97]},
      {stage2_9[7]},
      {stage2_10[14], stage2_10[15]},
      {stage3_11[7],stage3_10[22],stage3_9[23],stage3_8[31],stage3_7[39]}
   );
   gpc2116_5 gpc8651 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73], stage2_7[74]},
      {stage2_8[98]},
      {stage2_9[8]},
      {stage2_10[16], stage2_10[17]},
      {stage3_11[8],stage3_10[23],stage3_9[24],stage3_8[32],stage3_7[40]}
   );
   gpc615_5 gpc8652 (
      {stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78], stage2_7[79]},
      {stage2_8[99]},
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage3_11[9],stage3_10[24],stage3_9[25],stage3_8[33],stage3_7[41]}
   );
   gpc615_5 gpc8653 (
      {stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83], stage2_7[84]},
      {stage2_8[100]},
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage3_11[10],stage3_10[25],stage3_9[26],stage3_8[34],stage3_7[42]}
   );
   gpc606_5 gpc8654 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[0],stage3_11[11],stage3_10[26],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc8655 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[1],stage3_11[12],stage3_10[27],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc8656 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[2],stage3_11[13],stage3_10[28],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc8657 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[3],stage3_11[14],stage3_10[29],stage3_9[30],stage3_8[38]}
   );
   gpc606_5 gpc8658 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[4],stage3_11[15],stage3_10[30],stage3_9[31],stage3_8[39]}
   );
   gpc606_5 gpc8659 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[5],stage3_11[16],stage3_10[31],stage3_9[32],stage3_8[40]}
   );
   gpc606_5 gpc8660 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[6],stage3_11[17],stage3_10[32],stage3_9[33],stage3_8[41]}
   );
   gpc606_5 gpc8661 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[7],stage3_11[18],stage3_10[33],stage3_9[34],stage3_8[42]}
   );
   gpc606_5 gpc8662 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[8],stage3_11[19],stage3_10[34],stage3_9[35],stage3_8[43]}
   );
   gpc606_5 gpc8663 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], stage2_8[160]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[9],stage3_11[20],stage3_10[35],stage3_9[36],stage3_8[44]}
   );
   gpc606_5 gpc8664 (
      {stage2_8[161], stage2_8[162], stage2_8[163], stage2_8[164], stage2_8[165], stage2_8[166]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[10],stage3_11[21],stage3_10[36],stage3_9[37],stage3_8[45]}
   );
   gpc606_5 gpc8665 (
      {stage2_8[167], stage2_8[168], stage2_8[169], stage2_8[170], stage2_8[171], stage2_8[172]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[11],stage3_11[22],stage3_10[37],stage3_9[38],stage3_8[46]}
   );
   gpc606_5 gpc8666 (
      {stage2_9[21], stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[12],stage3_11[23],stage3_10[38],stage3_9[39]}
   );
   gpc606_5 gpc8667 (
      {stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30], stage2_9[31], stage2_9[32]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[13],stage3_11[24],stage3_10[39],stage3_9[40]}
   );
   gpc606_5 gpc8668 (
      {stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37], stage2_9[38]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[14],stage3_11[25],stage3_10[40],stage3_9[41]}
   );
   gpc606_5 gpc8669 (
      {stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43], stage2_9[44]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[15],stage3_11[26],stage3_10[41],stage3_9[42]}
   );
   gpc606_5 gpc8670 (
      {stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49], stage2_9[50]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[16],stage3_11[27],stage3_10[42],stage3_9[43]}
   );
   gpc606_5 gpc8671 (
      {stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[17],stage3_11[28],stage3_10[43],stage3_9[44]}
   );
   gpc606_5 gpc8672 (
      {stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[18],stage3_11[29],stage3_10[44],stage3_9[45]}
   );
   gpc606_5 gpc8673 (
      {stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67], stage2_9[68]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[19],stage3_11[30],stage3_10[45],stage3_9[46]}
   );
   gpc606_5 gpc8674 (
      {stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[20],stage3_11[31],stage3_10[46],stage3_9[47]}
   );
   gpc606_5 gpc8675 (
      {stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[21],stage3_11[32],stage3_10[47],stage3_9[48]}
   );
   gpc606_5 gpc8676 (
      {stage2_9[81], stage2_9[82], stage2_9[83], stage2_9[84], stage2_9[85], stage2_9[86]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[22],stage3_11[33],stage3_10[48],stage3_9[49]}
   );
   gpc606_5 gpc8677 (
      {stage2_9[87], stage2_9[88], stage2_9[89], stage2_9[90], stage2_9[91], stage2_9[92]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[23],stage3_11[34],stage3_10[49],stage3_9[50]}
   );
   gpc606_5 gpc8678 (
      {stage2_9[93], stage2_9[94], stage2_9[95], stage2_9[96], stage2_9[97], stage2_9[98]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[24],stage3_11[35],stage3_10[50],stage3_9[51]}
   );
   gpc606_5 gpc8679 (
      {stage2_9[99], stage2_9[100], stage2_9[101], stage2_9[102], stage2_9[103], stage2_9[104]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[25],stage3_11[36],stage3_10[51],stage3_9[52]}
   );
   gpc215_4 gpc8680 (
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94]},
      {stage2_11[84]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[14],stage3_12[26],stage3_11[37],stage3_10[52]}
   );
   gpc215_4 gpc8681 (
      {stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99]},
      {stage2_11[85]},
      {stage2_12[2], stage2_12[3]},
      {stage3_13[15],stage3_12[27],stage3_11[38],stage3_10[53]}
   );
   gpc215_4 gpc8682 (
      {stage2_10[100], stage2_10[101], stage2_10[102], stage2_10[103], stage2_10[104]},
      {stage2_11[86]},
      {stage2_12[4], stage2_12[5]},
      {stage3_13[16],stage3_12[28],stage3_11[39],stage3_10[54]}
   );
   gpc615_5 gpc8683 (
      {stage2_10[105], stage2_10[106], stage2_10[107], stage2_10[108], stage2_10[109]},
      {stage2_11[87]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[0],stage3_13[17],stage3_12[29],stage3_11[40],stage3_10[55]}
   );
   gpc615_5 gpc8684 (
      {stage2_10[110], stage2_10[111], stage2_10[112], stage2_10[113], stage2_10[114]},
      {stage2_11[88]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[1],stage3_13[18],stage3_12[30],stage3_11[41],stage3_10[56]}
   );
   gpc615_5 gpc8685 (
      {stage2_10[115], stage2_10[116], stage2_10[117], stage2_10[118], stage2_10[119]},
      {stage2_11[89]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[2],stage3_13[19],stage3_12[31],stage3_11[42],stage3_10[57]}
   );
   gpc615_5 gpc8686 (
      {stage2_10[120], stage2_10[121], stage2_10[122], stage2_10[123], stage2_10[124]},
      {stage2_11[90]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[3],stage3_13[20],stage3_12[32],stage3_11[43],stage3_10[58]}
   );
   gpc606_5 gpc8687 (
      {stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[4],stage3_13[21],stage3_12[33],stage3_11[44]}
   );
   gpc606_5 gpc8688 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[5],stage3_13[22],stage3_12[34],stage3_11[45]}
   );
   gpc606_5 gpc8689 (
      {stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[6],stage3_13[23],stage3_12[35],stage3_11[46]}
   );
   gpc606_5 gpc8690 (
      {stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[7],stage3_13[24],stage3_12[36],stage3_11[47]}
   );
   gpc615_5 gpc8691 (
      {stage2_11[115], stage2_11[116], stage2_11[117], stage2_11[118], stage2_11[119]},
      {stage2_12[30]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[8],stage3_13[25],stage3_12[37],stage3_11[48]}
   );
   gpc615_5 gpc8692 (
      {stage2_11[120], stage2_11[121], stage2_11[122], stage2_11[123], stage2_11[124]},
      {stage2_12[31]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[9],stage3_13[26],stage3_12[38],stage3_11[49]}
   );
   gpc606_5 gpc8693 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[6],stage3_14[10],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc8694 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[7],stage3_14[11],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc8695 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[8],stage3_14[12],stage3_13[29],stage3_12[41]}
   );
   gpc606_5 gpc8696 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[9],stage3_14[13],stage3_13[30],stage3_12[42]}
   );
   gpc606_5 gpc8697 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[10],stage3_14[14],stage3_13[31],stage3_12[43]}
   );
   gpc606_5 gpc8698 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[11],stage3_14[15],stage3_13[32],stage3_12[44]}
   );
   gpc606_5 gpc8699 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[12],stage3_14[16],stage3_13[33],stage3_12[45]}
   );
   gpc606_5 gpc8700 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[13],stage3_14[17],stage3_13[34],stage3_12[46]}
   );
   gpc606_5 gpc8701 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[14],stage3_14[18],stage3_13[35],stage3_12[47]}
   );
   gpc606_5 gpc8702 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[15],stage3_14[19],stage3_13[36],stage3_12[48]}
   );
   gpc623_5 gpc8703 (
      {stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_13[36], stage2_13[37]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[16],stage3_14[20],stage3_13[37],stage3_12[49]}
   );
   gpc623_5 gpc8704 (
      {stage2_12[95], stage2_12[96], stage2_12[97]},
      {stage2_13[38], stage2_13[39]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[17],stage3_14[21],stage3_13[38],stage3_12[50]}
   );
   gpc615_5 gpc8705 (
      {stage2_13[40], stage2_13[41], stage2_13[42], stage2_13[43], stage2_13[44]},
      {stage2_14[72]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[18],stage3_14[22],stage3_13[39]}
   );
   gpc615_5 gpc8706 (
      {stage2_13[45], stage2_13[46], stage2_13[47], stage2_13[48], stage2_13[49]},
      {stage2_14[73]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[19],stage3_14[23],stage3_13[40]}
   );
   gpc615_5 gpc8707 (
      {stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53], stage2_13[54]},
      {stage2_14[74]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[20],stage3_14[24],stage3_13[41]}
   );
   gpc615_5 gpc8708 (
      {stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_14[75]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[21],stage3_14[25],stage3_13[42]}
   );
   gpc615_5 gpc8709 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64]},
      {stage2_14[76]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[22],stage3_14[26],stage3_13[43]}
   );
   gpc615_5 gpc8710 (
      {stage2_13[65], stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69]},
      {stage2_14[77]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[23],stage3_14[27],stage3_13[44]}
   );
   gpc606_5 gpc8711 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[18],stage3_15[24],stage3_14[28]}
   );
   gpc606_5 gpc8712 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[19],stage3_15[25],stage3_14[29]}
   );
   gpc615_5 gpc8713 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94]},
      {stage2_15[36]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[20],stage3_15[26],stage3_14[30]}
   );
   gpc615_5 gpc8714 (
      {stage2_14[95], stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99]},
      {stage2_15[37]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[21],stage3_15[27],stage3_14[31]}
   );
   gpc615_5 gpc8715 (
      {stage2_14[100], stage2_14[101], stage2_14[102], stage2_14[103], stage2_14[104]},
      {stage2_15[38]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[22],stage3_15[28],stage3_14[32]}
   );
   gpc615_5 gpc8716 (
      {stage2_14[105], stage2_14[106], stage2_14[107], stage2_14[108], stage2_14[109]},
      {stage2_15[39]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[23],stage3_15[29],stage3_14[33]}
   );
   gpc615_5 gpc8717 (
      {stage2_14[110], stage2_14[111], stage2_14[112], stage2_14[113], stage2_14[114]},
      {stage2_15[40]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[24],stage3_15[30],stage3_14[34]}
   );
   gpc207_4 gpc8718 (
      {stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[7],stage3_17[13],stage3_16[25],stage3_15[31]}
   );
   gpc615_5 gpc8719 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[42]},
      {stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7]},
      {stage3_19[0],stage3_18[8],stage3_17[14],stage3_16[26],stage3_15[32]}
   );
   gpc615_5 gpc8720 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[43]},
      {stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13]},
      {stage3_19[1],stage3_18[9],stage3_17[15],stage3_16[27],stage3_15[33]}
   );
   gpc615_5 gpc8721 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[44]},
      {stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19]},
      {stage3_19[2],stage3_18[10],stage3_17[16],stage3_16[28],stage3_15[34]}
   );
   gpc615_5 gpc8722 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[45]},
      {stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25]},
      {stage3_19[3],stage3_18[11],stage3_17[17],stage3_16[29],stage3_15[35]}
   );
   gpc615_5 gpc8723 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[46]},
      {stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31]},
      {stage3_19[4],stage3_18[12],stage3_17[18],stage3_16[30],stage3_15[36]}
   );
   gpc615_5 gpc8724 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[47]},
      {stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37]},
      {stage3_19[5],stage3_18[13],stage3_17[19],stage3_16[31],stage3_15[37]}
   );
   gpc615_5 gpc8725 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[48]},
      {stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43]},
      {stage3_19[6],stage3_18[14],stage3_17[20],stage3_16[32],stage3_15[38]}
   );
   gpc615_5 gpc8726 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[49]},
      {stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49]},
      {stage3_19[7],stage3_18[15],stage3_17[21],stage3_16[33],stage3_15[39]}
   );
   gpc615_5 gpc8727 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[50]},
      {stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55]},
      {stage3_19[8],stage3_18[16],stage3_17[22],stage3_16[34],stage3_15[40]}
   );
   gpc615_5 gpc8728 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[51]},
      {stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61]},
      {stage3_19[9],stage3_18[17],stage3_17[23],stage3_16[35],stage3_15[41]}
   );
   gpc615_5 gpc8729 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[52]},
      {stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67]},
      {stage3_19[10],stage3_18[18],stage3_17[24],stage3_16[36],stage3_15[42]}
   );
   gpc615_5 gpc8730 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[53]},
      {stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73]},
      {stage3_19[11],stage3_18[19],stage3_17[25],stage3_16[37],stage3_15[43]}
   );
   gpc606_5 gpc8731 (
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[12],stage3_18[20],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc8732 (
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[13],stage3_18[21],stage3_17[27],stage3_16[39]}
   );
   gpc606_5 gpc8733 (
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[14],stage3_18[22],stage3_17[28],stage3_16[40]}
   );
   gpc606_5 gpc8734 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[15],stage3_18[23],stage3_17[29],stage3_16[41]}
   );
   gpc606_5 gpc8735 (
      {stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[16],stage3_18[24],stage3_17[30],stage3_16[42]}
   );
   gpc606_5 gpc8736 (
      {stage2_16[84], stage2_16[85], stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89]},
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage3_20[5],stage3_19[17],stage3_18[25],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc8737 (
      {stage2_16[90], stage2_16[91], stage2_16[92], stage2_16[93], stage2_16[94], stage2_16[95]},
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41]},
      {stage3_20[6],stage3_19[18],stage3_18[26],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc8738 (
      {stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[7],stage3_19[19],stage3_18[27],stage3_17[33]}
   );
   gpc2135_5 gpc8739 (
      {stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[1],stage3_20[8],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc8740 (
      {stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50], stage2_18[51]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[2],stage3_20[9],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc8741 (
      {stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55], stage2_18[56]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[3],stage3_20[10],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc8742 (
      {stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60], stage2_18[61]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[4],stage3_20[11],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc8743 (
      {stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[5],stage3_20[12],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc8744 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[6],stage3_20[13],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc8745 (
      {stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75], stage2_18[76]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[7],stage3_20[14],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc8746 (
      {stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80], stage2_18[81]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[8],stage3_20[15],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc8747 (
      {stage2_18[82], stage2_18[83], stage2_18[84], stage2_18[85], stage2_18[86]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[9],stage3_20[16],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc8748 (
      {stage2_18[87], stage2_18[88], stage2_18[89], stage2_18[90], stage2_18[91]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[10],stage3_20[17],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc8749 (
      {stage2_18[92], stage2_18[93], stage2_18[94], stage2_18[95], stage2_18[96]},
      {stage2_19[36], stage2_19[37], stage2_19[38]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[11],stage3_20[18],stage3_19[30],stage3_18[38]}
   );
   gpc2135_5 gpc8750 (
      {stage2_18[97], stage2_18[98], stage2_18[99], stage2_18[100], stage2_18[101]},
      {stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[12],stage3_20[19],stage3_19[31],stage3_18[39]}
   );
   gpc2135_5 gpc8751 (
      {stage2_18[102], stage2_18[103], stage2_18[104], stage2_18[105], stage2_18[106]},
      {stage2_19[42], stage2_19[43], stage2_19[44]},
      {stage2_20[12]},
      {stage2_21[24], stage2_21[25]},
      {stage3_22[12],stage3_21[13],stage3_20[20],stage3_19[32],stage3_18[40]}
   );
   gpc2135_5 gpc8752 (
      {stage2_18[107], stage2_18[108], stage2_18[109], stage2_18[110], stage2_18[111]},
      {stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[13]},
      {stage2_21[26], stage2_21[27]},
      {stage3_22[13],stage3_21[14],stage3_20[21],stage3_19[33],stage3_18[41]}
   );
   gpc2135_5 gpc8753 (
      {stage2_18[112], stage2_18[113], stage2_18[114], stage2_18[115], stage2_18[116]},
      {stage2_19[48], stage2_19[49], stage2_19[50]},
      {stage2_20[14]},
      {stage2_21[28], stage2_21[29]},
      {stage3_22[14],stage3_21[15],stage3_20[22],stage3_19[34],stage3_18[42]}
   );
   gpc2135_5 gpc8754 (
      {stage2_18[117], stage2_18[118], stage2_18[119], stage2_18[120], stage2_18[121]},
      {stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_20[15]},
      {stage2_21[30], stage2_21[31]},
      {stage3_22[15],stage3_21[16],stage3_20[23],stage3_19[35],stage3_18[43]}
   );
   gpc2135_5 gpc8755 (
      {stage2_18[122], stage2_18[123], stage2_18[124], stage2_18[125], stage2_18[126]},
      {stage2_19[54], stage2_19[55], stage2_19[56]},
      {stage2_20[16]},
      {stage2_21[32], stage2_21[33]},
      {stage3_22[16],stage3_21[17],stage3_20[24],stage3_19[36],stage3_18[44]}
   );
   gpc2135_5 gpc8756 (
      {stage2_18[127], stage2_18[128], stage2_18[129], stage2_18[130], stage2_18[131]},
      {stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage2_20[17]},
      {stage2_21[34], stage2_21[35]},
      {stage3_22[17],stage3_21[18],stage3_20[25],stage3_19[37],stage3_18[45]}
   );
   gpc2135_5 gpc8757 (
      {stage2_18[132], stage2_18[133], stage2_18[134], stage2_18[135], stage2_18[136]},
      {stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[18]},
      {stage2_21[36], stage2_21[37]},
      {stage3_22[18],stage3_21[19],stage3_20[26],stage3_19[38],stage3_18[46]}
   );
   gpc2135_5 gpc8758 (
      {stage2_18[137], stage2_18[138], stage2_18[139], stage2_18[140], stage2_18[141]},
      {stage2_19[63], stage2_19[64], stage2_19[65]},
      {stage2_20[19]},
      {stage2_21[38], stage2_21[39]},
      {stage3_22[19],stage3_21[20],stage3_20[27],stage3_19[39],stage3_18[47]}
   );
   gpc2135_5 gpc8759 (
      {stage2_18[142], stage2_18[143], stage2_18[144], stage2_18[145], stage2_18[146]},
      {stage2_19[66], stage2_19[67], stage2_19[68]},
      {stage2_20[20]},
      {stage2_21[40], stage2_21[41]},
      {stage3_22[20],stage3_21[21],stage3_20[28],stage3_19[40],stage3_18[48]}
   );
   gpc615_5 gpc8760 (
      {stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72], stage2_19[73]},
      {stage2_20[21]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[0],stage3_22[21],stage3_21[22],stage3_20[29],stage3_19[41]}
   );
   gpc615_5 gpc8761 (
      {stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77], stage2_19[78]},
      {stage2_20[22]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[1],stage3_22[22],stage3_21[23],stage3_20[30],stage3_19[42]}
   );
   gpc615_5 gpc8762 (
      {stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82], stage2_19[83]},
      {stage2_20[23]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[2],stage3_22[23],stage3_21[24],stage3_20[31],stage3_19[43]}
   );
   gpc615_5 gpc8763 (
      {stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87], stage2_19[88]},
      {stage2_20[24]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[3],stage3_22[24],stage3_21[25],stage3_20[32],stage3_19[44]}
   );
   gpc615_5 gpc8764 (
      {stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92], stage2_19[93]},
      {stage2_20[25]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[4],stage3_22[25],stage3_21[26],stage3_20[33],stage3_19[45]}
   );
   gpc606_5 gpc8765 (
      {stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30], stage2_20[31]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[26],stage3_21[27],stage3_20[34]}
   );
   gpc606_5 gpc8766 (
      {stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35], stage2_20[36], stage2_20[37]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[27],stage3_21[28],stage3_20[35]}
   );
   gpc606_5 gpc8767 (
      {stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[28],stage3_21[29],stage3_20[36]}
   );
   gpc606_5 gpc8768 (
      {stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47], stage2_20[48], stage2_20[49]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[8],stage3_22[29],stage3_21[30],stage3_20[37]}
   );
   gpc606_5 gpc8769 (
      {stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53], stage2_20[54], stage2_20[55]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[9],stage3_22[30],stage3_21[31],stage3_20[38]}
   );
   gpc606_5 gpc8770 (
      {stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59], stage2_20[60], stage2_20[61]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[10],stage3_22[31],stage3_21[32],stage3_20[39]}
   );
   gpc615_5 gpc8771 (
      {stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65], stage2_20[66]},
      {stage2_21[72]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[11],stage3_22[32],stage3_21[33],stage3_20[40]}
   );
   gpc615_5 gpc8772 (
      {stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage2_21[73]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage3_24[7],stage3_23[12],stage3_22[33],stage3_21[34],stage3_20[41]}
   );
   gpc606_5 gpc8773 (
      {stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77], stage2_21[78], stage2_21[79]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[8],stage3_23[13],stage3_22[34],stage3_21[35]}
   );
   gpc606_5 gpc8774 (
      {stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83], stage2_21[84], stage2_21[85]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[9],stage3_23[14],stage3_22[35],stage3_21[36]}
   );
   gpc615_5 gpc8775 (
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[10],stage3_23[15],stage3_22[36]}
   );
   gpc615_5 gpc8776 (
      {stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[11],stage3_23[16],stage3_22[37]}
   );
   gpc615_5 gpc8777 (
      {stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61], stage2_22[62]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[12],stage3_23[17],stage3_22[38]}
   );
   gpc615_5 gpc8778 (
      {stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66], stage2_22[67]},
      {stage2_23[15]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[5],stage3_24[13],stage3_23[18],stage3_22[39]}
   );
   gpc615_5 gpc8779 (
      {stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71], stage2_22[72]},
      {stage2_23[16]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[6],stage3_24[14],stage3_23[19],stage3_22[40]}
   );
   gpc615_5 gpc8780 (
      {stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76], stage2_22[77]},
      {stage2_23[17]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[7],stage3_24[15],stage3_23[20],stage3_22[41]}
   );
   gpc615_5 gpc8781 (
      {stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81], stage2_22[82]},
      {stage2_23[18]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[8],stage3_24[16],stage3_23[21],stage3_22[42]}
   );
   gpc615_5 gpc8782 (
      {stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86], stage2_22[87]},
      {stage2_23[19]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[9],stage3_24[17],stage3_23[22],stage3_22[43]}
   );
   gpc615_5 gpc8783 (
      {stage2_22[88], stage2_22[89], stage2_22[90], stage2_22[91], stage2_22[92]},
      {stage2_23[20]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[10],stage3_24[18],stage3_23[23],stage3_22[44]}
   );
   gpc615_5 gpc8784 (
      {stage2_22[93], stage2_22[94], stage2_22[95], stage2_22[96], stage2_22[97]},
      {stage2_23[21]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[11],stage3_24[19],stage3_23[24],stage3_22[45]}
   );
   gpc615_5 gpc8785 (
      {stage2_22[98], stage2_22[99], stage2_22[100], stage2_22[101], stage2_22[102]},
      {stage2_23[22]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[12],stage3_24[20],stage3_23[25],stage3_22[46]}
   );
   gpc615_5 gpc8786 (
      {stage2_22[103], stage2_22[104], stage2_22[105], stage2_22[106], stage2_22[107]},
      {stage2_23[23]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[13],stage3_24[21],stage3_23[26],stage3_22[47]}
   );
   gpc615_5 gpc8787 (
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28]},
      {stage2_24[72]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[12],stage3_25[14],stage3_24[22],stage3_23[27]}
   );
   gpc615_5 gpc8788 (
      {stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33]},
      {stage2_24[73]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[13],stage3_25[15],stage3_24[23],stage3_23[28]}
   );
   gpc615_5 gpc8789 (
      {stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage2_24[74]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[14],stage3_25[16],stage3_24[24],stage3_23[29]}
   );
   gpc615_5 gpc8790 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43]},
      {stage2_24[75]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[15],stage3_25[17],stage3_24[25],stage3_23[30]}
   );
   gpc615_5 gpc8791 (
      {stage2_23[44], stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48]},
      {stage2_24[76]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[16],stage3_25[18],stage3_24[26],stage3_23[31]}
   );
   gpc615_5 gpc8792 (
      {stage2_23[49], stage2_23[50], stage2_23[51], stage2_23[52], stage2_23[53]},
      {stage2_24[77]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[17],stage3_25[19],stage3_24[27],stage3_23[32]}
   );
   gpc615_5 gpc8793 (
      {stage2_23[54], stage2_23[55], stage2_23[56], stage2_23[57], stage2_23[58]},
      {stage2_24[78]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[18],stage3_25[20],stage3_24[28],stage3_23[33]}
   );
   gpc615_5 gpc8794 (
      {stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62], stage2_23[63]},
      {stage2_24[79]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[19],stage3_25[21],stage3_24[29],stage3_23[34]}
   );
   gpc615_5 gpc8795 (
      {stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_24[80]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[20],stage3_25[22],stage3_24[30],stage3_23[35]}
   );
   gpc615_5 gpc8796 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73]},
      {stage2_24[81]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[21],stage3_25[23],stage3_24[31],stage3_23[36]}
   );
   gpc615_5 gpc8797 (
      {stage2_23[74], stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78]},
      {stage2_24[82]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[22],stage3_25[24],stage3_24[32],stage3_23[37]}
   );
   gpc615_5 gpc8798 (
      {stage2_23[79], stage2_23[80], stage2_23[81], stage2_23[82], stage2_23[83]},
      {stage2_24[83]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[23],stage3_25[25],stage3_24[33],stage3_23[38]}
   );
   gpc615_5 gpc8799 (
      {stage2_23[84], stage2_23[85], stage2_23[86], stage2_23[87], stage2_23[88]},
      {stage2_24[84]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[24],stage3_25[26],stage3_24[34],stage3_23[39]}
   );
   gpc606_5 gpc8800 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[13],stage3_26[25],stage3_25[27]}
   );
   gpc606_5 gpc8801 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[1],stage3_27[14],stage3_26[26],stage3_25[28]}
   );
   gpc606_5 gpc8802 (
      {stage2_25[90], stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[2],stage3_27[15],stage3_26[27],stage3_25[29]}
   );
   gpc606_5 gpc8803 (
      {stage2_25[96], stage2_25[97], stage2_25[98], stage2_25[99], stage2_25[100], stage2_25[101]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[3],stage3_27[16],stage3_26[28],stage3_25[30]}
   );
   gpc117_4 gpc8804 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6]},
      {stage2_27[24]},
      {stage2_28[0]},
      {stage3_29[4],stage3_28[4],stage3_27[17],stage3_26[29]}
   );
   gpc117_4 gpc8805 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12], stage2_26[13]},
      {stage2_27[25]},
      {stage2_28[1]},
      {stage3_29[5],stage3_28[5],stage3_27[18],stage3_26[30]}
   );
   gpc117_4 gpc8806 (
      {stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_27[26]},
      {stage2_28[2]},
      {stage3_29[6],stage3_28[6],stage3_27[19],stage3_26[31]}
   );
   gpc117_4 gpc8807 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[27]},
      {stage2_28[3]},
      {stage3_29[7],stage3_28[7],stage3_27[20],stage3_26[32]}
   );
   gpc117_4 gpc8808 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34]},
      {stage2_27[28]},
      {stage2_28[4]},
      {stage3_29[8],stage3_28[8],stage3_27[21],stage3_26[33]}
   );
   gpc117_4 gpc8809 (
      {stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage2_27[29]},
      {stage2_28[5]},
      {stage3_29[9],stage3_28[9],stage3_27[22],stage3_26[34]}
   );
   gpc117_4 gpc8810 (
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48]},
      {stage2_27[30]},
      {stage2_28[6]},
      {stage3_29[10],stage3_28[10],stage3_27[23],stage3_26[35]}
   );
   gpc117_4 gpc8811 (
      {stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55]},
      {stage2_27[31]},
      {stage2_28[7]},
      {stage3_29[11],stage3_28[11],stage3_27[24],stage3_26[36]}
   );
   gpc117_4 gpc8812 (
      {stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[32]},
      {stage2_28[8]},
      {stage3_29[12],stage3_28[12],stage3_27[25],stage3_26[37]}
   );
   gpc117_4 gpc8813 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69]},
      {stage2_27[33]},
      {stage2_28[9]},
      {stage3_29[13],stage3_28[13],stage3_27[26],stage3_26[38]}
   );
   gpc117_4 gpc8814 (
      {stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76]},
      {stage2_27[34]},
      {stage2_28[10]},
      {stage3_29[14],stage3_28[14],stage3_27[27],stage3_26[39]}
   );
   gpc117_4 gpc8815 (
      {stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage2_27[35]},
      {stage2_28[11]},
      {stage3_29[15],stage3_28[15],stage3_27[28],stage3_26[40]}
   );
   gpc117_4 gpc8816 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88], stage2_26[89], stage2_26[90]},
      {stage2_27[36]},
      {stage2_28[12]},
      {stage3_29[16],stage3_28[16],stage3_27[29],stage3_26[41]}
   );
   gpc117_4 gpc8817 (
      {stage2_26[91], stage2_26[92], stage2_26[93], stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97]},
      {stage2_27[37]},
      {stage2_28[13]},
      {stage3_29[17],stage3_28[17],stage3_27[30],stage3_26[42]}
   );
   gpc117_4 gpc8818 (
      {stage2_26[98], stage2_26[99], stage2_26[100], stage2_26[101], stage2_26[102], stage2_26[103], stage2_26[104]},
      {stage2_27[38]},
      {stage2_28[14]},
      {stage3_29[18],stage3_28[18],stage3_27[31],stage3_26[43]}
   );
   gpc117_4 gpc8819 (
      {stage2_26[105], stage2_26[106], stage2_26[107], stage2_26[108], stage2_26[109], stage2_26[110], stage2_26[111]},
      {stage2_27[39]},
      {stage2_28[15]},
      {stage3_29[19],stage3_28[19],stage3_27[32],stage3_26[44]}
   );
   gpc117_4 gpc8820 (
      {stage2_26[112], stage2_26[113], stage2_26[114], stage2_26[115], stage2_26[116], stage2_26[117], stage2_26[118]},
      {stage2_27[40]},
      {stage2_28[16]},
      {stage3_29[20],stage3_28[20],stage3_27[33],stage3_26[45]}
   );
   gpc117_4 gpc8821 (
      {stage2_26[119], stage2_26[120], stage2_26[121], stage2_26[122], stage2_26[123], stage2_26[124], stage2_26[125]},
      {stage2_27[41]},
      {stage2_28[17]},
      {stage3_29[21],stage3_28[21],stage3_27[34],stage3_26[46]}
   );
   gpc7_3 gpc8822 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48]},
      {stage3_29[22],stage3_28[22],stage3_27[35]}
   );
   gpc7_3 gpc8823 (
      {stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55]},
      {stage3_29[23],stage3_28[23],stage3_27[36]}
   );
   gpc207_4 gpc8824 (
      {stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_29[0], stage2_29[1]},
      {stage3_30[0],stage3_29[24],stage3_28[24],stage3_27[37]}
   );
   gpc207_4 gpc8825 (
      {stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_29[2], stage2_29[3]},
      {stage3_30[1],stage3_29[25],stage3_28[25],stage3_27[38]}
   );
   gpc606_5 gpc8826 (
      {stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73], stage2_27[74], stage2_27[75]},
      {stage2_29[4], stage2_29[5], stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9]},
      {stage3_31[0],stage3_30[2],stage3_29[26],stage3_28[26],stage3_27[39]}
   );
   gpc606_5 gpc8827 (
      {stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80], stage2_27[81]},
      {stage2_29[10], stage2_29[11], stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15]},
      {stage3_31[1],stage3_30[3],stage3_29[27],stage3_28[27],stage3_27[40]}
   );
   gpc615_5 gpc8828 (
      {stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], 1'b0},
      {stage2_28[18]},
      {stage2_29[16], stage2_29[17], stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage3_31[2],stage3_30[4],stage3_29[28],stage3_28[28],stage3_27[41]}
   );
   gpc615_5 gpc8829 (
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_29[22]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[5],stage3_29[29],stage3_28[29]}
   );
   gpc615_5 gpc8830 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[23]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[6],stage3_29[30],stage3_28[30]}
   );
   gpc615_5 gpc8831 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[24]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[7],stage3_29[31],stage3_28[31]}
   );
   gpc615_5 gpc8832 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[25]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[8],stage3_29[32],stage3_28[32]}
   );
   gpc615_5 gpc8833 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[26]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[7],stage3_30[9],stage3_29[33],stage3_28[33]}
   );
   gpc1163_5 gpc8834 (
      {stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[5],stage3_31[8],stage3_30[10],stage3_29[34]}
   );
   gpc1163_5 gpc8835 (
      {stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[6],stage3_31[9],stage3_30[11],stage3_29[35]}
   );
   gpc1163_5 gpc8836 (
      {stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[7],stage3_31[10],stage3_30[12],stage3_29[36]}
   );
   gpc1163_5 gpc8837 (
      {stage2_29[36], stage2_29[37], stage2_29[38]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[8],stage3_31[11],stage3_30[13],stage3_29[37]}
   );
   gpc1163_5 gpc8838 (
      {stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[9],stage3_31[12],stage3_30[14],stage3_29[38]}
   );
   gpc606_5 gpc8839 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[10],stage3_31[13],stage3_30[15],stage3_29[39]}
   );
   gpc606_5 gpc8840 (
      {stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[11],stage3_31[14],stage3_30[16],stage3_29[40]}
   );
   gpc606_5 gpc8841 (
      {stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[12],stage3_31[15],stage3_30[17],stage3_29[41]}
   );
   gpc606_5 gpc8842 (
      {stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[13],stage3_31[16],stage3_30[18],stage3_29[42]}
   );
   gpc606_5 gpc8843 (
      {stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[14],stage3_31[17],stage3_30[19],stage3_29[43]}
   );
   gpc606_5 gpc8844 (
      {stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[15],stage3_31[18],stage3_30[20],stage3_29[44]}
   );
   gpc606_5 gpc8845 (
      {stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[16],stage3_31[19],stage3_30[21],stage3_29[45]}
   );
   gpc606_5 gpc8846 (
      {stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[17],stage3_31[20],stage3_30[22],stage3_29[46]}
   );
   gpc606_5 gpc8847 (
      {stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[18],stage3_31[21],stage3_30[23],stage3_29[47]}
   );
   gpc606_5 gpc8848 (
      {stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101]},
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage3_33[14],stage3_32[19],stage3_31[22],stage3_30[24],stage3_29[48]}
   );
   gpc1163_5 gpc8849 (
      {stage2_30[60], stage2_30[61], stage2_30[62]},
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_32[5]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[15],stage3_32[20],stage3_31[23],stage3_30[25]}
   );
   gpc615_5 gpc8850 (
      {stage2_30[63], stage2_30[64], stage2_30[65], stage2_30[66], stage2_30[67]},
      {stage2_31[71]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[16],stage3_32[21],stage3_31[24],stage3_30[26]}
   );
   gpc615_5 gpc8851 (
      {stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71], stage2_30[72]},
      {stage2_31[72]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[17],stage3_32[22],stage3_31[25],stage3_30[27]}
   );
   gpc615_5 gpc8852 (
      {stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[73]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[18],stage3_32[23],stage3_31[26],stage3_30[28]}
   );
   gpc615_5 gpc8853 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82]},
      {stage2_31[74]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[19],stage3_32[24],stage3_31[27],stage3_30[29]}
   );
   gpc615_5 gpc8854 (
      {stage2_30[83], stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87]},
      {stage2_31[75]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[20],stage3_32[25],stage3_31[28],stage3_30[30]}
   );
   gpc615_5 gpc8855 (
      {stage2_30[88], stage2_30[89], stage2_30[90], stage2_30[91], stage2_30[92]},
      {stage2_31[76]},
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40], stage2_32[41]},
      {stage3_34[6],stage3_33[21],stage3_32[26],stage3_31[29],stage3_30[31]}
   );
   gpc606_5 gpc8856 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[0],stage3_34[7],stage3_33[22],stage3_32[27],stage3_31[30]}
   );
   gpc606_5 gpc8857 (
      {stage2_31[83], stage2_31[84], stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88]},
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12]},
      {stage3_35[1],stage3_34[8],stage3_33[23],stage3_32[28],stage3_31[31]}
   );
   gpc606_5 gpc8858 (
      {stage2_31[89], stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18]},
      {stage3_35[2],stage3_34[9],stage3_33[24],stage3_32[29],stage3_31[32]}
   );
   gpc606_5 gpc8859 (
      {stage2_31[95], stage2_31[96], stage2_31[97], stage2_31[98], stage2_31[99], stage2_31[100]},
      {stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24]},
      {stage3_35[3],stage3_34[10],stage3_33[25],stage3_32[30],stage3_31[33]}
   );
   gpc606_5 gpc8860 (
      {stage2_31[101], stage2_31[102], stage2_31[103], stage2_31[104], stage2_31[105], stage2_31[106]},
      {stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29], stage2_33[30]},
      {stage3_35[4],stage3_34[11],stage3_33[26],stage3_32[31],stage3_31[34]}
   );
   gpc606_5 gpc8861 (
      {stage2_31[107], stage2_31[108], stage2_31[109], stage2_31[110], stage2_31[111], stage2_31[112]},
      {stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35], stage2_33[36]},
      {stage3_35[5],stage3_34[12],stage3_33[27],stage3_32[32],stage3_31[35]}
   );
   gpc606_5 gpc8862 (
      {stage2_31[113], stage2_31[114], stage2_31[115], stage2_31[116], stage2_31[117], stage2_31[118]},
      {stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41], stage2_33[42]},
      {stage3_35[6],stage3_34[13],stage3_33[28],stage3_32[33],stage3_31[36]}
   );
   gpc615_5 gpc8863 (
      {stage2_31[119], stage2_31[120], stage2_31[121], stage2_31[122], stage2_31[123]},
      {stage2_32[42]},
      {stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48]},
      {stage3_35[7],stage3_34[14],stage3_33[29],stage3_32[34],stage3_31[37]}
   );
   gpc1163_5 gpc8864 (
      {stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54]},
      {stage2_34[0]},
      {stage2_35[0]},
      {stage3_36[0],stage3_35[8],stage3_34[15],stage3_33[30],stage3_32[35]}
   );
   gpc1163_5 gpc8865 (
      {stage2_32[46], stage2_32[47], stage2_32[48]},
      {stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59], stage2_33[60]},
      {stage2_34[1]},
      {stage2_35[1]},
      {stage3_36[1],stage3_35[9],stage3_34[16],stage3_33[31],stage3_32[36]}
   );
   gpc1163_5 gpc8866 (
      {stage2_32[49], stage2_32[50], stage2_32[51]},
      {stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65], stage2_33[66]},
      {stage2_34[2]},
      {stage2_35[2]},
      {stage3_36[2],stage3_35[10],stage3_34[17],stage3_33[32],stage3_32[37]}
   );
   gpc1163_5 gpc8867 (
      {stage2_32[52], stage2_32[53], stage2_32[54]},
      {stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71], stage2_33[72]},
      {stage2_34[3]},
      {stage2_35[3]},
      {stage3_36[3],stage3_35[11],stage3_34[18],stage3_33[33],stage3_32[38]}
   );
   gpc1163_5 gpc8868 (
      {stage2_32[55], stage2_32[56], stage2_32[57]},
      {stage2_33[73], stage2_33[74], stage2_33[75], stage2_33[76], stage2_33[77], stage2_33[78]},
      {stage2_34[4]},
      {stage2_35[4]},
      {stage3_36[4],stage3_35[12],stage3_34[19],stage3_33[34],stage3_32[39]}
   );
   gpc1163_5 gpc8869 (
      {stage2_32[58], stage2_32[59], stage2_32[60]},
      {stage2_33[79], stage2_33[80], stage2_33[81], stage2_33[82], stage2_33[83], stage2_33[84]},
      {stage2_34[5]},
      {stage2_35[5]},
      {stage3_36[5],stage3_35[13],stage3_34[20],stage3_33[35],stage3_32[40]}
   );
   gpc1163_5 gpc8870 (
      {stage2_32[61], stage2_32[62], stage2_32[63]},
      {stage2_33[85], stage2_33[86], stage2_33[87], stage2_33[88], stage2_33[89], stage2_33[90]},
      {stage2_34[6]},
      {stage2_35[6]},
      {stage3_36[6],stage3_35[14],stage3_34[21],stage3_33[36],stage3_32[41]}
   );
   gpc606_5 gpc8871 (
      {stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68], stage2_32[69]},
      {stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11], stage2_34[12]},
      {stage3_36[7],stage3_35[15],stage3_34[22],stage3_33[37],stage3_32[42]}
   );
   gpc606_5 gpc8872 (
      {stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74], stage2_32[75]},
      {stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17], stage2_34[18]},
      {stage3_36[8],stage3_35[16],stage3_34[23],stage3_33[38],stage3_32[43]}
   );
   gpc606_5 gpc8873 (
      {stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80], stage2_32[81]},
      {stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23], stage2_34[24]},
      {stage3_36[9],stage3_35[17],stage3_34[24],stage3_33[39],stage3_32[44]}
   );
   gpc606_5 gpc8874 (
      {stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86], stage2_32[87]},
      {stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29], stage2_34[30]},
      {stage3_36[10],stage3_35[18],stage3_34[25],stage3_33[40],stage3_32[45]}
   );
   gpc606_5 gpc8875 (
      {stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92], stage2_32[93]},
      {stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35], stage2_34[36]},
      {stage3_36[11],stage3_35[19],stage3_34[26],stage3_33[41],stage3_32[46]}
   );
   gpc606_5 gpc8876 (
      {stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98], stage2_32[99]},
      {stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41], stage2_34[42]},
      {stage3_36[12],stage3_35[20],stage3_34[27],stage3_33[42],stage3_32[47]}
   );
   gpc606_5 gpc8877 (
      {stage2_32[100], stage2_32[101], stage2_32[102], stage2_32[103], stage2_32[104], stage2_32[105]},
      {stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47], stage2_34[48]},
      {stage3_36[13],stage3_35[21],stage3_34[28],stage3_33[43],stage3_32[48]}
   );
   gpc606_5 gpc8878 (
      {stage2_32[106], stage2_32[107], stage2_32[108], stage2_32[109], stage2_32[110], stage2_32[111]},
      {stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53], stage2_34[54]},
      {stage3_36[14],stage3_35[22],stage3_34[29],stage3_33[44],stage3_32[49]}
   );
   gpc615_5 gpc8879 (
      {stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage2_35[7]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[15],stage3_35[23],stage3_34[30]}
   );
   gpc615_5 gpc8880 (
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64]},
      {stage2_35[8]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[1],stage3_36[16],stage3_35[24],stage3_34[31]}
   );
   gpc615_5 gpc8881 (
      {stage2_34[65], stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69]},
      {stage2_35[9]},
      {stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage3_38[2],stage3_37[2],stage3_36[17],stage3_35[25],stage3_34[32]}
   );
   gpc615_5 gpc8882 (
      {stage2_34[70], stage2_34[71], stage2_34[72], stage2_34[73], stage2_34[74]},
      {stage2_35[10]},
      {stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21], stage2_36[22], stage2_36[23]},
      {stage3_38[3],stage3_37[3],stage3_36[18],stage3_35[26],stage3_34[33]}
   );
   gpc615_5 gpc8883 (
      {stage2_34[75], stage2_34[76], stage2_34[77], stage2_34[78], stage2_34[79]},
      {stage2_35[11]},
      {stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27], stage2_36[28], stage2_36[29]},
      {stage3_38[4],stage3_37[4],stage3_36[19],stage3_35[27],stage3_34[34]}
   );
   gpc615_5 gpc8884 (
      {stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83], stage2_34[84]},
      {stage2_35[12]},
      {stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35]},
      {stage3_38[5],stage3_37[5],stage3_36[20],stage3_35[28],stage3_34[35]}
   );
   gpc615_5 gpc8885 (
      {stage2_34[85], stage2_34[86], stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[13]},
      {stage2_36[36], stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41]},
      {stage3_38[6],stage3_37[6],stage3_36[21],stage3_35[29],stage3_34[36]}
   );
   gpc615_5 gpc8886 (
      {stage2_34[90], stage2_34[91], stage2_34[92], stage2_34[93], stage2_34[94]},
      {stage2_35[14]},
      {stage2_36[42], stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47]},
      {stage3_38[7],stage3_37[7],stage3_36[22],stage3_35[30],stage3_34[37]}
   );
   gpc615_5 gpc8887 (
      {stage2_34[95], stage2_34[96], stage2_34[97], stage2_34[98], stage2_34[99]},
      {stage2_35[15]},
      {stage2_36[48], stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53]},
      {stage3_38[8],stage3_37[8],stage3_36[23],stage3_35[31],stage3_34[38]}
   );
   gpc615_5 gpc8888 (
      {stage2_34[100], stage2_34[101], stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[16]},
      {stage2_36[54], stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59]},
      {stage3_38[9],stage3_37[9],stage3_36[24],stage3_35[32],stage3_34[39]}
   );
   gpc615_5 gpc8889 (
      {stage2_34[105], stage2_34[106], stage2_34[107], stage2_34[108], stage2_34[109]},
      {stage2_35[17]},
      {stage2_36[60], stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65]},
      {stage3_38[10],stage3_37[10],stage3_36[25],stage3_35[33],stage3_34[40]}
   );
   gpc615_5 gpc8890 (
      {stage2_34[110], stage2_34[111], stage2_34[112], stage2_34[113], stage2_34[114]},
      {stage2_35[18]},
      {stage2_36[66], stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71]},
      {stage3_38[11],stage3_37[11],stage3_36[26],stage3_35[34],stage3_34[41]}
   );
   gpc615_5 gpc8891 (
      {stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118], stage2_34[119]},
      {stage2_35[19]},
      {stage2_36[72], stage2_36[73], stage2_36[74], stage2_36[75], stage2_36[76], stage2_36[77]},
      {stage3_38[12],stage3_37[12],stage3_36[27],stage3_35[35],stage3_34[42]}
   );
   gpc615_5 gpc8892 (
      {stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123], stage2_34[124]},
      {stage2_35[20]},
      {stage2_36[78], stage2_36[79], stage2_36[80], stage2_36[81], stage2_36[82], stage2_36[83]},
      {stage3_38[13],stage3_37[13],stage3_36[28],stage3_35[36],stage3_34[43]}
   );
   gpc615_5 gpc8893 (
      {stage2_34[125], stage2_34[126], stage2_34[127], 1'b0, 1'b0},
      {stage2_35[21]},
      {stage2_36[84], stage2_36[85], stage2_36[86], stage2_36[87], stage2_36[88], stage2_36[89]},
      {stage3_38[14],stage3_37[14],stage3_36[29],stage3_35[37],stage3_34[44]}
   );
   gpc606_5 gpc8894 (
      {stage2_35[22], stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[15],stage3_37[15],stage3_36[30],stage3_35[38]}
   );
   gpc615_5 gpc8895 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[90]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[16],stage3_37[16],stage3_36[31],stage3_35[39]}
   );
   gpc615_5 gpc8896 (
      {stage2_35[33], stage2_35[34], stage2_35[35], stage2_35[36], stage2_35[37]},
      {stage2_36[91]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[17],stage3_37[17],stage3_36[32],stage3_35[40]}
   );
   gpc615_5 gpc8897 (
      {stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41], stage2_35[42]},
      {stage2_36[92]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[18],stage3_37[18],stage3_36[33],stage3_35[41]}
   );
   gpc615_5 gpc8898 (
      {stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[93]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[19],stage3_37[19],stage3_36[34],stage3_35[42]}
   );
   gpc615_5 gpc8899 (
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52]},
      {stage2_36[94]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[20],stage3_37[20],stage3_36[35],stage3_35[43]}
   );
   gpc615_5 gpc8900 (
      {stage2_35[53], stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57]},
      {stage2_36[95]},
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage3_39[6],stage3_38[21],stage3_37[21],stage3_36[36],stage3_35[44]}
   );
   gpc615_5 gpc8901 (
      {stage2_35[58], stage2_35[59], stage2_35[60], stage2_35[61], stage2_35[62]},
      {stage2_36[96]},
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage3_39[7],stage3_38[22],stage3_37[22],stage3_36[37],stage3_35[45]}
   );
   gpc615_5 gpc8902 (
      {stage2_35[63], stage2_35[64], stage2_35[65], stage2_35[66], stage2_35[67]},
      {stage2_36[97]},
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage3_39[8],stage3_38[23],stage3_37[23],stage3_36[38],stage3_35[46]}
   );
   gpc615_5 gpc8903 (
      {stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71], stage2_35[72]},
      {stage2_36[98]},
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58], stage2_37[59]},
      {stage3_39[9],stage3_38[24],stage3_37[24],stage3_36[39],stage3_35[47]}
   );
   gpc615_5 gpc8904 (
      {stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[99]},
      {stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63], stage2_37[64], stage2_37[65]},
      {stage3_39[10],stage3_38[25],stage3_37[25],stage3_36[40],stage3_35[48]}
   );
   gpc615_5 gpc8905 (
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82]},
      {stage2_36[100]},
      {stage2_37[66], stage2_37[67], stage2_37[68], stage2_37[69], stage2_37[70], stage2_37[71]},
      {stage3_39[11],stage3_38[26],stage3_37[26],stage3_36[41],stage3_35[49]}
   );
   gpc615_5 gpc8906 (
      {stage2_35[83], stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87]},
      {stage2_36[101]},
      {stage2_37[72], stage2_37[73], stage2_37[74], stage2_37[75], stage2_37[76], stage2_37[77]},
      {stage3_39[12],stage3_38[27],stage3_37[27],stage3_36[42],stage3_35[50]}
   );
   gpc615_5 gpc8907 (
      {stage2_35[88], stage2_35[89], stage2_35[90], stage2_35[91], stage2_35[92]},
      {stage2_36[102]},
      {stage2_37[78], stage2_37[79], stage2_37[80], stage2_37[81], stage2_37[82], stage2_37[83]},
      {stage3_39[13],stage3_38[28],stage3_37[28],stage3_36[43],stage3_35[51]}
   );
   gpc615_5 gpc8908 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97]},
      {stage2_36[103]},
      {stage2_37[84], stage2_37[85], stage2_37[86], stage2_37[87], stage2_37[88], stage2_37[89]},
      {stage3_39[14],stage3_38[29],stage3_37[29],stage3_36[44],stage3_35[52]}
   );
   gpc615_5 gpc8909 (
      {stage2_35[98], stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102]},
      {stage2_36[104]},
      {stage2_37[90], stage2_37[91], stage2_37[92], stage2_37[93], stage2_37[94], stage2_37[95]},
      {stage3_39[15],stage3_38[30],stage3_37[30],stage3_36[45],stage3_35[53]}
   );
   gpc615_5 gpc8910 (
      {stage2_35[103], stage2_35[104], stage2_35[105], stage2_35[106], stage2_35[107]},
      {stage2_36[105]},
      {stage2_37[96], stage2_37[97], stage2_37[98], stage2_37[99], stage2_37[100], stage2_37[101]},
      {stage3_39[16],stage3_38[31],stage3_37[31],stage3_36[46],stage3_35[54]}
   );
   gpc615_5 gpc8911 (
      {stage2_35[108], stage2_35[109], stage2_35[110], stage2_35[111], stage2_35[112]},
      {stage2_36[106]},
      {stage2_37[102], stage2_37[103], stage2_37[104], stage2_37[105], stage2_37[106], stage2_37[107]},
      {stage3_39[17],stage3_38[32],stage3_37[32],stage3_36[47],stage3_35[55]}
   );
   gpc615_5 gpc8912 (
      {stage2_35[113], stage2_35[114], stage2_35[115], stage2_35[116], stage2_35[117]},
      {stage2_36[107]},
      {stage2_37[108], stage2_37[109], stage2_37[110], stage2_37[111], stage2_37[112], stage2_37[113]},
      {stage3_39[18],stage3_38[33],stage3_37[33],stage3_36[48],stage3_35[56]}
   );
   gpc606_5 gpc8913 (
      {stage2_36[108], stage2_36[109], stage2_36[110], stage2_36[111], stage2_36[112], stage2_36[113]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[19],stage3_38[34],stage3_37[34],stage3_36[49]}
   );
   gpc615_5 gpc8914 (
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10]},
      {stage2_39[0]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[1],stage3_39[20],stage3_38[35]}
   );
   gpc615_5 gpc8915 (
      {stage2_38[11], stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15]},
      {stage2_39[1]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[1],stage3_40[2],stage3_39[21],stage3_38[36]}
   );
   gpc615_5 gpc8916 (
      {stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_39[2]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[2],stage3_40[3],stage3_39[22],stage3_38[37]}
   );
   gpc615_5 gpc8917 (
      {stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage2_39[3]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[3],stage3_40[4],stage3_39[23],stage3_38[38]}
   );
   gpc615_5 gpc8918 (
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30]},
      {stage2_39[4]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[4],stage3_40[5],stage3_39[24],stage3_38[39]}
   );
   gpc615_5 gpc8919 (
      {stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage2_39[5]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[5],stage3_40[6],stage3_39[25],stage3_38[40]}
   );
   gpc615_5 gpc8920 (
      {stage2_38[36], stage2_38[37], stage2_38[38], stage2_38[39], stage2_38[40]},
      {stage2_39[6]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[6],stage3_40[7],stage3_39[26],stage3_38[41]}
   );
   gpc615_5 gpc8921 (
      {stage2_38[41], stage2_38[42], stage2_38[43], stage2_38[44], stage2_38[45]},
      {stage2_39[7]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[7],stage3_40[8],stage3_39[27],stage3_38[42]}
   );
   gpc615_5 gpc8922 (
      {stage2_38[46], stage2_38[47], stage2_38[48], stage2_38[49], stage2_38[50]},
      {stage2_39[8]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[8],stage3_40[9],stage3_39[28],stage3_38[43]}
   );
   gpc615_5 gpc8923 (
      {stage2_38[51], stage2_38[52], stage2_38[53], stage2_38[54], stage2_38[55]},
      {stage2_39[9]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[9],stage3_40[10],stage3_39[29],stage3_38[44]}
   );
   gpc615_5 gpc8924 (
      {stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59], stage2_38[60]},
      {stage2_39[10]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[10],stage3_40[11],stage3_39[30],stage3_38[45]}
   );
   gpc615_5 gpc8925 (
      {stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_39[11]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[11],stage3_40[12],stage3_39[31],stage3_38[46]}
   );
   gpc615_5 gpc8926 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70]},
      {stage2_39[12]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[12],stage3_40[13],stage3_39[32],stage3_38[47]}
   );
   gpc615_5 gpc8927 (
      {stage2_38[71], stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75]},
      {stage2_39[13]},
      {stage2_40[78], stage2_40[79], stage2_40[80], stage2_40[81], stage2_40[82], stage2_40[83]},
      {stage3_42[13],stage3_41[13],stage3_40[14],stage3_39[33],stage3_38[48]}
   );
   gpc615_5 gpc8928 (
      {stage2_38[76], stage2_38[77], stage2_38[78], stage2_38[79], stage2_38[80]},
      {stage2_39[14]},
      {stage2_40[84], stage2_40[85], stage2_40[86], stage2_40[87], stage2_40[88], stage2_40[89]},
      {stage3_42[14],stage3_41[14],stage3_40[15],stage3_39[34],stage3_38[49]}
   );
   gpc615_5 gpc8929 (
      {stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_40[90]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[15],stage3_41[15],stage3_40[16],stage3_39[35]}
   );
   gpc615_5 gpc8930 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24]},
      {stage2_40[91]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[16],stage3_41[16],stage3_40[17],stage3_39[36]}
   );
   gpc615_5 gpc8931 (
      {stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage2_40[92]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[17],stage3_41[17],stage3_40[18],stage3_39[37]}
   );
   gpc615_5 gpc8932 (
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34]},
      {stage2_40[93]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[18],stage3_41[18],stage3_40[19],stage3_39[38]}
   );
   gpc615_5 gpc8933 (
      {stage2_39[35], stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39]},
      {stage2_40[94]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[19],stage3_41[19],stage3_40[20],stage3_39[39]}
   );
   gpc615_5 gpc8934 (
      {stage2_39[40], stage2_39[41], stage2_39[42], stage2_39[43], stage2_39[44]},
      {stage2_40[95]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[20],stage3_41[20],stage3_40[21],stage3_39[40]}
   );
   gpc615_5 gpc8935 (
      {stage2_39[45], stage2_39[46], stage2_39[47], stage2_39[48], stage2_39[49]},
      {stage2_40[96]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[21],stage3_41[21],stage3_40[22],stage3_39[41]}
   );
   gpc615_5 gpc8936 (
      {stage2_39[50], stage2_39[51], stage2_39[52], stage2_39[53], stage2_39[54]},
      {stage2_40[97]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[22],stage3_41[22],stage3_40[23],stage3_39[42]}
   );
   gpc615_5 gpc8937 (
      {stage2_39[55], stage2_39[56], stage2_39[57], stage2_39[58], stage2_39[59]},
      {stage2_40[98]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[23],stage3_41[23],stage3_40[24],stage3_39[43]}
   );
   gpc615_5 gpc8938 (
      {stage2_39[60], stage2_39[61], stage2_39[62], stage2_39[63], stage2_39[64]},
      {stage2_40[99]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[24],stage3_41[24],stage3_40[25],stage3_39[44]}
   );
   gpc615_5 gpc8939 (
      {stage2_39[65], stage2_39[66], stage2_39[67], stage2_39[68], stage2_39[69]},
      {stage2_40[100]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[25],stage3_41[25],stage3_40[26],stage3_39[45]}
   );
   gpc615_5 gpc8940 (
      {stage2_39[70], stage2_39[71], stage2_39[72], stage2_39[73], stage2_39[74]},
      {stage2_40[101]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[26],stage3_41[26],stage3_40[27],stage3_39[46]}
   );
   gpc615_5 gpc8941 (
      {stage2_39[75], stage2_39[76], stage2_39[77], stage2_39[78], stage2_39[79]},
      {stage2_40[102]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[27],stage3_41[27],stage3_40[28],stage3_39[47]}
   );
   gpc615_5 gpc8942 (
      {stage2_39[80], stage2_39[81], stage2_39[82], stage2_39[83], stage2_39[84]},
      {stage2_40[103]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[28],stage3_41[28],stage3_40[29],stage3_39[48]}
   );
   gpc615_5 gpc8943 (
      {stage2_39[85], stage2_39[86], stage2_39[87], stage2_39[88], stage2_39[89]},
      {stage2_40[104]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[29],stage3_41[29],stage3_40[30],stage3_39[49]}
   );
   gpc615_5 gpc8944 (
      {stage2_39[90], stage2_39[91], stage2_39[92], stage2_39[93], stage2_39[94]},
      {stage2_40[105]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[30],stage3_41[30],stage3_40[31],stage3_39[50]}
   );
   gpc615_5 gpc8945 (
      {stage2_39[95], stage2_39[96], stage2_39[97], stage2_39[98], stage2_39[99]},
      {stage2_40[106]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[31],stage3_41[31],stage3_40[32],stage3_39[51]}
   );
   gpc606_5 gpc8946 (
      {stage2_40[107], stage2_40[108], stage2_40[109], stage2_40[110], stage2_40[111], stage2_40[112]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[32],stage3_41[32],stage3_40[33]}
   );
   gpc606_5 gpc8947 (
      {stage2_40[113], stage2_40[114], stage2_40[115], stage2_40[116], stage2_40[117], stage2_40[118]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[33],stage3_41[33],stage3_40[34]}
   );
   gpc606_5 gpc8948 (
      {stage2_40[119], stage2_40[120], stage2_40[121], stage2_40[122], stage2_40[123], stage2_40[124]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[19],stage3_42[34],stage3_41[34],stage3_40[35]}
   );
   gpc606_5 gpc8949 (
      {stage2_40[125], stage2_40[126], stage2_40[127], stage2_40[128], stage2_40[129], stage2_40[130]},
      {stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21], stage2_42[22], stage2_42[23]},
      {stage3_44[3],stage3_43[20],stage3_42[35],stage3_41[35],stage3_40[36]}
   );
   gpc615_5 gpc8950 (
      {stage2_42[24], stage2_42[25], stage2_42[26], stage2_42[27], stage2_42[28]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[21],stage3_42[36]}
   );
   gpc615_5 gpc8951 (
      {stage2_42[29], stage2_42[30], stage2_42[31], stage2_42[32], stage2_42[33]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[22],stage3_42[37]}
   );
   gpc615_5 gpc8952 (
      {stage2_42[34], stage2_42[35], stage2_42[36], stage2_42[37], stage2_42[38]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[6],stage3_43[23],stage3_42[38]}
   );
   gpc615_5 gpc8953 (
      {stage2_42[39], stage2_42[40], stage2_42[41], stage2_42[42], stage2_42[43]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[7],stage3_43[24],stage3_42[39]}
   );
   gpc615_5 gpc8954 (
      {stage2_42[44], stage2_42[45], stage2_42[46], stage2_42[47], stage2_42[48]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[8],stage3_43[25],stage3_42[40]}
   );
   gpc615_5 gpc8955 (
      {stage2_42[49], stage2_42[50], stage2_42[51], stage2_42[52], stage2_42[53]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[9],stage3_43[26],stage3_42[41]}
   );
   gpc615_5 gpc8956 (
      {stage2_42[54], stage2_42[55], stage2_42[56], stage2_42[57], stage2_42[58]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[10],stage3_43[27],stage3_42[42]}
   );
   gpc615_5 gpc8957 (
      {stage2_42[59], stage2_42[60], stage2_42[61], stage2_42[62], stage2_42[63]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[11],stage3_43[28],stage3_42[43]}
   );
   gpc615_5 gpc8958 (
      {stage2_42[64], stage2_42[65], stage2_42[66], stage2_42[67], stage2_42[68]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[12],stage3_43[29],stage3_42[44]}
   );
   gpc615_5 gpc8959 (
      {stage2_42[69], stage2_42[70], stage2_42[71], stage2_42[72], stage2_42[73]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[13],stage3_43[30],stage3_42[45]}
   );
   gpc606_5 gpc8960 (
      {stage2_43[10], stage2_43[11], stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[10],stage3_45[10],stage3_44[14],stage3_43[31]}
   );
   gpc606_5 gpc8961 (
      {stage2_43[16], stage2_43[17], stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[11],stage3_45[11],stage3_44[15],stage3_43[32]}
   );
   gpc606_5 gpc8962 (
      {stage2_43[22], stage2_43[23], stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[12],stage3_45[12],stage3_44[16],stage3_43[33]}
   );
   gpc606_5 gpc8963 (
      {stage2_43[28], stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[13],stage3_45[13],stage3_44[17],stage3_43[34]}
   );
   gpc606_5 gpc8964 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38], stage2_43[39]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[14],stage3_45[14],stage3_44[18],stage3_43[35]}
   );
   gpc606_5 gpc8965 (
      {stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[15],stage3_45[15],stage3_44[19],stage3_43[36]}
   );
   gpc606_5 gpc8966 (
      {stage2_43[46], stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[16],stage3_45[16],stage3_44[20],stage3_43[37]}
   );
   gpc606_5 gpc8967 (
      {stage2_43[52], stage2_43[53], stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[17],stage3_45[17],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc8968 (
      {stage2_43[58], stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62]},
      {stage2_44[60]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[18],stage3_45[18],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc8969 (
      {stage2_43[63], stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67]},
      {stage2_44[61]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[19],stage3_45[19],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc8970 (
      {stage2_43[68], stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72]},
      {stage2_44[62]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[20],stage3_45[20],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc8971 (
      {stage2_43[73], stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77]},
      {stage2_44[63]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[21],stage3_45[21],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc8972 (
      {stage2_43[78], stage2_43[79], stage2_43[80], stage2_43[81], stage2_43[82]},
      {stage2_44[64]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[22],stage3_45[22],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc8973 (
      {stage2_43[83], stage2_43[84], stage2_43[85], stage2_43[86], stage2_43[87]},
      {stage2_44[65]},
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage3_47[13],stage3_46[23],stage3_45[23],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc8974 (
      {stage2_43[88], stage2_43[89], stage2_43[90], stage2_43[91], stage2_43[92]},
      {stage2_44[66]},
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage3_47[14],stage3_46[24],stage3_45[24],stage3_44[28],stage3_43[45]}
   );
   gpc615_5 gpc8975 (
      {stage2_43[93], stage2_43[94], stage2_43[95], stage2_43[96], stage2_43[97]},
      {stage2_44[67]},
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage3_47[15],stage3_46[25],stage3_45[25],stage3_44[29],stage3_43[46]}
   );
   gpc606_5 gpc8976 (
      {stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71], stage2_44[72], stage2_44[73]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[16],stage3_46[26],stage3_45[26],stage3_44[30]}
   );
   gpc606_5 gpc8977 (
      {stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77], stage2_44[78], stage2_44[79]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[17],stage3_46[27],stage3_45[27],stage3_44[31]}
   );
   gpc606_5 gpc8978 (
      {stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83], stage2_44[84], stage2_44[85]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[18],stage3_46[28],stage3_45[28],stage3_44[32]}
   );
   gpc606_5 gpc8979 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[3],stage3_47[19],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc8980 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[4],stage3_47[20],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc8981 (
      {stage2_45[108], stage2_45[109], stage2_45[110], stage2_45[111], stage2_45[112], stage2_45[113]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[5],stage3_47[21],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc8982 (
      {stage2_45[114], stage2_45[115], stage2_45[116], stage2_45[117], stage2_45[118], stage2_45[119]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[6],stage3_47[22],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc8983 (
      {stage2_45[120], stage2_45[121], stage2_45[122], stage2_45[123], stage2_45[124], stage2_45[125]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[7],stage3_47[23],stage3_46[33],stage3_45[33]}
   );
   gpc615_5 gpc8984 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[30]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[5],stage3_48[8],stage3_47[24],stage3_46[34]}
   );
   gpc615_5 gpc8985 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[31]},
      {stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage3_50[1],stage3_49[6],stage3_48[9],stage3_47[25],stage3_46[35]}
   );
   gpc615_5 gpc8986 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[32]},
      {stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17]},
      {stage3_50[2],stage3_49[7],stage3_48[10],stage3_47[26],stage3_46[36]}
   );
   gpc615_5 gpc8987 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[33]},
      {stage2_48[18], stage2_48[19], stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23]},
      {stage3_50[3],stage3_49[8],stage3_48[11],stage3_47[27],stage3_46[37]}
   );
   gpc615_5 gpc8988 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[34]},
      {stage2_48[24], stage2_48[25], stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29]},
      {stage3_50[4],stage3_49[9],stage3_48[12],stage3_47[28],stage3_46[38]}
   );
   gpc615_5 gpc8989 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[35]},
      {stage2_48[30], stage2_48[31], stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35]},
      {stage3_50[5],stage3_49[10],stage3_48[13],stage3_47[29],stage3_46[39]}
   );
   gpc615_5 gpc8990 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[36]},
      {stage2_48[36], stage2_48[37], stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41]},
      {stage3_50[6],stage3_49[11],stage3_48[14],stage3_47[30],stage3_46[40]}
   );
   gpc615_5 gpc8991 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[37]},
      {stage2_48[42], stage2_48[43], stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47]},
      {stage3_50[7],stage3_49[12],stage3_48[15],stage3_47[31],stage3_46[41]}
   );
   gpc615_5 gpc8992 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[38]},
      {stage2_48[48], stage2_48[49], stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53]},
      {stage3_50[8],stage3_49[13],stage3_48[16],stage3_47[32],stage3_46[42]}
   );
   gpc615_5 gpc8993 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[39]},
      {stage2_48[54], stage2_48[55], stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59]},
      {stage3_50[9],stage3_49[14],stage3_48[17],stage3_47[33],stage3_46[43]}
   );
   gpc615_5 gpc8994 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[40]},
      {stage2_48[60], stage2_48[61], stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65]},
      {stage3_50[10],stage3_49[15],stage3_48[18],stage3_47[34],stage3_46[44]}
   );
   gpc615_5 gpc8995 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[41]},
      {stage2_48[66], stage2_48[67], stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71]},
      {stage3_50[11],stage3_49[16],stage3_48[19],stage3_47[35],stage3_46[45]}
   );
   gpc615_5 gpc8996 (
      {stage2_46[78], stage2_46[79], stage2_46[80], stage2_46[81], stage2_46[82]},
      {stage2_47[42]},
      {stage2_48[72], stage2_48[73], stage2_48[74], stage2_48[75], stage2_48[76], stage2_48[77]},
      {stage3_50[12],stage3_49[17],stage3_48[20],stage3_47[36],stage3_46[46]}
   );
   gpc615_5 gpc8997 (
      {stage2_46[83], stage2_46[84], stage2_46[85], stage2_46[86], stage2_46[87]},
      {stage2_47[43]},
      {stage2_48[78], stage2_48[79], stage2_48[80], stage2_48[81], stage2_48[82], stage2_48[83]},
      {stage3_50[13],stage3_49[18],stage3_48[21],stage3_47[37],stage3_46[47]}
   );
   gpc615_5 gpc8998 (
      {stage2_46[88], stage2_46[89], stage2_46[90], stage2_46[91], stage2_46[92]},
      {stage2_47[44]},
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage3_50[14],stage3_49[19],stage3_48[22],stage3_47[38],stage3_46[48]}
   );
   gpc1163_5 gpc8999 (
      {stage2_47[45], stage2_47[46], stage2_47[47]},
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_49[0]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[15],stage3_49[20],stage3_48[23],stage3_47[39]}
   );
   gpc1163_5 gpc9000 (
      {stage2_47[48], stage2_47[49], stage2_47[50]},
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_49[1]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[16],stage3_49[21],stage3_48[24],stage3_47[40]}
   );
   gpc1163_5 gpc9001 (
      {stage2_47[51], stage2_47[52], stage2_47[53]},
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_49[2]},
      {stage2_50[2]},
      {stage3_51[2],stage3_50[17],stage3_49[22],stage3_48[25],stage3_47[41]}
   );
   gpc1163_5 gpc9002 (
      {stage2_47[54], stage2_47[55], stage2_47[56]},
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_49[3]},
      {stage2_50[3]},
      {stage3_51[3],stage3_50[18],stage3_49[23],stage3_48[26],stage3_47[42]}
   );
   gpc1163_5 gpc9003 (
      {stage2_47[57], stage2_47[58], stage2_47[59]},
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_49[4]},
      {stage2_50[4]},
      {stage3_51[4],stage3_50[19],stage3_49[24],stage3_48[27],stage3_47[43]}
   );
   gpc1163_5 gpc9004 (
      {stage2_47[60], stage2_47[61], stage2_47[62]},
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_49[5]},
      {stage2_50[5]},
      {stage3_51[5],stage3_50[20],stage3_49[25],stage3_48[28],stage3_47[44]}
   );
   gpc615_5 gpc9005 (
      {stage2_47[63], stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67]},
      {stage2_48[126]},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[6],stage3_50[21],stage3_49[26],stage3_48[29],stage3_47[45]}
   );
   gpc615_5 gpc9006 (
      {stage2_47[68], stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72]},
      {stage2_48[127]},
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage3_51[7],stage3_50[22],stage3_49[27],stage3_48[30],stage3_47[46]}
   );
   gpc615_5 gpc9007 (
      {stage2_47[73], stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77]},
      {stage2_48[128]},
      {stage2_49[18], stage2_49[19], stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23]},
      {stage3_51[8],stage3_50[23],stage3_49[28],stage3_48[31],stage3_47[47]}
   );
   gpc615_5 gpc9008 (
      {stage2_47[78], stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82]},
      {stage2_48[129]},
      {stage2_49[24], stage2_49[25], stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29]},
      {stage3_51[9],stage3_50[24],stage3_49[29],stage3_48[32],stage3_47[48]}
   );
   gpc606_5 gpc9009 (
      {stage2_48[130], stage2_48[131], stage2_48[132], stage2_48[133], stage2_48[134], stage2_48[135]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[0],stage3_51[10],stage3_50[25],stage3_49[30],stage3_48[33]}
   );
   gpc606_5 gpc9010 (
      {stage2_48[136], stage2_48[137], stage2_48[138], stage2_48[139], stage2_48[140], stage2_48[141]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[1],stage3_51[11],stage3_50[26],stage3_49[31],stage3_48[34]}
   );
   gpc606_5 gpc9011 (
      {stage2_48[142], stage2_48[143], stage2_48[144], stage2_48[145], stage2_48[146], stage2_48[147]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[2],stage3_51[12],stage3_50[27],stage3_49[32],stage3_48[35]}
   );
   gpc606_5 gpc9012 (
      {stage2_48[148], stage2_48[149], stage2_48[150], stage2_48[151], stage2_48[152], stage2_48[153]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[3],stage3_51[13],stage3_50[28],stage3_49[33],stage3_48[36]}
   );
   gpc606_5 gpc9013 (
      {stage2_49[30], stage2_49[31], stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[4],stage3_51[14],stage3_50[29],stage3_49[34]}
   );
   gpc606_5 gpc9014 (
      {stage2_49[36], stage2_49[37], stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[5],stage3_51[15],stage3_50[30],stage3_49[35]}
   );
   gpc606_5 gpc9015 (
      {stage2_49[42], stage2_49[43], stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[6],stage3_51[16],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc9016 (
      {stage2_49[48], stage2_49[49], stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[7],stage3_51[17],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc9017 (
      {stage2_49[54], stage2_49[55], stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[8],stage3_51[18],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc9018 (
      {stage2_49[60], stage2_49[61], stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[9],stage3_51[19],stage3_50[34],stage3_49[39]}
   );
   gpc606_5 gpc9019 (
      {stage2_49[66], stage2_49[67], stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71]},
      {stage2_51[36], stage2_51[37], stage2_51[38], stage2_51[39], stage2_51[40], stage2_51[41]},
      {stage3_53[6],stage3_52[10],stage3_51[20],stage3_50[35],stage3_49[40]}
   );
   gpc606_5 gpc9020 (
      {stage2_49[72], stage2_49[73], stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77]},
      {stage2_51[42], stage2_51[43], stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47]},
      {stage3_53[7],stage3_52[11],stage3_51[21],stage3_50[36],stage3_49[41]}
   );
   gpc606_5 gpc9021 (
      {stage2_49[78], stage2_49[79], stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83]},
      {stage2_51[48], stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage3_53[8],stage3_52[12],stage3_51[22],stage3_50[37],stage3_49[42]}
   );
   gpc606_5 gpc9022 (
      {stage2_49[84], stage2_49[85], stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89]},
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58], stage2_51[59]},
      {stage3_53[9],stage3_52[13],stage3_51[23],stage3_50[38],stage3_49[43]}
   );
   gpc606_5 gpc9023 (
      {stage2_49[90], stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_51[60], stage2_51[61], stage2_51[62], stage2_51[63], stage2_51[64], stage2_51[65]},
      {stage3_53[10],stage3_52[14],stage3_51[24],stage3_50[39],stage3_49[44]}
   );
   gpc2135_5 gpc9024 (
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34]},
      {stage2_51[66], stage2_51[67], stage2_51[68]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[11],stage3_52[15],stage3_51[25],stage3_50[40]}
   );
   gpc1406_5 gpc9025 (
      {stage2_50[35], stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40]},
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4]},
      {stage2_53[2]},
      {stage3_54[1],stage3_53[12],stage3_52[16],stage3_51[26],stage3_50[41]}
   );
   gpc1406_5 gpc9026 (
      {stage2_50[41], stage2_50[42], stage2_50[43], stage2_50[44], stage2_50[45], stage2_50[46]},
      {stage2_52[5], stage2_52[6], stage2_52[7], stage2_52[8]},
      {stage2_53[3]},
      {stage3_54[2],stage3_53[13],stage3_52[17],stage3_51[27],stage3_50[42]}
   );
   gpc1406_5 gpc9027 (
      {stage2_50[47], stage2_50[48], stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52]},
      {stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12]},
      {stage2_53[4]},
      {stage3_54[3],stage3_53[14],stage3_52[18],stage3_51[28],stage3_50[43]}
   );
   gpc606_5 gpc9028 (
      {stage2_50[53], stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17], stage2_52[18]},
      {stage3_54[4],stage3_53[15],stage3_52[19],stage3_51[29],stage3_50[44]}
   );
   gpc606_5 gpc9029 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63], stage2_50[64]},
      {stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23], stage2_52[24]},
      {stage3_54[5],stage3_53[16],stage3_52[20],stage3_51[30],stage3_50[45]}
   );
   gpc606_5 gpc9030 (
      {stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68], stage2_50[69], stage2_50[70]},
      {stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29], stage2_52[30]},
      {stage3_54[6],stage3_53[17],stage3_52[21],stage3_51[31],stage3_50[46]}
   );
   gpc606_5 gpc9031 (
      {stage2_50[71], stage2_50[72], stage2_50[73], stage2_50[74], stage2_50[75], stage2_50[76]},
      {stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35], stage2_52[36]},
      {stage3_54[7],stage3_53[18],stage3_52[22],stage3_51[32],stage3_50[47]}
   );
   gpc606_5 gpc9032 (
      {stage2_50[77], stage2_50[78], stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82]},
      {stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41], stage2_52[42]},
      {stage3_54[8],stage3_53[19],stage3_52[23],stage3_51[33],stage3_50[48]}
   );
   gpc606_5 gpc9033 (
      {stage2_50[83], stage2_50[84], stage2_50[85], stage2_50[86], stage2_50[87], stage2_50[88]},
      {stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47], stage2_52[48]},
      {stage3_54[9],stage3_53[20],stage3_52[24],stage3_51[34],stage3_50[49]}
   );
   gpc606_5 gpc9034 (
      {stage2_50[89], stage2_50[90], stage2_50[91], stage2_50[92], stage2_50[93], stage2_50[94]},
      {stage2_52[49], stage2_52[50], stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54]},
      {stage3_54[10],stage3_53[21],stage3_52[25],stage3_51[35],stage3_50[50]}
   );
   gpc606_5 gpc9035 (
      {stage2_50[95], stage2_50[96], stage2_50[97], stage2_50[98], stage2_50[99], stage2_50[100]},
      {stage2_52[55], stage2_52[56], stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60]},
      {stage3_54[11],stage3_53[22],stage3_52[26],stage3_51[36],stage3_50[51]}
   );
   gpc606_5 gpc9036 (
      {stage2_50[101], stage2_50[102], stage2_50[103], stage2_50[104], stage2_50[105], stage2_50[106]},
      {stage2_52[61], stage2_52[62], stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66]},
      {stage3_54[12],stage3_53[23],stage3_52[27],stage3_51[37],stage3_50[52]}
   );
   gpc606_5 gpc9037 (
      {stage2_50[107], stage2_50[108], stage2_50[109], stage2_50[110], stage2_50[111], stage2_50[112]},
      {stage2_52[67], stage2_52[68], stage2_52[69], stage2_52[70], stage2_52[71], stage2_52[72]},
      {stage3_54[13],stage3_53[24],stage3_52[28],stage3_51[38],stage3_50[53]}
   );
   gpc606_5 gpc9038 (
      {stage2_50[113], stage2_50[114], stage2_50[115], stage2_50[116], stage2_50[117], stage2_50[118]},
      {stage2_52[73], stage2_52[74], stage2_52[75], stage2_52[76], stage2_52[77], stage2_52[78]},
      {stage3_54[14],stage3_53[25],stage3_52[29],stage3_51[39],stage3_50[54]}
   );
   gpc606_5 gpc9039 (
      {stage2_50[119], stage2_50[120], stage2_50[121], stage2_50[122], stage2_50[123], stage2_50[124]},
      {stage2_52[79], stage2_52[80], stage2_52[81], stage2_52[82], stage2_52[83], stage2_52[84]},
      {stage3_54[15],stage3_53[26],stage3_52[30],stage3_51[40],stage3_50[55]}
   );
   gpc606_5 gpc9040 (
      {stage2_50[125], stage2_50[126], stage2_50[127], stage2_50[128], stage2_50[129], stage2_50[130]},
      {stage2_52[85], stage2_52[86], stage2_52[87], stage2_52[88], stage2_52[89], stage2_52[90]},
      {stage3_54[16],stage3_53[27],stage3_52[31],stage3_51[41],stage3_50[56]}
   );
   gpc606_5 gpc9041 (
      {stage2_50[131], stage2_50[132], stage2_50[133], stage2_50[134], stage2_50[135], stage2_50[136]},
      {stage2_52[91], stage2_52[92], stage2_52[93], stage2_52[94], stage2_52[95], stage2_52[96]},
      {stage3_54[17],stage3_53[28],stage3_52[32],stage3_51[42],stage3_50[57]}
   );
   gpc606_5 gpc9042 (
      {stage2_50[137], stage2_50[138], stage2_50[139], stage2_50[140], stage2_50[141], stage2_50[142]},
      {stage2_52[97], stage2_52[98], stage2_52[99], stage2_52[100], stage2_52[101], stage2_52[102]},
      {stage3_54[18],stage3_53[29],stage3_52[33],stage3_51[43],stage3_50[58]}
   );
   gpc606_5 gpc9043 (
      {stage2_50[143], stage2_50[144], stage2_50[145], stage2_50[146], stage2_50[147], stage2_50[148]},
      {stage2_52[103], stage2_52[104], stage2_52[105], stage2_52[106], stage2_52[107], stage2_52[108]},
      {stage3_54[19],stage3_53[30],stage3_52[34],stage3_51[44],stage3_50[59]}
   );
   gpc606_5 gpc9044 (
      {stage2_51[69], stage2_51[70], stage2_51[71], stage2_51[72], stage2_51[73], stage2_51[74]},
      {stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10]},
      {stage3_55[0],stage3_54[20],stage3_53[31],stage3_52[35],stage3_51[45]}
   );
   gpc606_5 gpc9045 (
      {stage2_51[75], stage2_51[76], stage2_51[77], stage2_51[78], stage2_51[79], stage2_51[80]},
      {stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16]},
      {stage3_55[1],stage3_54[21],stage3_53[32],stage3_52[36],stage3_51[46]}
   );
   gpc606_5 gpc9046 (
      {stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[2],stage3_54[22],stage3_53[33]}
   );
   gpc606_5 gpc9047 (
      {stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[3],stage3_54[23],stage3_53[34]}
   );
   gpc606_5 gpc9048 (
      {stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[4],stage3_54[24],stage3_53[35]}
   );
   gpc606_5 gpc9049 (
      {stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[3],stage3_55[5],stage3_54[25],stage3_53[36]}
   );
   gpc606_5 gpc9050 (
      {stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[4],stage3_55[6],stage3_54[26],stage3_53[37]}
   );
   gpc606_5 gpc9051 (
      {stage2_53[47], stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[5],stage3_55[7],stage3_54[27],stage3_53[38]}
   );
   gpc606_5 gpc9052 (
      {stage2_53[53], stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[6],stage3_55[8],stage3_54[28],stage3_53[39]}
   );
   gpc606_5 gpc9053 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63], stage2_53[64]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[7],stage3_55[9],stage3_54[29],stage3_53[40]}
   );
   gpc606_5 gpc9054 (
      {stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68], stage2_53[69], stage2_53[70]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[8],stage3_55[10],stage3_54[30],stage3_53[41]}
   );
   gpc606_5 gpc9055 (
      {stage2_53[71], stage2_53[72], stage2_53[73], stage2_53[74], stage2_53[75], stage2_53[76]},
      {stage2_55[54], stage2_55[55], stage2_55[56], stage2_55[57], stage2_55[58], stage2_55[59]},
      {stage3_57[9],stage3_56[9],stage3_55[11],stage3_54[31],stage3_53[42]}
   );
   gpc606_5 gpc9056 (
      {stage2_53[77], stage2_53[78], stage2_53[79], stage2_53[80], stage2_53[81], stage2_53[82]},
      {stage2_55[60], stage2_55[61], stage2_55[62], stage2_55[63], stage2_55[64], stage2_55[65]},
      {stage3_57[10],stage3_56[10],stage3_55[12],stage3_54[32],stage3_53[43]}
   );
   gpc606_5 gpc9057 (
      {stage2_53[83], stage2_53[84], stage2_53[85], stage2_53[86], stage2_53[87], stage2_53[88]},
      {stage2_55[66], stage2_55[67], stage2_55[68], stage2_55[69], stage2_55[70], stage2_55[71]},
      {stage3_57[11],stage3_56[11],stage3_55[13],stage3_54[33],stage3_53[44]}
   );
   gpc606_5 gpc9058 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[12],stage3_56[12],stage3_55[14],stage3_54[34]}
   );
   gpc606_5 gpc9059 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[13],stage3_56[13],stage3_55[15],stage3_54[35]}
   );
   gpc606_5 gpc9060 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[14],stage3_56[14],stage3_55[16],stage3_54[36]}
   );
   gpc606_5 gpc9061 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22], stage2_54[23]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[15],stage3_56[15],stage3_55[17],stage3_54[37]}
   );
   gpc606_5 gpc9062 (
      {stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[16],stage3_56[16],stage3_55[18],stage3_54[38]}
   );
   gpc606_5 gpc9063 (
      {stage2_54[30], stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[17],stage3_56[17],stage3_55[19],stage3_54[39]}
   );
   gpc606_5 gpc9064 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40], stage2_54[41]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[18],stage3_56[18],stage3_55[20],stage3_54[40]}
   );
   gpc606_5 gpc9065 (
      {stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45], stage2_54[46], stage2_54[47]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[19],stage3_56[19],stage3_55[21],stage3_54[41]}
   );
   gpc606_5 gpc9066 (
      {stage2_54[48], stage2_54[49], stage2_54[50], stage2_54[51], stage2_54[52], stage2_54[53]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[20],stage3_56[20],stage3_55[22],stage3_54[42]}
   );
   gpc606_5 gpc9067 (
      {stage2_54[54], stage2_54[55], stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[21],stage3_56[21],stage3_55[23],stage3_54[43]}
   );
   gpc606_5 gpc9068 (
      {stage2_54[60], stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[22],stage3_56[22],stage3_55[24],stage3_54[44]}
   );
   gpc606_5 gpc9069 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70], stage2_54[71]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[23],stage3_56[23],stage3_55[25],stage3_54[45]}
   );
   gpc606_5 gpc9070 (
      {stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75], stage2_54[76], stage2_54[77]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[24],stage3_56[24],stage3_55[26],stage3_54[46]}
   );
   gpc606_5 gpc9071 (
      {stage2_54[78], stage2_54[79], stage2_54[80], stage2_54[81], stage2_54[82], stage2_54[83]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[25],stage3_56[25],stage3_55[27],stage3_54[47]}
   );
   gpc606_5 gpc9072 (
      {stage2_54[84], stage2_54[85], stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[26],stage3_56[26],stage3_55[28],stage3_54[48]}
   );
   gpc606_5 gpc9073 (
      {stage2_54[90], stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[27],stage3_56[27],stage3_55[29],stage3_54[49]}
   );
   gpc606_5 gpc9074 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], stage2_54[100], stage2_54[101]},
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100], stage2_56[101]},
      {stage3_58[16],stage3_57[28],stage3_56[28],stage3_55[30],stage3_54[50]}
   );
   gpc606_5 gpc9075 (
      {stage2_54[102], stage2_54[103], stage2_54[104], stage2_54[105], stage2_54[106], stage2_54[107]},
      {stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105], stage2_56[106], stage2_56[107]},
      {stage3_58[17],stage3_57[29],stage3_56[29],stage3_55[31],stage3_54[51]}
   );
   gpc606_5 gpc9076 (
      {stage2_54[108], stage2_54[109], stage2_54[110], stage2_54[111], stage2_54[112], stage2_54[113]},
      {stage2_56[108], stage2_56[109], stage2_56[110], stage2_56[111], stage2_56[112], stage2_56[113]},
      {stage3_58[18],stage3_57[30],stage3_56[30],stage3_55[32],stage3_54[52]}
   );
   gpc606_5 gpc9077 (
      {stage2_55[72], stage2_55[73], stage2_55[74], stage2_55[75], stage2_55[76], stage2_55[77]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[19],stage3_57[31],stage3_56[31],stage3_55[33]}
   );
   gpc606_5 gpc9078 (
      {stage2_55[78], stage2_55[79], stage2_55[80], stage2_55[81], stage2_55[82], stage2_55[83]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[20],stage3_57[32],stage3_56[32],stage3_55[34]}
   );
   gpc606_5 gpc9079 (
      {stage2_55[84], stage2_55[85], stage2_55[86], stage2_55[87], stage2_55[88], stage2_55[89]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[21],stage3_57[33],stage3_56[33],stage3_55[35]}
   );
   gpc606_5 gpc9080 (
      {stage2_55[90], stage2_55[91], stage2_55[92], stage2_55[93], stage2_55[94], stage2_55[95]},
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage3_59[3],stage3_58[22],stage3_57[34],stage3_56[34],stage3_55[36]}
   );
   gpc606_5 gpc9081 (
      {stage2_55[96], stage2_55[97], stage2_55[98], stage2_55[99], stage2_55[100], stage2_55[101]},
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage3_59[4],stage3_58[23],stage3_57[35],stage3_56[35],stage3_55[37]}
   );
   gpc606_5 gpc9082 (
      {stage2_56[114], stage2_56[115], stage2_56[116], stage2_56[117], stage2_56[118], stage2_56[119]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[5],stage3_58[24],stage3_57[36],stage3_56[36]}
   );
   gpc606_5 gpc9083 (
      {stage2_56[120], stage2_56[121], stage2_56[122], stage2_56[123], stage2_56[124], stage2_56[125]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[6],stage3_58[25],stage3_57[37],stage3_56[37]}
   );
   gpc606_5 gpc9084 (
      {stage2_56[126], stage2_56[127], stage2_56[128], stage2_56[129], stage2_56[130], stage2_56[131]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[7],stage3_58[26],stage3_57[38],stage3_56[38]}
   );
   gpc606_5 gpc9085 (
      {stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33], stage2_57[34], stage2_57[35]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[3],stage3_59[8],stage3_58[27],stage3_57[39]}
   );
   gpc606_5 gpc9086 (
      {stage2_57[36], stage2_57[37], stage2_57[38], stage2_57[39], stage2_57[40], stage2_57[41]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[4],stage3_59[9],stage3_58[28],stage3_57[40]}
   );
   gpc606_5 gpc9087 (
      {stage2_57[42], stage2_57[43], stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[5],stage3_59[10],stage3_58[29],stage3_57[41]}
   );
   gpc606_5 gpc9088 (
      {stage2_57[48], stage2_57[49], stage2_57[50], stage2_57[51], stage2_57[52], stage2_57[53]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[6],stage3_59[11],stage3_58[30],stage3_57[42]}
   );
   gpc606_5 gpc9089 (
      {stage2_57[54], stage2_57[55], stage2_57[56], stage2_57[57], stage2_57[58], stage2_57[59]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[7],stage3_59[12],stage3_58[31],stage3_57[43]}
   );
   gpc606_5 gpc9090 (
      {stage2_57[60], stage2_57[61], stage2_57[62], stage2_57[63], stage2_57[64], stage2_57[65]},
      {stage2_59[30], stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35]},
      {stage3_61[5],stage3_60[8],stage3_59[13],stage3_58[32],stage3_57[44]}
   );
   gpc606_5 gpc9091 (
      {stage2_57[66], stage2_57[67], stage2_57[68], stage2_57[69], stage2_57[70], stage2_57[71]},
      {stage2_59[36], stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41]},
      {stage3_61[6],stage3_60[9],stage3_59[14],stage3_58[33],stage3_57[45]}
   );
   gpc207_4 gpc9092 (
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23], stage2_58[24]},
      {stage2_60[0], stage2_60[1]},
      {stage3_61[7],stage3_60[10],stage3_59[15],stage3_58[34]}
   );
   gpc207_4 gpc9093 (
      {stage2_58[25], stage2_58[26], stage2_58[27], stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31]},
      {stage2_60[2], stage2_60[3]},
      {stage3_61[8],stage3_60[11],stage3_59[16],stage3_58[35]}
   );
   gpc207_4 gpc9094 (
      {stage2_58[32], stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37], stage2_58[38]},
      {stage2_60[4], stage2_60[5]},
      {stage3_61[9],stage3_60[12],stage3_59[17],stage3_58[36]}
   );
   gpc207_4 gpc9095 (
      {stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42], stage2_58[43], stage2_58[44], stage2_58[45]},
      {stage2_60[6], stage2_60[7]},
      {stage3_61[10],stage3_60[13],stage3_59[18],stage3_58[37]}
   );
   gpc207_4 gpc9096 (
      {stage2_58[46], stage2_58[47], stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_60[8], stage2_60[9]},
      {stage3_61[11],stage3_60[14],stage3_59[19],stage3_58[38]}
   );
   gpc207_4 gpc9097 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57], stage2_58[58], stage2_58[59]},
      {stage2_60[10], stage2_60[11]},
      {stage3_61[12],stage3_60[15],stage3_59[20],stage3_58[39]}
   );
   gpc207_4 gpc9098 (
      {stage2_58[60], stage2_58[61], stage2_58[62], stage2_58[63], stage2_58[64], stage2_58[65], stage2_58[66]},
      {stage2_60[12], stage2_60[13]},
      {stage3_61[13],stage3_60[16],stage3_59[21],stage3_58[40]}
   );
   gpc207_4 gpc9099 (
      {stage2_58[67], stage2_58[68], stage2_58[69], stage2_58[70], stage2_58[71], stage2_58[72], stage2_58[73]},
      {stage2_60[14], stage2_60[15]},
      {stage3_61[14],stage3_60[17],stage3_59[22],stage3_58[41]}
   );
   gpc615_5 gpc9100 (
      {stage2_58[74], stage2_58[75], stage2_58[76], stage2_58[77], stage2_58[78]},
      {stage2_59[42]},
      {stage2_60[16], stage2_60[17], stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21]},
      {stage3_62[0],stage3_61[15],stage3_60[18],stage3_59[23],stage3_58[42]}
   );
   gpc606_5 gpc9101 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[1],stage3_61[16],stage3_60[19],stage3_59[24]}
   );
   gpc606_5 gpc9102 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[2],stage3_61[17],stage3_60[20],stage3_59[25]}
   );
   gpc606_5 gpc9103 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59], stage2_59[60]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[3],stage3_61[18],stage3_60[21],stage3_59[26]}
   );
   gpc606_5 gpc9104 (
      {stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64], stage2_59[65], stage2_59[66]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[4],stage3_61[19],stage3_60[22],stage3_59[27]}
   );
   gpc606_5 gpc9105 (
      {stage2_59[67], stage2_59[68], stage2_59[69], stage2_59[70], stage2_59[71], stage2_59[72]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[5],stage3_61[20],stage3_60[23],stage3_59[28]}
   );
   gpc606_5 gpc9106 (
      {stage2_59[73], stage2_59[74], stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[6],stage3_61[21],stage3_60[24],stage3_59[29]}
   );
   gpc606_5 gpc9107 (
      {stage2_59[79], stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[7],stage3_61[22],stage3_60[25],stage3_59[30]}
   );
   gpc606_5 gpc9108 (
      {stage2_59[85], stage2_59[86], stage2_59[87], stage2_59[88], stage2_59[89], stage2_59[90]},
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage3_63[7],stage3_62[8],stage3_61[23],stage3_60[26],stage3_59[31]}
   );
   gpc606_5 gpc9109 (
      {stage2_59[91], stage2_59[92], stage2_59[93], stage2_59[94], stage2_59[95], stage2_59[96]},
      {stage2_61[48], stage2_61[49], stage2_61[50], stage2_61[51], stage2_61[52], stage2_61[53]},
      {stage3_63[8],stage3_62[9],stage3_61[24],stage3_60[27],stage3_59[32]}
   );
   gpc606_5 gpc9110 (
      {stage2_59[97], stage2_59[98], stage2_59[99], stage2_59[100], stage2_59[101], stage2_59[102]},
      {stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58], stage2_61[59]},
      {stage3_63[9],stage3_62[10],stage3_61[25],stage3_60[28],stage3_59[33]}
   );
   gpc606_5 gpc9111 (
      {stage2_59[103], stage2_59[104], stage2_59[105], stage2_59[106], stage2_59[107], stage2_59[108]},
      {stage2_61[60], stage2_61[61], stage2_61[62], stage2_61[63], stage2_61[64], stage2_61[65]},
      {stage3_63[10],stage3_62[11],stage3_61[26],stage3_60[29],stage3_59[34]}
   );
   gpc606_5 gpc9112 (
      {stage2_59[109], stage2_59[110], stage2_59[111], stage2_59[112], stage2_59[113], stage2_59[114]},
      {stage2_61[66], stage2_61[67], stage2_61[68], stage2_61[69], stage2_61[70], stage2_61[71]},
      {stage3_63[11],stage3_62[12],stage3_61[27],stage3_60[30],stage3_59[35]}
   );
   gpc606_5 gpc9113 (
      {stage2_59[115], stage2_59[116], stage2_59[117], stage2_59[118], stage2_59[119], stage2_59[120]},
      {stage2_61[72], stage2_61[73], stage2_61[74], stage2_61[75], stage2_61[76], stage2_61[77]},
      {stage3_63[12],stage3_62[13],stage3_61[28],stage3_60[31],stage3_59[36]}
   );
   gpc606_5 gpc9114 (
      {stage2_59[121], stage2_59[122], stage2_59[123], stage2_59[124], stage2_59[125], stage2_59[126]},
      {stage2_61[78], stage2_61[79], stage2_61[80], stage2_61[81], stage2_61[82], stage2_61[83]},
      {stage3_63[13],stage3_62[14],stage3_61[29],stage3_60[32],stage3_59[37]}
   );
   gpc606_5 gpc9115 (
      {stage2_59[127], stage2_59[128], stage2_59[129], stage2_59[130], stage2_59[131], stage2_59[132]},
      {stage2_61[84], stage2_61[85], stage2_61[86], stage2_61[87], stage2_61[88], stage2_61[89]},
      {stage3_63[14],stage3_62[15],stage3_61[30],stage3_60[33],stage3_59[38]}
   );
   gpc606_5 gpc9116 (
      {stage2_60[22], stage2_60[23], stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[15],stage3_62[16],stage3_61[31],stage3_60[34]}
   );
   gpc606_5 gpc9117 (
      {stage2_60[28], stage2_60[29], stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[16],stage3_62[17],stage3_61[32],stage3_60[35]}
   );
   gpc606_5 gpc9118 (
      {stage2_60[34], stage2_60[35], stage2_60[36], stage2_60[37], stage2_60[38], stage2_60[39]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[17],stage3_62[18],stage3_61[33],stage3_60[36]}
   );
   gpc606_5 gpc9119 (
      {stage2_60[40], stage2_60[41], stage2_60[42], stage2_60[43], stage2_60[44], stage2_60[45]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[18],stage3_62[19],stage3_61[34],stage3_60[37]}
   );
   gpc606_5 gpc9120 (
      {stage2_60[46], stage2_60[47], stage2_60[48], stage2_60[49], stage2_60[50], stage2_60[51]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[19],stage3_62[20],stage3_61[35],stage3_60[38]}
   );
   gpc606_5 gpc9121 (
      {stage2_60[52], stage2_60[53], stage2_60[54], stage2_60[55], stage2_60[56], stage2_60[57]},
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34], stage2_62[35]},
      {stage3_64[5],stage3_63[20],stage3_62[21],stage3_61[36],stage3_60[39]}
   );
   gpc606_5 gpc9122 (
      {stage2_60[58], stage2_60[59], stage2_60[60], stage2_60[61], stage2_60[62], stage2_60[63]},
      {stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39], stage2_62[40], stage2_62[41]},
      {stage3_64[6],stage3_63[21],stage3_62[22],stage3_61[37],stage3_60[40]}
   );
   gpc606_5 gpc9123 (
      {stage2_60[64], stage2_60[65], stage2_60[66], stage2_60[67], stage2_60[68], stage2_60[69]},
      {stage2_62[42], stage2_62[43], stage2_62[44], stage2_62[45], stage2_62[46], stage2_62[47]},
      {stage3_64[7],stage3_63[22],stage3_62[23],stage3_61[38],stage3_60[41]}
   );
   gpc606_5 gpc9124 (
      {stage2_60[70], stage2_60[71], stage2_60[72], stage2_60[73], stage2_60[74], stage2_60[75]},
      {stage2_62[48], stage2_62[49], stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53]},
      {stage3_64[8],stage3_63[23],stage3_62[24],stage3_61[39],stage3_60[42]}
   );
   gpc606_5 gpc9125 (
      {stage2_60[76], stage2_60[77], stage2_60[78], stage2_60[79], stage2_60[80], stage2_60[81]},
      {stage2_62[54], stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage3_64[9],stage3_63[24],stage3_62[25],stage3_61[40],stage3_60[43]}
   );
   gpc606_5 gpc9126 (
      {stage2_60[82], stage2_60[83], stage2_60[84], stage2_60[85], stage2_60[86], stage2_60[87]},
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64], stage2_62[65]},
      {stage3_64[10],stage3_63[25],stage3_62[26],stage3_61[41],stage3_60[44]}
   );
   gpc606_5 gpc9127 (
      {stage2_60[88], stage2_60[89], stage2_60[90], stage2_60[91], stage2_60[92], stage2_60[93]},
      {stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69], stage2_62[70], stage2_62[71]},
      {stage3_64[11],stage3_63[26],stage3_62[27],stage3_61[42],stage3_60[45]}
   );
   gpc606_5 gpc9128 (
      {stage2_60[94], stage2_60[95], stage2_60[96], stage2_60[97], stage2_60[98], stage2_60[99]},
      {stage2_62[72], stage2_62[73], stage2_62[74], stage2_62[75], stage2_62[76], stage2_62[77]},
      {stage3_64[12],stage3_63[27],stage3_62[28],stage3_61[43],stage3_60[46]}
   );
   gpc606_5 gpc9129 (
      {stage2_60[100], stage2_60[101], stage2_60[102], stage2_60[103], stage2_60[104], stage2_60[105]},
      {stage2_62[78], stage2_62[79], stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83]},
      {stage3_64[13],stage3_63[28],stage3_62[29],stage3_61[44],stage3_60[47]}
   );
   gpc606_5 gpc9130 (
      {stage2_62[84], stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[0],stage3_64[14],stage3_63[29],stage3_62[30]}
   );
   gpc606_5 gpc9131 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94], stage2_62[95]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[1],stage3_64[15],stage3_63[30],stage3_62[31]}
   );
   gpc606_5 gpc9132 (
      {stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99], stage2_62[100], stage2_62[101]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[2],stage3_64[16],stage3_63[31],stage3_62[32]}
   );
   gpc606_5 gpc9133 (
      {stage2_62[102], stage2_62[103], stage2_62[104], stage2_62[105], stage2_62[106], stage2_62[107]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[3],stage3_64[17],stage3_63[32],stage3_62[33]}
   );
   gpc606_5 gpc9134 (
      {stage2_62[108], stage2_62[109], stage2_62[110], stage2_62[111], stage2_62[112], stage2_62[113]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[4],stage3_64[18],stage3_63[33],stage3_62[34]}
   );
   gpc606_5 gpc9135 (
      {stage2_62[114], stage2_62[115], stage2_62[116], stage2_62[117], stage2_62[118], stage2_62[119]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[5],stage3_64[19],stage3_63[34],stage3_62[35]}
   );
   gpc606_5 gpc9136 (
      {stage2_62[120], stage2_62[121], stage2_62[122], stage2_62[123], stage2_62[124], stage2_62[125]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[6],stage3_64[20],stage3_63[35],stage3_62[36]}
   );
   gpc606_5 gpc9137 (
      {stage2_62[126], stage2_62[127], stage2_62[128], stage2_62[129], stage2_62[130], stage2_62[131]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[7],stage3_64[21],stage3_63[36],stage3_62[37]}
   );
   gpc606_5 gpc9138 (
      {stage2_62[132], stage2_62[133], stage2_62[134], stage2_62[135], stage2_62[136], stage2_62[137]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[8],stage3_64[22],stage3_63[37],stage3_62[38]}
   );
   gpc606_5 gpc9139 (
      {stage2_62[138], stage2_62[139], stage2_62[140], stage2_62[141], stage2_62[142], stage2_62[143]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[9],stage3_64[23],stage3_63[38],stage3_62[39]}
   );
   gpc117_4 gpc9140 (
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage2_64[60]},
      {stage2_65[0]},
      {stage3_66[10],stage3_65[10],stage3_64[24],stage3_63[39]}
   );
   gpc117_4 gpc9141 (
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12], stage2_63[13]},
      {stage2_64[61]},
      {stage2_65[1]},
      {stage3_66[11],stage3_65[11],stage3_64[25],stage3_63[40]}
   );
   gpc117_4 gpc9142 (
      {stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18], stage2_63[19], stage2_63[20]},
      {stage2_64[62]},
      {stage2_65[2]},
      {stage3_66[12],stage3_65[12],stage3_64[26],stage3_63[41]}
   );
   gpc117_4 gpc9143 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[63]},
      {stage2_65[3]},
      {stage3_66[13],stage3_65[13],stage3_64[27],stage3_63[42]}
   );
   gpc117_4 gpc9144 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[64]},
      {stage2_65[4]},
      {stage3_66[14],stage3_65[14],stage3_64[28],stage3_63[43]}
   );
   gpc606_5 gpc9145 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40]},
      {stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9], stage2_65[10]},
      {stage3_67[0],stage3_66[15],stage3_65[15],stage3_64[29],stage3_63[44]}
   );
   gpc606_5 gpc9146 (
      {stage2_63[41], stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46]},
      {stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14], stage2_65[15], stage2_65[16]},
      {stage3_67[1],stage3_66[16],stage3_65[16],stage3_64[30],stage3_63[45]}
   );
   gpc606_5 gpc9147 (
      {stage2_63[47], stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52]},
      {stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20], stage2_65[21], stage2_65[22]},
      {stage3_67[2],stage3_66[17],stage3_65[17],stage3_64[31],stage3_63[46]}
   );
   gpc606_5 gpc9148 (
      {stage2_63[53], stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58]},
      {stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26], stage2_65[27], stage2_65[28]},
      {stage3_67[3],stage3_66[18],stage3_65[18],stage3_64[32],stage3_63[47]}
   );
   gpc606_5 gpc9149 (
      {stage2_63[59], stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64]},
      {stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32], stage2_65[33], stage2_65[34]},
      {stage3_67[4],stage3_66[19],stage3_65[19],stage3_64[33],stage3_63[48]}
   );
   gpc606_5 gpc9150 (
      {stage2_63[65], stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70]},
      {stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38], stage2_65[39], stage2_65[40]},
      {stage3_67[5],stage3_66[20],stage3_65[20],stage3_64[34],stage3_63[49]}
   );
   gpc606_5 gpc9151 (
      {stage2_63[71], stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76]},
      {stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44], stage2_65[45], stage2_65[46]},
      {stage3_67[6],stage3_66[21],stage3_65[21],stage3_64[35],stage3_63[50]}
   );
   gpc606_5 gpc9152 (
      {stage2_63[77], stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82]},
      {stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50], stage2_65[51], stage2_65[52]},
      {stage3_67[7],stage3_66[22],stage3_65[22],stage3_64[36],stage3_63[51]}
   );
   gpc606_5 gpc9153 (
      {stage2_63[83], stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88]},
      {stage2_65[53], stage2_65[54], stage2_65[55], stage2_65[56], stage2_65[57], stage2_65[58]},
      {stage3_67[8],stage3_66[23],stage3_65[23],stage3_64[37],stage3_63[52]}
   );
   gpc606_5 gpc9154 (
      {stage2_63[89], stage2_63[90], stage2_63[91], stage2_63[92], stage2_63[93], stage2_63[94]},
      {stage2_65[59], stage2_65[60], stage2_65[61], stage2_65[62], stage2_65[63], stage2_65[64]},
      {stage3_67[9],stage3_66[24],stage3_65[24],stage3_64[38],stage3_63[53]}
   );
   gpc606_5 gpc9155 (
      {stage2_64[65], stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[10],stage3_66[25],stage3_65[25],stage3_64[39]}
   );
   gpc606_5 gpc9156 (
      {stage2_64[71], stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[11],stage3_66[26],stage3_65[26],stage3_64[40]}
   );
   gpc606_5 gpc9157 (
      {stage2_64[77], stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[12],stage3_66[27],stage3_65[27],stage3_64[41]}
   );
   gpc606_5 gpc9158 (
      {stage2_64[83], stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[13],stage3_66[28],stage3_65[28],stage3_64[42]}
   );
   gpc606_5 gpc9159 (
      {stage2_64[89], stage2_64[90], stage2_64[91], stage2_64[92], stage2_64[93], stage2_64[94]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[14],stage3_66[29],stage3_65[29],stage3_64[43]}
   );
   gpc1_1 gpc9160 (
      {stage2_0[29]},
      {stage3_0[6]}
   );
   gpc1_1 gpc9161 (
      {stage2_0[30]},
      {stage3_0[7]}
   );
   gpc1_1 gpc9162 (
      {stage2_0[31]},
      {stage3_0[8]}
   );
   gpc1_1 gpc9163 (
      {stage2_0[32]},
      {stage3_0[9]}
   );
   gpc1_1 gpc9164 (
      {stage2_0[33]},
      {stage3_0[10]}
   );
   gpc1_1 gpc9165 (
      {stage2_1[22]},
      {stage3_1[9]}
   );
   gpc1_1 gpc9166 (
      {stage2_1[23]},
      {stage3_1[10]}
   );
   gpc1_1 gpc9167 (
      {stage2_1[24]},
      {stage3_1[11]}
   );
   gpc1_1 gpc9168 (
      {stage2_1[25]},
      {stage3_1[12]}
   );
   gpc1_1 gpc9169 (
      {stage2_1[26]},
      {stage3_1[13]}
   );
   gpc1_1 gpc9170 (
      {stage2_1[27]},
      {stage3_1[14]}
   );
   gpc1_1 gpc9171 (
      {stage2_1[28]},
      {stage3_1[15]}
   );
   gpc1_1 gpc9172 (
      {stage2_1[29]},
      {stage3_1[16]}
   );
   gpc1_1 gpc9173 (
      {stage2_1[30]},
      {stage3_1[17]}
   );
   gpc1_1 gpc9174 (
      {stage2_1[31]},
      {stage3_1[18]}
   );
   gpc1_1 gpc9175 (
      {stage2_1[32]},
      {stage3_1[19]}
   );
   gpc1_1 gpc9176 (
      {stage2_1[33]},
      {stage3_1[20]}
   );
   gpc1_1 gpc9177 (
      {stage2_1[34]},
      {stage3_1[21]}
   );
   gpc1_1 gpc9178 (
      {stage2_1[35]},
      {stage3_1[22]}
   );
   gpc1_1 gpc9179 (
      {stage2_1[36]},
      {stage3_1[23]}
   );
   gpc1_1 gpc9180 (
      {stage2_1[37]},
      {stage3_1[24]}
   );
   gpc1_1 gpc9181 (
      {stage2_1[38]},
      {stage3_1[25]}
   );
   gpc1_1 gpc9182 (
      {stage2_7[85]},
      {stage3_7[43]}
   );
   gpc1_1 gpc9183 (
      {stage2_7[86]},
      {stage3_7[44]}
   );
   gpc1_1 gpc9184 (
      {stage2_7[87]},
      {stage3_7[45]}
   );
   gpc1_1 gpc9185 (
      {stage2_7[88]},
      {stage3_7[46]}
   );
   gpc1_1 gpc9186 (
      {stage2_7[89]},
      {stage3_7[47]}
   );
   gpc1_1 gpc9187 (
      {stage2_7[90]},
      {stage3_7[48]}
   );
   gpc1_1 gpc9188 (
      {stage2_7[91]},
      {stage3_7[49]}
   );
   gpc1_1 gpc9189 (
      {stage2_7[92]},
      {stage3_7[50]}
   );
   gpc1_1 gpc9190 (
      {stage2_7[93]},
      {stage3_7[51]}
   );
   gpc1_1 gpc9191 (
      {stage2_7[94]},
      {stage3_7[52]}
   );
   gpc1_1 gpc9192 (
      {stage2_7[95]},
      {stage3_7[53]}
   );
   gpc1_1 gpc9193 (
      {stage2_7[96]},
      {stage3_7[54]}
   );
   gpc1_1 gpc9194 (
      {stage2_10[125]},
      {stage3_10[59]}
   );
   gpc1_1 gpc9195 (
      {stage2_10[126]},
      {stage3_10[60]}
   );
   gpc1_1 gpc9196 (
      {stage2_10[127]},
      {stage3_10[61]}
   );
   gpc1_1 gpc9197 (
      {stage2_10[128]},
      {stage3_10[62]}
   );
   gpc1_1 gpc9198 (
      {stage2_10[129]},
      {stage3_10[63]}
   );
   gpc1_1 gpc9199 (
      {stage2_10[130]},
      {stage3_10[64]}
   );
   gpc1_1 gpc9200 (
      {stage2_10[131]},
      {stage3_10[65]}
   );
   gpc1_1 gpc9201 (
      {stage2_10[132]},
      {stage3_10[66]}
   );
   gpc1_1 gpc9202 (
      {stage2_10[133]},
      {stage3_10[67]}
   );
   gpc1_1 gpc9203 (
      {stage2_11[125]},
      {stage3_11[50]}
   );
   gpc1_1 gpc9204 (
      {stage2_11[126]},
      {stage3_11[51]}
   );
   gpc1_1 gpc9205 (
      {stage2_11[127]},
      {stage3_11[52]}
   );
   gpc1_1 gpc9206 (
      {stage2_11[128]},
      {stage3_11[53]}
   );
   gpc1_1 gpc9207 (
      {stage2_11[129]},
      {stage3_11[54]}
   );
   gpc1_1 gpc9208 (
      {stage2_11[130]},
      {stage3_11[55]}
   );
   gpc1_1 gpc9209 (
      {stage2_11[131]},
      {stage3_11[56]}
   );
   gpc1_1 gpc9210 (
      {stage2_11[132]},
      {stage3_11[57]}
   );
   gpc1_1 gpc9211 (
      {stage2_11[133]},
      {stage3_11[58]}
   );
   gpc1_1 gpc9212 (
      {stage2_11[134]},
      {stage3_11[59]}
   );
   gpc1_1 gpc9213 (
      {stage2_11[135]},
      {stage3_11[60]}
   );
   gpc1_1 gpc9214 (
      {stage2_12[98]},
      {stage3_12[51]}
   );
   gpc1_1 gpc9215 (
      {stage2_12[99]},
      {stage3_12[52]}
   );
   gpc1_1 gpc9216 (
      {stage2_12[100]},
      {stage3_12[53]}
   );
   gpc1_1 gpc9217 (
      {stage2_12[101]},
      {stage3_12[54]}
   );
   gpc1_1 gpc9218 (
      {stage2_12[102]},
      {stage3_12[55]}
   );
   gpc1_1 gpc9219 (
      {stage2_12[103]},
      {stage3_12[56]}
   );
   gpc1_1 gpc9220 (
      {stage2_12[104]},
      {stage3_12[57]}
   );
   gpc1_1 gpc9221 (
      {stage2_12[105]},
      {stage3_12[58]}
   );
   gpc1_1 gpc9222 (
      {stage2_12[106]},
      {stage3_12[59]}
   );
   gpc1_1 gpc9223 (
      {stage2_12[107]},
      {stage3_12[60]}
   );
   gpc1_1 gpc9224 (
      {stage2_12[108]},
      {stage3_12[61]}
   );
   gpc1_1 gpc9225 (
      {stage2_12[109]},
      {stage3_12[62]}
   );
   gpc1_1 gpc9226 (
      {stage2_12[110]},
      {stage3_12[63]}
   );
   gpc1_1 gpc9227 (
      {stage2_12[111]},
      {stage3_12[64]}
   );
   gpc1_1 gpc9228 (
      {stage2_12[112]},
      {stage3_12[65]}
   );
   gpc1_1 gpc9229 (
      {stage2_12[113]},
      {stage3_12[66]}
   );
   gpc1_1 gpc9230 (
      {stage2_12[114]},
      {stage3_12[67]}
   );
   gpc1_1 gpc9231 (
      {stage2_12[115]},
      {stage3_12[68]}
   );
   gpc1_1 gpc9232 (
      {stage2_12[116]},
      {stage3_12[69]}
   );
   gpc1_1 gpc9233 (
      {stage2_12[117]},
      {stage3_12[70]}
   );
   gpc1_1 gpc9234 (
      {stage2_12[118]},
      {stage3_12[71]}
   );
   gpc1_1 gpc9235 (
      {stage2_12[119]},
      {stage3_12[72]}
   );
   gpc1_1 gpc9236 (
      {stage2_12[120]},
      {stage3_12[73]}
   );
   gpc1_1 gpc9237 (
      {stage2_12[121]},
      {stage3_12[74]}
   );
   gpc1_1 gpc9238 (
      {stage2_12[122]},
      {stage3_12[75]}
   );
   gpc1_1 gpc9239 (
      {stage2_12[123]},
      {stage3_12[76]}
   );
   gpc1_1 gpc9240 (
      {stage2_12[124]},
      {stage3_12[77]}
   );
   gpc1_1 gpc9241 (
      {stage2_12[125]},
      {stage3_12[78]}
   );
   gpc1_1 gpc9242 (
      {stage2_12[126]},
      {stage3_12[79]}
   );
   gpc1_1 gpc9243 (
      {stage2_12[127]},
      {stage3_12[80]}
   );
   gpc1_1 gpc9244 (
      {stage2_13[70]},
      {stage3_13[45]}
   );
   gpc1_1 gpc9245 (
      {stage2_13[71]},
      {stage3_13[46]}
   );
   gpc1_1 gpc9246 (
      {stage2_15[108]},
      {stage3_15[44]}
   );
   gpc1_1 gpc9247 (
      {stage2_15[109]},
      {stage3_15[45]}
   );
   gpc1_1 gpc9248 (
      {stage2_15[110]},
      {stage3_15[46]}
   );
   gpc1_1 gpc9249 (
      {stage2_15[111]},
      {stage3_15[47]}
   );
   gpc1_1 gpc9250 (
      {stage2_15[112]},
      {stage3_15[48]}
   );
   gpc1_1 gpc9251 (
      {stage2_15[113]},
      {stage3_15[49]}
   );
   gpc1_1 gpc9252 (
      {stage2_15[114]},
      {stage3_15[50]}
   );
   gpc1_1 gpc9253 (
      {stage2_16[96]},
      {stage3_16[45]}
   );
   gpc1_1 gpc9254 (
      {stage2_16[97]},
      {stage3_16[46]}
   );
   gpc1_1 gpc9255 (
      {stage2_16[98]},
      {stage3_16[47]}
   );
   gpc1_1 gpc9256 (
      {stage2_16[99]},
      {stage3_16[48]}
   );
   gpc1_1 gpc9257 (
      {stage2_16[100]},
      {stage3_16[49]}
   );
   gpc1_1 gpc9258 (
      {stage2_16[101]},
      {stage3_16[50]}
   );
   gpc1_1 gpc9259 (
      {stage2_16[102]},
      {stage3_16[51]}
   );
   gpc1_1 gpc9260 (
      {stage2_16[103]},
      {stage3_16[52]}
   );
   gpc1_1 gpc9261 (
      {stage2_16[104]},
      {stage3_16[53]}
   );
   gpc1_1 gpc9262 (
      {stage2_16[105]},
      {stage3_16[54]}
   );
   gpc1_1 gpc9263 (
      {stage2_16[106]},
      {stage3_16[55]}
   );
   gpc1_1 gpc9264 (
      {stage2_16[107]},
      {stage3_16[56]}
   );
   gpc1_1 gpc9265 (
      {stage2_16[108]},
      {stage3_16[57]}
   );
   gpc1_1 gpc9266 (
      {stage2_16[109]},
      {stage3_16[58]}
   );
   gpc1_1 gpc9267 (
      {stage2_17[80]},
      {stage3_17[34]}
   );
   gpc1_1 gpc9268 (
      {stage2_17[81]},
      {stage3_17[35]}
   );
   gpc1_1 gpc9269 (
      {stage2_17[82]},
      {stage3_17[36]}
   );
   gpc1_1 gpc9270 (
      {stage2_17[83]},
      {stage3_17[37]}
   );
   gpc1_1 gpc9271 (
      {stage2_17[84]},
      {stage3_17[38]}
   );
   gpc1_1 gpc9272 (
      {stage2_17[85]},
      {stage3_17[39]}
   );
   gpc1_1 gpc9273 (
      {stage2_17[86]},
      {stage3_17[40]}
   );
   gpc1_1 gpc9274 (
      {stage2_17[87]},
      {stage3_17[41]}
   );
   gpc1_1 gpc9275 (
      {stage2_17[88]},
      {stage3_17[42]}
   );
   gpc1_1 gpc9276 (
      {stage2_17[89]},
      {stage3_17[43]}
   );
   gpc1_1 gpc9277 (
      {stage2_18[147]},
      {stage3_18[49]}
   );
   gpc1_1 gpc9278 (
      {stage2_18[148]},
      {stage3_18[50]}
   );
   gpc1_1 gpc9279 (
      {stage2_18[149]},
      {stage3_18[51]}
   );
   gpc1_1 gpc9280 (
      {stage2_18[150]},
      {stage3_18[52]}
   );
   gpc1_1 gpc9281 (
      {stage2_18[151]},
      {stage3_18[53]}
   );
   gpc1_1 gpc9282 (
      {stage2_18[152]},
      {stage3_18[54]}
   );
   gpc1_1 gpc9283 (
      {stage2_18[153]},
      {stage3_18[55]}
   );
   gpc1_1 gpc9284 (
      {stage2_18[154]},
      {stage3_18[56]}
   );
   gpc1_1 gpc9285 (
      {stage2_18[155]},
      {stage3_18[57]}
   );
   gpc1_1 gpc9286 (
      {stage2_18[156]},
      {stage3_18[58]}
   );
   gpc1_1 gpc9287 (
      {stage2_18[157]},
      {stage3_18[59]}
   );
   gpc1_1 gpc9288 (
      {stage2_18[158]},
      {stage3_18[60]}
   );
   gpc1_1 gpc9289 (
      {stage2_18[159]},
      {stage3_18[61]}
   );
   gpc1_1 gpc9290 (
      {stage2_18[160]},
      {stage3_18[62]}
   );
   gpc1_1 gpc9291 (
      {stage2_18[161]},
      {stage3_18[63]}
   );
   gpc1_1 gpc9292 (
      {stage2_20[72]},
      {stage3_20[42]}
   );
   gpc1_1 gpc9293 (
      {stage2_20[73]},
      {stage3_20[43]}
   );
   gpc1_1 gpc9294 (
      {stage2_20[74]},
      {stage3_20[44]}
   );
   gpc1_1 gpc9295 (
      {stage2_20[75]},
      {stage3_20[45]}
   );
   gpc1_1 gpc9296 (
      {stage2_20[76]},
      {stage3_20[46]}
   );
   gpc1_1 gpc9297 (
      {stage2_20[77]},
      {stage3_20[47]}
   );
   gpc1_1 gpc9298 (
      {stage2_20[78]},
      {stage3_20[48]}
   );
   gpc1_1 gpc9299 (
      {stage2_20[79]},
      {stage3_20[49]}
   );
   gpc1_1 gpc9300 (
      {stage2_20[80]},
      {stage3_20[50]}
   );
   gpc1_1 gpc9301 (
      {stage2_20[81]},
      {stage3_20[51]}
   );
   gpc1_1 gpc9302 (
      {stage2_20[82]},
      {stage3_20[52]}
   );
   gpc1_1 gpc9303 (
      {stage2_20[83]},
      {stage3_20[53]}
   );
   gpc1_1 gpc9304 (
      {stage2_20[84]},
      {stage3_20[54]}
   );
   gpc1_1 gpc9305 (
      {stage2_20[85]},
      {stage3_20[55]}
   );
   gpc1_1 gpc9306 (
      {stage2_20[86]},
      {stage3_20[56]}
   );
   gpc1_1 gpc9307 (
      {stage2_20[87]},
      {stage3_20[57]}
   );
   gpc1_1 gpc9308 (
      {stage2_21[86]},
      {stage3_21[37]}
   );
   gpc1_1 gpc9309 (
      {stage2_21[87]},
      {stage3_21[38]}
   );
   gpc1_1 gpc9310 (
      {stage2_21[88]},
      {stage3_21[39]}
   );
   gpc1_1 gpc9311 (
      {stage2_21[89]},
      {stage3_21[40]}
   );
   gpc1_1 gpc9312 (
      {stage2_21[90]},
      {stage3_21[41]}
   );
   gpc1_1 gpc9313 (
      {stage2_21[91]},
      {stage3_21[42]}
   );
   gpc1_1 gpc9314 (
      {stage2_21[92]},
      {stage3_21[43]}
   );
   gpc1_1 gpc9315 (
      {stage2_21[93]},
      {stage3_21[44]}
   );
   gpc1_1 gpc9316 (
      {stage2_21[94]},
      {stage3_21[45]}
   );
   gpc1_1 gpc9317 (
      {stage2_21[95]},
      {stage3_21[46]}
   );
   gpc1_1 gpc9318 (
      {stage2_21[96]},
      {stage3_21[47]}
   );
   gpc1_1 gpc9319 (
      {stage2_21[97]},
      {stage3_21[48]}
   );
   gpc1_1 gpc9320 (
      {stage2_21[98]},
      {stage3_21[49]}
   );
   gpc1_1 gpc9321 (
      {stage2_21[99]},
      {stage3_21[50]}
   );
   gpc1_1 gpc9322 (
      {stage2_21[100]},
      {stage3_21[51]}
   );
   gpc1_1 gpc9323 (
      {stage2_21[101]},
      {stage3_21[52]}
   );
   gpc1_1 gpc9324 (
      {stage2_21[102]},
      {stage3_21[53]}
   );
   gpc1_1 gpc9325 (
      {stage2_21[103]},
      {stage3_21[54]}
   );
   gpc1_1 gpc9326 (
      {stage2_21[104]},
      {stage3_21[55]}
   );
   gpc1_1 gpc9327 (
      {stage2_21[105]},
      {stage3_21[56]}
   );
   gpc1_1 gpc9328 (
      {stage2_21[106]},
      {stage3_21[57]}
   );
   gpc1_1 gpc9329 (
      {stage2_21[107]},
      {stage3_21[58]}
   );
   gpc1_1 gpc9330 (
      {stage2_21[108]},
      {stage3_21[59]}
   );
   gpc1_1 gpc9331 (
      {stage2_21[109]},
      {stage3_21[60]}
   );
   gpc1_1 gpc9332 (
      {stage2_21[110]},
      {stage3_21[61]}
   );
   gpc1_1 gpc9333 (
      {stage2_21[111]},
      {stage3_21[62]}
   );
   gpc1_1 gpc9334 (
      {stage2_22[108]},
      {stage3_22[48]}
   );
   gpc1_1 gpc9335 (
      {stage2_22[109]},
      {stage3_22[49]}
   );
   gpc1_1 gpc9336 (
      {stage2_23[89]},
      {stage3_23[40]}
   );
   gpc1_1 gpc9337 (
      {stage2_23[90]},
      {stage3_23[41]}
   );
   gpc1_1 gpc9338 (
      {stage2_23[91]},
      {stage3_23[42]}
   );
   gpc1_1 gpc9339 (
      {stage2_23[92]},
      {stage3_23[43]}
   );
   gpc1_1 gpc9340 (
      {stage2_23[93]},
      {stage3_23[44]}
   );
   gpc1_1 gpc9341 (
      {stage2_23[94]},
      {stage3_23[45]}
   );
   gpc1_1 gpc9342 (
      {stage2_23[95]},
      {stage3_23[46]}
   );
   gpc1_1 gpc9343 (
      {stage2_23[96]},
      {stage3_23[47]}
   );
   gpc1_1 gpc9344 (
      {stage2_23[97]},
      {stage3_23[48]}
   );
   gpc1_1 gpc9345 (
      {stage2_25[102]},
      {stage3_25[31]}
   );
   gpc1_1 gpc9346 (
      {stage2_25[103]},
      {stage3_25[32]}
   );
   gpc1_1 gpc9347 (
      {stage2_25[104]},
      {stage3_25[33]}
   );
   gpc1_1 gpc9348 (
      {stage2_25[105]},
      {stage3_25[34]}
   );
   gpc1_1 gpc9349 (
      {stage2_25[106]},
      {stage3_25[35]}
   );
   gpc1_1 gpc9350 (
      {stage2_25[107]},
      {stage3_25[36]}
   );
   gpc1_1 gpc9351 (
      {stage2_25[108]},
      {stage3_25[37]}
   );
   gpc1_1 gpc9352 (
      {stage2_25[109]},
      {stage3_25[38]}
   );
   gpc1_1 gpc9353 (
      {stage2_25[110]},
      {stage3_25[39]}
   );
   gpc1_1 gpc9354 (
      {stage2_25[111]},
      {stage3_25[40]}
   );
   gpc1_1 gpc9355 (
      {stage2_25[112]},
      {stage3_25[41]}
   );
   gpc1_1 gpc9356 (
      {stage2_25[113]},
      {stage3_25[42]}
   );
   gpc1_1 gpc9357 (
      {stage2_25[114]},
      {stage3_25[43]}
   );
   gpc1_1 gpc9358 (
      {stage2_25[115]},
      {stage3_25[44]}
   );
   gpc1_1 gpc9359 (
      {stage2_25[116]},
      {stage3_25[45]}
   );
   gpc1_1 gpc9360 (
      {stage2_25[117]},
      {stage3_25[46]}
   );
   gpc1_1 gpc9361 (
      {stage2_25[118]},
      {stage3_25[47]}
   );
   gpc1_1 gpc9362 (
      {stage2_25[119]},
      {stage3_25[48]}
   );
   gpc1_1 gpc9363 (
      {stage2_25[120]},
      {stage3_25[49]}
   );
   gpc1_1 gpc9364 (
      {stage2_25[121]},
      {stage3_25[50]}
   );
   gpc1_1 gpc9365 (
      {stage2_25[122]},
      {stage3_25[51]}
   );
   gpc1_1 gpc9366 (
      {stage2_26[126]},
      {stage3_26[47]}
   );
   gpc1_1 gpc9367 (
      {stage2_26[127]},
      {stage3_26[48]}
   );
   gpc1_1 gpc9368 (
      {stage2_26[128]},
      {stage3_26[49]}
   );
   gpc1_1 gpc9369 (
      {stage2_26[129]},
      {stage3_26[50]}
   );
   gpc1_1 gpc9370 (
      {stage2_26[130]},
      {stage3_26[51]}
   );
   gpc1_1 gpc9371 (
      {stage2_28[44]},
      {stage3_28[34]}
   );
   gpc1_1 gpc9372 (
      {stage2_28[45]},
      {stage3_28[35]}
   );
   gpc1_1 gpc9373 (
      {stage2_28[46]},
      {stage3_28[36]}
   );
   gpc1_1 gpc9374 (
      {stage2_28[47]},
      {stage3_28[37]}
   );
   gpc1_1 gpc9375 (
      {stage2_28[48]},
      {stage3_28[38]}
   );
   gpc1_1 gpc9376 (
      {stage2_28[49]},
      {stage3_28[39]}
   );
   gpc1_1 gpc9377 (
      {stage2_28[50]},
      {stage3_28[40]}
   );
   gpc1_1 gpc9378 (
      {stage2_28[51]},
      {stage3_28[41]}
   );
   gpc1_1 gpc9379 (
      {stage2_28[52]},
      {stage3_28[42]}
   );
   gpc1_1 gpc9380 (
      {stage2_28[53]},
      {stage3_28[43]}
   );
   gpc1_1 gpc9381 (
      {stage2_28[54]},
      {stage3_28[44]}
   );
   gpc1_1 gpc9382 (
      {stage2_28[55]},
      {stage3_28[45]}
   );
   gpc1_1 gpc9383 (
      {stage2_28[56]},
      {stage3_28[46]}
   );
   gpc1_1 gpc9384 (
      {stage2_28[57]},
      {stage3_28[47]}
   );
   gpc1_1 gpc9385 (
      {stage2_28[58]},
      {stage3_28[48]}
   );
   gpc1_1 gpc9386 (
      {stage2_28[59]},
      {stage3_28[49]}
   );
   gpc1_1 gpc9387 (
      {stage2_28[60]},
      {stage3_28[50]}
   );
   gpc1_1 gpc9388 (
      {stage2_28[61]},
      {stage3_28[51]}
   );
   gpc1_1 gpc9389 (
      {stage2_28[62]},
      {stage3_28[52]}
   );
   gpc1_1 gpc9390 (
      {stage2_28[63]},
      {stage3_28[53]}
   );
   gpc1_1 gpc9391 (
      {stage2_28[64]},
      {stage3_28[54]}
   );
   gpc1_1 gpc9392 (
      {stage2_28[65]},
      {stage3_28[55]}
   );
   gpc1_1 gpc9393 (
      {stage2_28[66]},
      {stage3_28[56]}
   );
   gpc1_1 gpc9394 (
      {stage2_28[67]},
      {stage3_28[57]}
   );
   gpc1_1 gpc9395 (
      {stage2_28[68]},
      {stage3_28[58]}
   );
   gpc1_1 gpc9396 (
      {stage2_28[69]},
      {stage3_28[59]}
   );
   gpc1_1 gpc9397 (
      {stage2_28[70]},
      {stage3_28[60]}
   );
   gpc1_1 gpc9398 (
      {stage2_28[71]},
      {stage3_28[61]}
   );
   gpc1_1 gpc9399 (
      {stage2_28[72]},
      {stage3_28[62]}
   );
   gpc1_1 gpc9400 (
      {stage2_28[73]},
      {stage3_28[63]}
   );
   gpc1_1 gpc9401 (
      {stage2_28[74]},
      {stage3_28[64]}
   );
   gpc1_1 gpc9402 (
      {stage2_28[75]},
      {stage3_28[65]}
   );
   gpc1_1 gpc9403 (
      {stage2_28[76]},
      {stage3_28[66]}
   );
   gpc1_1 gpc9404 (
      {stage2_28[77]},
      {stage3_28[67]}
   );
   gpc1_1 gpc9405 (
      {stage2_28[78]},
      {stage3_28[68]}
   );
   gpc1_1 gpc9406 (
      {stage2_28[79]},
      {stage3_28[69]}
   );
   gpc1_1 gpc9407 (
      {stage2_29[102]},
      {stage3_29[49]}
   );
   gpc1_1 gpc9408 (
      {stage2_29[103]},
      {stage3_29[50]}
   );
   gpc1_1 gpc9409 (
      {stage2_29[104]},
      {stage3_29[51]}
   );
   gpc1_1 gpc9410 (
      {stage2_29[105]},
      {stage3_29[52]}
   );
   gpc1_1 gpc9411 (
      {stage2_29[106]},
      {stage3_29[53]}
   );
   gpc1_1 gpc9412 (
      {stage2_29[107]},
      {stage3_29[54]}
   );
   gpc1_1 gpc9413 (
      {stage2_29[108]},
      {stage3_29[55]}
   );
   gpc1_1 gpc9414 (
      {stage2_29[109]},
      {stage3_29[56]}
   );
   gpc1_1 gpc9415 (
      {stage2_29[110]},
      {stage3_29[57]}
   );
   gpc1_1 gpc9416 (
      {stage2_29[111]},
      {stage3_29[58]}
   );
   gpc1_1 gpc9417 (
      {stage2_30[93]},
      {stage3_30[32]}
   );
   gpc1_1 gpc9418 (
      {stage2_30[94]},
      {stage3_30[33]}
   );
   gpc1_1 gpc9419 (
      {stage2_30[95]},
      {stage3_30[34]}
   );
   gpc1_1 gpc9420 (
      {stage2_30[96]},
      {stage3_30[35]}
   );
   gpc1_1 gpc9421 (
      {stage2_30[97]},
      {stage3_30[36]}
   );
   gpc1_1 gpc9422 (
      {stage2_30[98]},
      {stage3_30[37]}
   );
   gpc1_1 gpc9423 (
      {stage2_30[99]},
      {stage3_30[38]}
   );
   gpc1_1 gpc9424 (
      {stage2_31[124]},
      {stage3_31[38]}
   );
   gpc1_1 gpc9425 (
      {stage2_31[125]},
      {stage3_31[39]}
   );
   gpc1_1 gpc9426 (
      {stage2_31[126]},
      {stage3_31[40]}
   );
   gpc1_1 gpc9427 (
      {stage2_31[127]},
      {stage3_31[41]}
   );
   gpc1_1 gpc9428 (
      {stage2_32[112]},
      {stage3_32[50]}
   );
   gpc1_1 gpc9429 (
      {stage2_32[113]},
      {stage3_32[51]}
   );
   gpc1_1 gpc9430 (
      {stage2_32[114]},
      {stage3_32[52]}
   );
   gpc1_1 gpc9431 (
      {stage2_32[115]},
      {stage3_32[53]}
   );
   gpc1_1 gpc9432 (
      {stage2_32[116]},
      {stage3_32[54]}
   );
   gpc1_1 gpc9433 (
      {stage2_32[117]},
      {stage3_32[55]}
   );
   gpc1_1 gpc9434 (
      {stage2_33[91]},
      {stage3_33[45]}
   );
   gpc1_1 gpc9435 (
      {stage2_33[92]},
      {stage3_33[46]}
   );
   gpc1_1 gpc9436 (
      {stage2_33[93]},
      {stage3_33[47]}
   );
   gpc1_1 gpc9437 (
      {stage2_33[94]},
      {stage3_33[48]}
   );
   gpc1_1 gpc9438 (
      {stage2_33[95]},
      {stage3_33[49]}
   );
   gpc1_1 gpc9439 (
      {stage2_33[96]},
      {stage3_33[50]}
   );
   gpc1_1 gpc9440 (
      {stage2_33[97]},
      {stage3_33[51]}
   );
   gpc1_1 gpc9441 (
      {stage2_33[98]},
      {stage3_33[52]}
   );
   gpc1_1 gpc9442 (
      {stage2_33[99]},
      {stage3_33[53]}
   );
   gpc1_1 gpc9443 (
      {stage2_33[100]},
      {stage3_33[54]}
   );
   gpc1_1 gpc9444 (
      {stage2_33[101]},
      {stage3_33[55]}
   );
   gpc1_1 gpc9445 (
      {stage2_33[102]},
      {stage3_33[56]}
   );
   gpc1_1 gpc9446 (
      {stage2_33[103]},
      {stage3_33[57]}
   );
   gpc1_1 gpc9447 (
      {stage2_33[104]},
      {stage3_33[58]}
   );
   gpc1_1 gpc9448 (
      {stage2_33[105]},
      {stage3_33[59]}
   );
   gpc1_1 gpc9449 (
      {stage2_33[106]},
      {stage3_33[60]}
   );
   gpc1_1 gpc9450 (
      {stage2_33[107]},
      {stage3_33[61]}
   );
   gpc1_1 gpc9451 (
      {stage2_33[108]},
      {stage3_33[62]}
   );
   gpc1_1 gpc9452 (
      {stage2_36[114]},
      {stage3_36[50]}
   );
   gpc1_1 gpc9453 (
      {stage2_36[115]},
      {stage3_36[51]}
   );
   gpc1_1 gpc9454 (
      {stage2_36[116]},
      {stage3_36[52]}
   );
   gpc1_1 gpc9455 (
      {stage2_36[117]},
      {stage3_36[53]}
   );
   gpc1_1 gpc9456 (
      {stage2_36[118]},
      {stage3_36[54]}
   );
   gpc1_1 gpc9457 (
      {stage2_36[119]},
      {stage3_36[55]}
   );
   gpc1_1 gpc9458 (
      {stage2_38[81]},
      {stage3_38[50]}
   );
   gpc1_1 gpc9459 (
      {stage2_38[82]},
      {stage3_38[51]}
   );
   gpc1_1 gpc9460 (
      {stage2_38[83]},
      {stage3_38[52]}
   );
   gpc1_1 gpc9461 (
      {stage2_38[84]},
      {stage3_38[53]}
   );
   gpc1_1 gpc9462 (
      {stage2_38[85]},
      {stage3_38[54]}
   );
   gpc1_1 gpc9463 (
      {stage2_38[86]},
      {stage3_38[55]}
   );
   gpc1_1 gpc9464 (
      {stage2_38[87]},
      {stage3_38[56]}
   );
   gpc1_1 gpc9465 (
      {stage2_38[88]},
      {stage3_38[57]}
   );
   gpc1_1 gpc9466 (
      {stage2_38[89]},
      {stage3_38[58]}
   );
   gpc1_1 gpc9467 (
      {stage2_38[90]},
      {stage3_38[59]}
   );
   gpc1_1 gpc9468 (
      {stage2_38[91]},
      {stage3_38[60]}
   );
   gpc1_1 gpc9469 (
      {stage2_38[92]},
      {stage3_38[61]}
   );
   gpc1_1 gpc9470 (
      {stage2_38[93]},
      {stage3_38[62]}
   );
   gpc1_1 gpc9471 (
      {stage2_38[94]},
      {stage3_38[63]}
   );
   gpc1_1 gpc9472 (
      {stage2_38[95]},
      {stage3_38[64]}
   );
   gpc1_1 gpc9473 (
      {stage2_38[96]},
      {stage3_38[65]}
   );
   gpc1_1 gpc9474 (
      {stage2_38[97]},
      {stage3_38[66]}
   );
   gpc1_1 gpc9475 (
      {stage2_38[98]},
      {stage3_38[67]}
   );
   gpc1_1 gpc9476 (
      {stage2_38[99]},
      {stage3_38[68]}
   );
   gpc1_1 gpc9477 (
      {stage2_39[100]},
      {stage3_39[52]}
   );
   gpc1_1 gpc9478 (
      {stage2_39[101]},
      {stage3_39[53]}
   );
   gpc1_1 gpc9479 (
      {stage2_39[102]},
      {stage3_39[54]}
   );
   gpc1_1 gpc9480 (
      {stage2_39[103]},
      {stage3_39[55]}
   );
   gpc1_1 gpc9481 (
      {stage2_39[104]},
      {stage3_39[56]}
   );
   gpc1_1 gpc9482 (
      {stage2_39[105]},
      {stage3_39[57]}
   );
   gpc1_1 gpc9483 (
      {stage2_39[106]},
      {stage3_39[58]}
   );
   gpc1_1 gpc9484 (
      {stage2_39[107]},
      {stage3_39[59]}
   );
   gpc1_1 gpc9485 (
      {stage2_40[131]},
      {stage3_40[37]}
   );
   gpc1_1 gpc9486 (
      {stage2_40[132]},
      {stage3_40[38]}
   );
   gpc1_1 gpc9487 (
      {stage2_40[133]},
      {stage3_40[39]}
   );
   gpc1_1 gpc9488 (
      {stage2_40[134]},
      {stage3_40[40]}
   );
   gpc1_1 gpc9489 (
      {stage2_40[135]},
      {stage3_40[41]}
   );
   gpc1_1 gpc9490 (
      {stage2_40[136]},
      {stage3_40[42]}
   );
   gpc1_1 gpc9491 (
      {stage2_40[137]},
      {stage3_40[43]}
   );
   gpc1_1 gpc9492 (
      {stage2_40[138]},
      {stage3_40[44]}
   );
   gpc1_1 gpc9493 (
      {stage2_40[139]},
      {stage3_40[45]}
   );
   gpc1_1 gpc9494 (
      {stage2_41[102]},
      {stage3_41[36]}
   );
   gpc1_1 gpc9495 (
      {stage2_41[103]},
      {stage3_41[37]}
   );
   gpc1_1 gpc9496 (
      {stage2_41[104]},
      {stage3_41[38]}
   );
   gpc1_1 gpc9497 (
      {stage2_41[105]},
      {stage3_41[39]}
   );
   gpc1_1 gpc9498 (
      {stage2_41[106]},
      {stage3_41[40]}
   );
   gpc1_1 gpc9499 (
      {stage2_41[107]},
      {stage3_41[41]}
   );
   gpc1_1 gpc9500 (
      {stage2_41[108]},
      {stage3_41[42]}
   );
   gpc1_1 gpc9501 (
      {stage2_41[109]},
      {stage3_41[43]}
   );
   gpc1_1 gpc9502 (
      {stage2_41[110]},
      {stage3_41[44]}
   );
   gpc1_1 gpc9503 (
      {stage2_41[111]},
      {stage3_41[45]}
   );
   gpc1_1 gpc9504 (
      {stage2_41[112]},
      {stage3_41[46]}
   );
   gpc1_1 gpc9505 (
      {stage2_41[113]},
      {stage3_41[47]}
   );
   gpc1_1 gpc9506 (
      {stage2_41[114]},
      {stage3_41[48]}
   );
   gpc1_1 gpc9507 (
      {stage2_41[115]},
      {stage3_41[49]}
   );
   gpc1_1 gpc9508 (
      {stage2_41[116]},
      {stage3_41[50]}
   );
   gpc1_1 gpc9509 (
      {stage2_41[117]},
      {stage3_41[51]}
   );
   gpc1_1 gpc9510 (
      {stage2_41[118]},
      {stage3_41[52]}
   );
   gpc1_1 gpc9511 (
      {stage2_41[119]},
      {stage3_41[53]}
   );
   gpc1_1 gpc9512 (
      {stage2_41[120]},
      {stage3_41[54]}
   );
   gpc1_1 gpc9513 (
      {stage2_41[121]},
      {stage3_41[55]}
   );
   gpc1_1 gpc9514 (
      {stage2_41[122]},
      {stage3_41[56]}
   );
   gpc1_1 gpc9515 (
      {stage2_42[74]},
      {stage3_42[46]}
   );
   gpc1_1 gpc9516 (
      {stage2_42[75]},
      {stage3_42[47]}
   );
   gpc1_1 gpc9517 (
      {stage2_42[76]},
      {stage3_42[48]}
   );
   gpc1_1 gpc9518 (
      {stage2_42[77]},
      {stage3_42[49]}
   );
   gpc1_1 gpc9519 (
      {stage2_42[78]},
      {stage3_42[50]}
   );
   gpc1_1 gpc9520 (
      {stage2_42[79]},
      {stage3_42[51]}
   );
   gpc1_1 gpc9521 (
      {stage2_42[80]},
      {stage3_42[52]}
   );
   gpc1_1 gpc9522 (
      {stage2_42[81]},
      {stage3_42[53]}
   );
   gpc1_1 gpc9523 (
      {stage2_43[98]},
      {stage3_43[47]}
   );
   gpc1_1 gpc9524 (
      {stage2_43[99]},
      {stage3_43[48]}
   );
   gpc1_1 gpc9525 (
      {stage2_43[100]},
      {stage3_43[49]}
   );
   gpc1_1 gpc9526 (
      {stage2_43[101]},
      {stage3_43[50]}
   );
   gpc1_1 gpc9527 (
      {stage2_43[102]},
      {stage3_43[51]}
   );
   gpc1_1 gpc9528 (
      {stage2_43[103]},
      {stage3_43[52]}
   );
   gpc1_1 gpc9529 (
      {stage2_43[104]},
      {stage3_43[53]}
   );
   gpc1_1 gpc9530 (
      {stage2_43[105]},
      {stage3_43[54]}
   );
   gpc1_1 gpc9531 (
      {stage2_43[106]},
      {stage3_43[55]}
   );
   gpc1_1 gpc9532 (
      {stage2_43[107]},
      {stage3_43[56]}
   );
   gpc1_1 gpc9533 (
      {stage2_43[108]},
      {stage3_43[57]}
   );
   gpc1_1 gpc9534 (
      {stage2_43[109]},
      {stage3_43[58]}
   );
   gpc1_1 gpc9535 (
      {stage2_43[110]},
      {stage3_43[59]}
   );
   gpc1_1 gpc9536 (
      {stage2_44[86]},
      {stage3_44[33]}
   );
   gpc1_1 gpc9537 (
      {stage2_44[87]},
      {stage3_44[34]}
   );
   gpc1_1 gpc9538 (
      {stage2_44[88]},
      {stage3_44[35]}
   );
   gpc1_1 gpc9539 (
      {stage2_44[89]},
      {stage3_44[36]}
   );
   gpc1_1 gpc9540 (
      {stage2_44[90]},
      {stage3_44[37]}
   );
   gpc1_1 gpc9541 (
      {stage2_44[91]},
      {stage3_44[38]}
   );
   gpc1_1 gpc9542 (
      {stage2_44[92]},
      {stage3_44[39]}
   );
   gpc1_1 gpc9543 (
      {stage2_44[93]},
      {stage3_44[40]}
   );
   gpc1_1 gpc9544 (
      {stage2_44[94]},
      {stage3_44[41]}
   );
   gpc1_1 gpc9545 (
      {stage2_44[95]},
      {stage3_44[42]}
   );
   gpc1_1 gpc9546 (
      {stage2_44[96]},
      {stage3_44[43]}
   );
   gpc1_1 gpc9547 (
      {stage2_44[97]},
      {stage3_44[44]}
   );
   gpc1_1 gpc9548 (
      {stage2_44[98]},
      {stage3_44[45]}
   );
   gpc1_1 gpc9549 (
      {stage2_44[99]},
      {stage3_44[46]}
   );
   gpc1_1 gpc9550 (
      {stage2_44[100]},
      {stage3_44[47]}
   );
   gpc1_1 gpc9551 (
      {stage2_44[101]},
      {stage3_44[48]}
   );
   gpc1_1 gpc9552 (
      {stage2_44[102]},
      {stage3_44[49]}
   );
   gpc1_1 gpc9553 (
      {stage2_44[103]},
      {stage3_44[50]}
   );
   gpc1_1 gpc9554 (
      {stage2_44[104]},
      {stage3_44[51]}
   );
   gpc1_1 gpc9555 (
      {stage2_44[105]},
      {stage3_44[52]}
   );
   gpc1_1 gpc9556 (
      {stage2_44[106]},
      {stage3_44[53]}
   );
   gpc1_1 gpc9557 (
      {stage2_44[107]},
      {stage3_44[54]}
   );
   gpc1_1 gpc9558 (
      {stage2_44[108]},
      {stage3_44[55]}
   );
   gpc1_1 gpc9559 (
      {stage2_44[109]},
      {stage3_44[56]}
   );
   gpc1_1 gpc9560 (
      {stage2_44[110]},
      {stage3_44[57]}
   );
   gpc1_1 gpc9561 (
      {stage2_44[111]},
      {stage3_44[58]}
   );
   gpc1_1 gpc9562 (
      {stage2_44[112]},
      {stage3_44[59]}
   );
   gpc1_1 gpc9563 (
      {stage2_44[113]},
      {stage3_44[60]}
   );
   gpc1_1 gpc9564 (
      {stage2_44[114]},
      {stage3_44[61]}
   );
   gpc1_1 gpc9565 (
      {stage2_44[115]},
      {stage3_44[62]}
   );
   gpc1_1 gpc9566 (
      {stage2_44[116]},
      {stage3_44[63]}
   );
   gpc1_1 gpc9567 (
      {stage2_44[117]},
      {stage3_44[64]}
   );
   gpc1_1 gpc9568 (
      {stage2_44[118]},
      {stage3_44[65]}
   );
   gpc1_1 gpc9569 (
      {stage2_44[119]},
      {stage3_44[66]}
   );
   gpc1_1 gpc9570 (
      {stage2_44[120]},
      {stage3_44[67]}
   );
   gpc1_1 gpc9571 (
      {stage2_44[121]},
      {stage3_44[68]}
   );
   gpc1_1 gpc9572 (
      {stage2_44[122]},
      {stage3_44[69]}
   );
   gpc1_1 gpc9573 (
      {stage2_44[123]},
      {stage3_44[70]}
   );
   gpc1_1 gpc9574 (
      {stage2_44[124]},
      {stage3_44[71]}
   );
   gpc1_1 gpc9575 (
      {stage2_44[125]},
      {stage3_44[72]}
   );
   gpc1_1 gpc9576 (
      {stage2_44[126]},
      {stage3_44[73]}
   );
   gpc1_1 gpc9577 (
      {stage2_44[127]},
      {stage3_44[74]}
   );
   gpc1_1 gpc9578 (
      {stage2_44[128]},
      {stage3_44[75]}
   );
   gpc1_1 gpc9579 (
      {stage2_44[129]},
      {stage3_44[76]}
   );
   gpc1_1 gpc9580 (
      {stage2_44[130]},
      {stage3_44[77]}
   );
   gpc1_1 gpc9581 (
      {stage2_44[131]},
      {stage3_44[78]}
   );
   gpc1_1 gpc9582 (
      {stage2_44[132]},
      {stage3_44[79]}
   );
   gpc1_1 gpc9583 (
      {stage2_44[133]},
      {stage3_44[80]}
   );
   gpc1_1 gpc9584 (
      {stage2_44[134]},
      {stage3_44[81]}
   );
   gpc1_1 gpc9585 (
      {stage2_44[135]},
      {stage3_44[82]}
   );
   gpc1_1 gpc9586 (
      {stage2_44[136]},
      {stage3_44[83]}
   );
   gpc1_1 gpc9587 (
      {stage2_44[137]},
      {stage3_44[84]}
   );
   gpc1_1 gpc9588 (
      {stage2_45[126]},
      {stage3_45[34]}
   );
   gpc1_1 gpc9589 (
      {stage2_45[127]},
      {stage3_45[35]}
   );
   gpc1_1 gpc9590 (
      {stage2_45[128]},
      {stage3_45[36]}
   );
   gpc1_1 gpc9591 (
      {stage2_45[129]},
      {stage3_45[37]}
   );
   gpc1_1 gpc9592 (
      {stage2_45[130]},
      {stage3_45[38]}
   );
   gpc1_1 gpc9593 (
      {stage2_45[131]},
      {stage3_45[39]}
   );
   gpc1_1 gpc9594 (
      {stage2_47[83]},
      {stage3_47[49]}
   );
   gpc1_1 gpc9595 (
      {stage2_47[84]},
      {stage3_47[50]}
   );
   gpc1_1 gpc9596 (
      {stage2_47[85]},
      {stage3_47[51]}
   );
   gpc1_1 gpc9597 (
      {stage2_47[86]},
      {stage3_47[52]}
   );
   gpc1_1 gpc9598 (
      {stage2_47[87]},
      {stage3_47[53]}
   );
   gpc1_1 gpc9599 (
      {stage2_47[88]},
      {stage3_47[54]}
   );
   gpc1_1 gpc9600 (
      {stage2_47[89]},
      {stage3_47[55]}
   );
   gpc1_1 gpc9601 (
      {stage2_47[90]},
      {stage3_47[56]}
   );
   gpc1_1 gpc9602 (
      {stage2_47[91]},
      {stage3_47[57]}
   );
   gpc1_1 gpc9603 (
      {stage2_47[92]},
      {stage3_47[58]}
   );
   gpc1_1 gpc9604 (
      {stage2_47[93]},
      {stage3_47[59]}
   );
   gpc1_1 gpc9605 (
      {stage2_47[94]},
      {stage3_47[60]}
   );
   gpc1_1 gpc9606 (
      {stage2_47[95]},
      {stage3_47[61]}
   );
   gpc1_1 gpc9607 (
      {stage2_47[96]},
      {stage3_47[62]}
   );
   gpc1_1 gpc9608 (
      {stage2_47[97]},
      {stage3_47[63]}
   );
   gpc1_1 gpc9609 (
      {stage2_47[98]},
      {stage3_47[64]}
   );
   gpc1_1 gpc9610 (
      {stage2_47[99]},
      {stage3_47[65]}
   );
   gpc1_1 gpc9611 (
      {stage2_47[100]},
      {stage3_47[66]}
   );
   gpc1_1 gpc9612 (
      {stage2_47[101]},
      {stage3_47[67]}
   );
   gpc1_1 gpc9613 (
      {stage2_47[102]},
      {stage3_47[68]}
   );
   gpc1_1 gpc9614 (
      {stage2_47[103]},
      {stage3_47[69]}
   );
   gpc1_1 gpc9615 (
      {stage2_47[104]},
      {stage3_47[70]}
   );
   gpc1_1 gpc9616 (
      {stage2_47[105]},
      {stage3_47[71]}
   );
   gpc1_1 gpc9617 (
      {stage2_47[106]},
      {stage3_47[72]}
   );
   gpc1_1 gpc9618 (
      {stage2_47[107]},
      {stage3_47[73]}
   );
   gpc1_1 gpc9619 (
      {stage2_49[96]},
      {stage3_49[45]}
   );
   gpc1_1 gpc9620 (
      {stage2_49[97]},
      {stage3_49[46]}
   );
   gpc1_1 gpc9621 (
      {stage2_49[98]},
      {stage3_49[47]}
   );
   gpc1_1 gpc9622 (
      {stage2_49[99]},
      {stage3_49[48]}
   );
   gpc1_1 gpc9623 (
      {stage2_49[100]},
      {stage3_49[49]}
   );
   gpc1_1 gpc9624 (
      {stage2_49[101]},
      {stage3_49[50]}
   );
   gpc1_1 gpc9625 (
      {stage2_49[102]},
      {stage3_49[51]}
   );
   gpc1_1 gpc9626 (
      {stage2_49[103]},
      {stage3_49[52]}
   );
   gpc1_1 gpc9627 (
      {stage2_49[104]},
      {stage3_49[53]}
   );
   gpc1_1 gpc9628 (
      {stage2_49[105]},
      {stage3_49[54]}
   );
   gpc1_1 gpc9629 (
      {stage2_49[106]},
      {stage3_49[55]}
   );
   gpc1_1 gpc9630 (
      {stage2_49[107]},
      {stage3_49[56]}
   );
   gpc1_1 gpc9631 (
      {stage2_49[108]},
      {stage3_49[57]}
   );
   gpc1_1 gpc9632 (
      {stage2_49[109]},
      {stage3_49[58]}
   );
   gpc1_1 gpc9633 (
      {stage2_49[110]},
      {stage3_49[59]}
   );
   gpc1_1 gpc9634 (
      {stage2_49[111]},
      {stage3_49[60]}
   );
   gpc1_1 gpc9635 (
      {stage2_49[112]},
      {stage3_49[61]}
   );
   gpc1_1 gpc9636 (
      {stage2_49[113]},
      {stage3_49[62]}
   );
   gpc1_1 gpc9637 (
      {stage2_49[114]},
      {stage3_49[63]}
   );
   gpc1_1 gpc9638 (
      {stage2_49[115]},
      {stage3_49[64]}
   );
   gpc1_1 gpc9639 (
      {stage2_50[149]},
      {stage3_50[60]}
   );
   gpc1_1 gpc9640 (
      {stage2_50[150]},
      {stage3_50[61]}
   );
   gpc1_1 gpc9641 (
      {stage2_50[151]},
      {stage3_50[62]}
   );
   gpc1_1 gpc9642 (
      {stage2_50[152]},
      {stage3_50[63]}
   );
   gpc1_1 gpc9643 (
      {stage2_51[81]},
      {stage3_51[47]}
   );
   gpc1_1 gpc9644 (
      {stage2_51[82]},
      {stage3_51[48]}
   );
   gpc1_1 gpc9645 (
      {stage2_51[83]},
      {stage3_51[49]}
   );
   gpc1_1 gpc9646 (
      {stage2_51[84]},
      {stage3_51[50]}
   );
   gpc1_1 gpc9647 (
      {stage2_51[85]},
      {stage3_51[51]}
   );
   gpc1_1 gpc9648 (
      {stage2_51[86]},
      {stage3_51[52]}
   );
   gpc1_1 gpc9649 (
      {stage2_51[87]},
      {stage3_51[53]}
   );
   gpc1_1 gpc9650 (
      {stage2_52[109]},
      {stage3_52[37]}
   );
   gpc1_1 gpc9651 (
      {stage2_52[110]},
      {stage3_52[38]}
   );
   gpc1_1 gpc9652 (
      {stage2_52[111]},
      {stage3_52[39]}
   );
   gpc1_1 gpc9653 (
      {stage2_52[112]},
      {stage3_52[40]}
   );
   gpc1_1 gpc9654 (
      {stage2_52[113]},
      {stage3_52[41]}
   );
   gpc1_1 gpc9655 (
      {stage2_52[114]},
      {stage3_52[42]}
   );
   gpc1_1 gpc9656 (
      {stage2_52[115]},
      {stage3_52[43]}
   );
   gpc1_1 gpc9657 (
      {stage2_52[116]},
      {stage3_52[44]}
   );
   gpc1_1 gpc9658 (
      {stage2_52[117]},
      {stage3_52[45]}
   );
   gpc1_1 gpc9659 (
      {stage2_52[118]},
      {stage3_52[46]}
   );
   gpc1_1 gpc9660 (
      {stage2_52[119]},
      {stage3_52[47]}
   );
   gpc1_1 gpc9661 (
      {stage2_52[120]},
      {stage3_52[48]}
   );
   gpc1_1 gpc9662 (
      {stage2_52[121]},
      {stage3_52[49]}
   );
   gpc1_1 gpc9663 (
      {stage2_52[122]},
      {stage3_52[50]}
   );
   gpc1_1 gpc9664 (
      {stage2_52[123]},
      {stage3_52[51]}
   );
   gpc1_1 gpc9665 (
      {stage2_52[124]},
      {stage3_52[52]}
   );
   gpc1_1 gpc9666 (
      {stage2_52[125]},
      {stage3_52[53]}
   );
   gpc1_1 gpc9667 (
      {stage2_52[126]},
      {stage3_52[54]}
   );
   gpc1_1 gpc9668 (
      {stage2_52[127]},
      {stage3_52[55]}
   );
   gpc1_1 gpc9669 (
      {stage2_53[89]},
      {stage3_53[45]}
   );
   gpc1_1 gpc9670 (
      {stage2_53[90]},
      {stage3_53[46]}
   );
   gpc1_1 gpc9671 (
      {stage2_53[91]},
      {stage3_53[47]}
   );
   gpc1_1 gpc9672 (
      {stage2_53[92]},
      {stage3_53[48]}
   );
   gpc1_1 gpc9673 (
      {stage2_53[93]},
      {stage3_53[49]}
   );
   gpc1_1 gpc9674 (
      {stage2_53[94]},
      {stage3_53[50]}
   );
   gpc1_1 gpc9675 (
      {stage2_53[95]},
      {stage3_53[51]}
   );
   gpc1_1 gpc9676 (
      {stage2_53[96]},
      {stage3_53[52]}
   );
   gpc1_1 gpc9677 (
      {stage2_54[114]},
      {stage3_54[53]}
   );
   gpc1_1 gpc9678 (
      {stage2_54[115]},
      {stage3_54[54]}
   );
   gpc1_1 gpc9679 (
      {stage2_54[116]},
      {stage3_54[55]}
   );
   gpc1_1 gpc9680 (
      {stage2_54[117]},
      {stage3_54[56]}
   );
   gpc1_1 gpc9681 (
      {stage2_54[118]},
      {stage3_54[57]}
   );
   gpc1_1 gpc9682 (
      {stage2_54[119]},
      {stage3_54[58]}
   );
   gpc1_1 gpc9683 (
      {stage2_54[120]},
      {stage3_54[59]}
   );
   gpc1_1 gpc9684 (
      {stage2_54[121]},
      {stage3_54[60]}
   );
   gpc1_1 gpc9685 (
      {stage2_54[122]},
      {stage3_54[61]}
   );
   gpc1_1 gpc9686 (
      {stage2_54[123]},
      {stage3_54[62]}
   );
   gpc1_1 gpc9687 (
      {stage2_55[102]},
      {stage3_55[38]}
   );
   gpc1_1 gpc9688 (
      {stage2_55[103]},
      {stage3_55[39]}
   );
   gpc1_1 gpc9689 (
      {stage2_55[104]},
      {stage3_55[40]}
   );
   gpc1_1 gpc9690 (
      {stage2_55[105]},
      {stage3_55[41]}
   );
   gpc1_1 gpc9691 (
      {stage2_55[106]},
      {stage3_55[42]}
   );
   gpc1_1 gpc9692 (
      {stage2_55[107]},
      {stage3_55[43]}
   );
   gpc1_1 gpc9693 (
      {stage2_55[108]},
      {stage3_55[44]}
   );
   gpc1_1 gpc9694 (
      {stage2_55[109]},
      {stage3_55[45]}
   );
   gpc1_1 gpc9695 (
      {stage2_55[110]},
      {stage3_55[46]}
   );
   gpc1_1 gpc9696 (
      {stage2_57[72]},
      {stage3_57[46]}
   );
   gpc1_1 gpc9697 (
      {stage2_57[73]},
      {stage3_57[47]}
   );
   gpc1_1 gpc9698 (
      {stage2_57[74]},
      {stage3_57[48]}
   );
   gpc1_1 gpc9699 (
      {stage2_57[75]},
      {stage3_57[49]}
   );
   gpc1_1 gpc9700 (
      {stage2_57[76]},
      {stage3_57[50]}
   );
   gpc1_1 gpc9701 (
      {stage2_57[77]},
      {stage3_57[51]}
   );
   gpc1_1 gpc9702 (
      {stage2_57[78]},
      {stage3_57[52]}
   );
   gpc1_1 gpc9703 (
      {stage2_58[79]},
      {stage3_58[43]}
   );
   gpc1_1 gpc9704 (
      {stage2_58[80]},
      {stage3_58[44]}
   );
   gpc1_1 gpc9705 (
      {stage2_58[81]},
      {stage3_58[45]}
   );
   gpc1_1 gpc9706 (
      {stage2_58[82]},
      {stage3_58[46]}
   );
   gpc1_1 gpc9707 (
      {stage2_58[83]},
      {stage3_58[47]}
   );
   gpc1_1 gpc9708 (
      {stage2_58[84]},
      {stage3_58[48]}
   );
   gpc1_1 gpc9709 (
      {stage2_59[133]},
      {stage3_59[39]}
   );
   gpc1_1 gpc9710 (
      {stage2_59[134]},
      {stage3_59[40]}
   );
   gpc1_1 gpc9711 (
      {stage2_59[135]},
      {stage3_59[41]}
   );
   gpc1_1 gpc9712 (
      {stage2_59[136]},
      {stage3_59[42]}
   );
   gpc1_1 gpc9713 (
      {stage2_59[137]},
      {stage3_59[43]}
   );
   gpc1_1 gpc9714 (
      {stage2_59[138]},
      {stage3_59[44]}
   );
   gpc1_1 gpc9715 (
      {stage2_59[139]},
      {stage3_59[45]}
   );
   gpc1_1 gpc9716 (
      {stage2_60[106]},
      {stage3_60[48]}
   );
   gpc1_1 gpc9717 (
      {stage2_60[107]},
      {stage3_60[49]}
   );
   gpc1_1 gpc9718 (
      {stage2_60[108]},
      {stage3_60[50]}
   );
   gpc1_1 gpc9719 (
      {stage2_60[109]},
      {stage3_60[51]}
   );
   gpc1_1 gpc9720 (
      {stage2_60[110]},
      {stage3_60[52]}
   );
   gpc1_1 gpc9721 (
      {stage2_61[90]},
      {stage3_61[45]}
   );
   gpc1_1 gpc9722 (
      {stage2_61[91]},
      {stage3_61[46]}
   );
   gpc1_1 gpc9723 (
      {stage2_61[92]},
      {stage3_61[47]}
   );
   gpc1_1 gpc9724 (
      {stage2_61[93]},
      {stage3_61[48]}
   );
   gpc1_1 gpc9725 (
      {stage2_61[94]},
      {stage3_61[49]}
   );
   gpc1_1 gpc9726 (
      {stage2_61[95]},
      {stage3_61[50]}
   );
   gpc1_1 gpc9727 (
      {stage2_61[96]},
      {stage3_61[51]}
   );
   gpc1_1 gpc9728 (
      {stage2_61[97]},
      {stage3_61[52]}
   );
   gpc1_1 gpc9729 (
      {stage2_61[98]},
      {stage3_61[53]}
   );
   gpc1_1 gpc9730 (
      {stage2_61[99]},
      {stage3_61[54]}
   );
   gpc1_1 gpc9731 (
      {stage2_61[100]},
      {stage3_61[55]}
   );
   gpc1_1 gpc9732 (
      {stage2_61[101]},
      {stage3_61[56]}
   );
   gpc1_1 gpc9733 (
      {stage2_62[144]},
      {stage3_62[40]}
   );
   gpc1_1 gpc9734 (
      {stage2_63[95]},
      {stage3_63[54]}
   );
   gpc1_1 gpc9735 (
      {stage2_63[96]},
      {stage3_63[55]}
   );
   gpc1_1 gpc9736 (
      {stage2_63[97]},
      {stage3_63[56]}
   );
   gpc1_1 gpc9737 (
      {stage2_63[98]},
      {stage3_63[57]}
   );
   gpc1_1 gpc9738 (
      {stage2_63[99]},
      {stage3_63[58]}
   );
   gpc1_1 gpc9739 (
      {stage2_63[100]},
      {stage3_63[59]}
   );
   gpc1_1 gpc9740 (
      {stage2_63[101]},
      {stage3_63[60]}
   );
   gpc1_1 gpc9741 (
      {stage2_63[102]},
      {stage3_63[61]}
   );
   gpc1_1 gpc9742 (
      {stage2_63[103]},
      {stage3_63[62]}
   );
   gpc1_1 gpc9743 (
      {stage2_63[104]},
      {stage3_63[63]}
   );
   gpc1_1 gpc9744 (
      {stage2_63[105]},
      {stage3_63[64]}
   );
   gpc1_1 gpc9745 (
      {stage2_63[106]},
      {stage3_63[65]}
   );
   gpc1_1 gpc9746 (
      {stage2_63[107]},
      {stage3_63[66]}
   );
   gpc1_1 gpc9747 (
      {stage2_63[108]},
      {stage3_63[67]}
   );
   gpc1_1 gpc9748 (
      {stage2_63[109]},
      {stage3_63[68]}
   );
   gpc1_1 gpc9749 (
      {stage2_63[110]},
      {stage3_63[69]}
   );
   gpc1_1 gpc9750 (
      {stage2_63[111]},
      {stage3_63[70]}
   );
   gpc1_1 gpc9751 (
      {stage2_63[112]},
      {stage3_63[71]}
   );
   gpc1_1 gpc9752 (
      {stage2_64[95]},
      {stage3_64[44]}
   );
   gpc1_1 gpc9753 (
      {stage2_64[96]},
      {stage3_64[45]}
   );
   gpc1_1 gpc9754 (
      {stage2_64[97]},
      {stage3_64[46]}
   );
   gpc1_1 gpc9755 (
      {stage2_64[98]},
      {stage3_64[47]}
   );
   gpc1_1 gpc9756 (
      {stage2_64[99]},
      {stage3_64[48]}
   );
   gpc1_1 gpc9757 (
      {stage2_64[100]},
      {stage3_64[49]}
   );
   gpc1_1 gpc9758 (
      {stage2_64[101]},
      {stage3_64[50]}
   );
   gpc1_1 gpc9759 (
      {stage2_65[65]},
      {stage3_65[30]}
   );
   gpc1_1 gpc9760 (
      {stage2_65[66]},
      {stage3_65[31]}
   );
   gpc1_1 gpc9761 (
      {stage2_65[67]},
      {stage3_65[32]}
   );
   gpc1_1 gpc9762 (
      {stage2_66[30]},
      {stage3_66[30]}
   );
   gpc1_1 gpc9763 (
      {stage2_66[31]},
      {stage3_66[31]}
   );
   gpc1_1 gpc9764 (
      {stage2_66[32]},
      {stage3_66[32]}
   );
   gpc1_1 gpc9765 (
      {stage2_66[33]},
      {stage3_66[33]}
   );
   gpc1_1 gpc9766 (
      {stage2_66[34]},
      {stage3_66[34]}
   );
   gpc1_1 gpc9767 (
      {stage2_66[35]},
      {stage3_66[35]}
   );
   gpc1_1 gpc9768 (
      {stage2_66[36]},
      {stage3_66[36]}
   );
   gpc1_1 gpc9769 (
      {stage2_66[37]},
      {stage3_66[37]}
   );
   gpc1_1 gpc9770 (
      {stage2_66[38]},
      {stage3_66[38]}
   );
   gpc1_1 gpc9771 (
      {stage2_66[39]},
      {stage3_66[39]}
   );
   gpc1_1 gpc9772 (
      {stage2_66[40]},
      {stage3_66[40]}
   );
   gpc1_1 gpc9773 (
      {stage2_66[41]},
      {stage3_66[41]}
   );
   gpc1_1 gpc9774 (
      {stage2_66[42]},
      {stage3_66[42]}
   );
   gpc1_1 gpc9775 (
      {stage2_66[43]},
      {stage3_66[43]}
   );
   gpc1_1 gpc9776 (
      {stage2_66[44]},
      {stage3_66[44]}
   );
   gpc1_1 gpc9777 (
      {stage2_66[45]},
      {stage3_66[45]}
   );
   gpc1_1 gpc9778 (
      {stage2_66[46]},
      {stage3_66[46]}
   );
   gpc1_1 gpc9779 (
      {stage2_66[47]},
      {stage3_66[47]}
   );
   gpc1_1 gpc9780 (
      {stage2_66[48]},
      {stage3_66[48]}
   );
   gpc1_1 gpc9781 (
      {stage2_66[49]},
      {stage3_66[49]}
   );
   gpc1_1 gpc9782 (
      {stage2_66[50]},
      {stage3_66[50]}
   );
   gpc1_1 gpc9783 (
      {stage2_66[51]},
      {stage3_66[51]}
   );
   gpc1_1 gpc9784 (
      {stage2_66[52]},
      {stage3_66[52]}
   );
   gpc1_1 gpc9785 (
      {stage2_66[53]},
      {stage3_66[53]}
   );
   gpc606_5 gpc9786 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc9787 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc9788 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc9789 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc9790 (
      {stage3_1[18], stage3_1[19], stage3_1[20], stage3_1[21], stage3_1[22], stage3_1[23]},
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc9791 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc9792 (
      {stage3_3[24], stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc9793 (
      {stage3_3[29], stage3_3[30], stage3_3[31], stage3_3[32], stage3_3[33]},
      {stage3_4[7]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc9794 (
      {stage3_3[34], stage3_3[35], stage3_3[36], stage3_3[37], stage3_3[38]},
      {stage3_4[8]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[3],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc9795 (
      {stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[4],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc9796 (
      {stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[5],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc9797 (
      {stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[5],stage4_6[6],stage4_5[10],stage4_4[11]}
   );
   gpc606_5 gpc9798 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[3],stage4_7[6],stage4_6[7],stage4_5[11],stage4_4[12]}
   );
   gpc606_5 gpc9799 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[4],stage4_7[7],stage4_6[8],stage4_5[12],stage4_4[13]}
   );
   gpc606_5 gpc9800 (
      {stage3_4[39], stage3_4[40], stage3_4[41], stage3_4[42], stage3_4[43], stage3_4[44]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[5],stage4_7[8],stage4_6[9],stage4_5[13],stage4_4[14]}
   );
   gpc606_5 gpc9801 (
      {stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48], stage3_4[49], stage3_4[50]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[6],stage4_7[9],stage4_6[10],stage4_5[14],stage4_4[15]}
   );
   gpc606_5 gpc9802 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[7],stage4_7[10],stage4_6[11],stage4_5[15]}
   );
   gpc615_5 gpc9803 (
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[8],stage4_7[11],stage4_6[12]}
   );
   gpc615_5 gpc9804 (
      {stage3_6[47], stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[9],stage4_7[12],stage4_6[13]}
   );
   gpc615_5 gpc9805 (
      {stage3_6[52], stage3_6[53], stage3_6[54], stage3_6[55], stage3_6[56]},
      {stage3_7[8]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[10],stage4_7[13],stage4_6[14]}
   );
   gpc615_5 gpc9806 (
      {stage3_6[57], stage3_6[58], stage3_6[59], stage3_6[60], stage3_6[61]},
      {stage3_7[9]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[4],stage4_8[11],stage4_7[14],stage4_6[15]}
   );
   gpc615_5 gpc9807 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[24]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[4],stage4_9[5],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc9808 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[25]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[5],stage4_9[6],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc9809 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[26]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[6],stage4_9[7],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc9810 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[27]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[7],stage4_9[8],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc9811 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[28]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[8],stage4_9[9],stage4_8[16],stage4_7[19]}
   );
   gpc606_5 gpc9812 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[5],stage4_10[9],stage4_9[10]}
   );
   gpc606_5 gpc9813 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[6],stage4_10[10],stage4_9[11]}
   );
   gpc606_5 gpc9814 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[7],stage4_10[11],stage4_9[12]}
   );
   gpc606_5 gpc9815 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], 1'b0},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[8],stage4_10[12],stage4_9[13]}
   );
   gpc615_5 gpc9816 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[24]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[4],stage4_12[4],stage4_11[9],stage4_10[13]}
   );
   gpc615_5 gpc9817 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[25]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[5],stage4_12[5],stage4_11[10],stage4_10[14]}
   );
   gpc615_5 gpc9818 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[26]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[6],stage4_12[6],stage4_11[11],stage4_10[15]}
   );
   gpc615_5 gpc9819 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[27]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[7],stage4_12[7],stage4_11[12],stage4_10[16]}
   );
   gpc615_5 gpc9820 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24]},
      {stage3_11[28]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[8],stage4_12[8],stage4_11[13],stage4_10[17]}
   );
   gpc615_5 gpc9821 (
      {stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29]},
      {stage3_11[29]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[9],stage4_12[9],stage4_11[14],stage4_10[18]}
   );
   gpc615_5 gpc9822 (
      {stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33], stage3_10[34]},
      {stage3_11[30]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[10],stage4_12[10],stage4_11[15],stage4_10[19]}
   );
   gpc615_5 gpc9823 (
      {stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38], stage3_10[39]},
      {stage3_11[31]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[11],stage4_12[11],stage4_11[16],stage4_10[20]}
   );
   gpc615_5 gpc9824 (
      {stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43], stage3_10[44]},
      {stage3_11[32]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[12],stage4_12[12],stage4_11[17],stage4_10[21]}
   );
   gpc615_5 gpc9825 (
      {stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48], stage3_10[49]},
      {stage3_11[33]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[13],stage4_12[13],stage4_11[18],stage4_10[22]}
   );
   gpc615_5 gpc9826 (
      {stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53], stage3_10[54]},
      {stage3_11[34]},
      {stage3_12[60], stage3_12[61], stage3_12[62], stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage4_14[10],stage4_13[14],stage4_12[14],stage4_11[19],stage4_10[23]}
   );
   gpc615_5 gpc9827 (
      {stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58], stage3_10[59]},
      {stage3_11[35]},
      {stage3_12[66], stage3_12[67], stage3_12[68], stage3_12[69], stage3_12[70], stage3_12[71]},
      {stage4_14[11],stage4_13[15],stage4_12[15],stage4_11[20],stage4_10[24]}
   );
   gpc615_5 gpc9828 (
      {stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63], stage3_10[64]},
      {stage3_11[36]},
      {stage3_12[72], stage3_12[73], stage3_12[74], stage3_12[75], stage3_12[76], stage3_12[77]},
      {stage4_14[12],stage4_13[16],stage4_12[16],stage4_11[21],stage4_10[25]}
   );
   gpc615_5 gpc9829 (
      {stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[78]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[13],stage4_13[17],stage4_12[17],stage4_11[22]}
   );
   gpc615_5 gpc9830 (
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46]},
      {stage3_12[79]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[14],stage4_13[18],stage4_12[18],stage4_11[23]}
   );
   gpc615_5 gpc9831 (
      {stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51]},
      {stage3_12[80]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[15],stage4_13[19],stage4_12[19],stage4_11[24]}
   );
   gpc117_4 gpc9832 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[3],stage4_14[16],stage4_13[20]}
   );
   gpc606_5 gpc9833 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6]},
      {stage4_17[0],stage4_16[1],stage4_15[4],stage4_14[17],stage4_13[21]}
   );
   gpc606_5 gpc9834 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage4_17[1],stage4_16[2],stage4_15[5],stage4_14[18],stage4_13[22]}
   );
   gpc606_5 gpc9835 (
      {stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42]},
      {stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18]},
      {stage4_17[2],stage4_16[3],stage4_15[6],stage4_14[19],stage4_13[23]}
   );
   gpc615_5 gpc9836 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_15[19]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[3],stage4_16[4],stage4_15[7],stage4_14[20]}
   );
   gpc615_5 gpc9837 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[20]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[4],stage4_16[5],stage4_15[8],stage4_14[21]}
   );
   gpc615_5 gpc9838 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[21]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[5],stage4_16[6],stage4_15[9],stage4_14[22]}
   );
   gpc615_5 gpc9839 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[22]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[6],stage4_16[7],stage4_15[10],stage4_14[23]}
   );
   gpc615_5 gpc9840 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[23]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[7],stage4_16[8],stage4_15[11],stage4_14[24]}
   );
   gpc615_5 gpc9841 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[24]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[8],stage4_16[9],stage4_15[12],stage4_14[25]}
   );
   gpc615_5 gpc9842 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[9],stage4_16[10],stage4_15[13]}
   );
   gpc615_5 gpc9843 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[37]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[7],stage4_17[10],stage4_16[11],stage4_15[14]}
   );
   gpc615_5 gpc9844 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[38]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[8],stage4_17[11],stage4_16[12],stage4_15[15]}
   );
   gpc615_5 gpc9845 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[39]},
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage4_19[3],stage4_18[9],stage4_17[12],stage4_16[13],stage4_15[16]}
   );
   gpc606_5 gpc9846 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[4],stage4_18[10],stage4_17[13]}
   );
   gpc606_5 gpc9847 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[5],stage4_18[11],stage4_17[14]}
   );
   gpc207_4 gpc9848 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[2],stage4_20[2],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc9849 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[3],stage4_20[3],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc9850 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[4],stage4_20[4],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc9851 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[5],stage4_20[5],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc9852 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[6],stage4_20[6],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc9853 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[7],stage4_20[7],stage4_19[11],stage4_18[17]}
   );
   gpc615_5 gpc9854 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46]},
      {stage3_19[12]},
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage4_22[0],stage4_21[8],stage4_20[8],stage4_19[12],stage4_18[18]}
   );
   gpc615_5 gpc9855 (
      {stage3_18[47], stage3_18[48], stage3_18[49], stage3_18[50], stage3_18[51]},
      {stage3_19[13]},
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage4_22[1],stage4_21[9],stage4_20[9],stage4_19[13],stage4_18[19]}
   );
   gpc606_5 gpc9856 (
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[2],stage4_21[10],stage4_20[10],stage4_19[14]}
   );
   gpc606_5 gpc9857 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[3],stage4_21[11],stage4_20[11],stage4_19[15]}
   );
   gpc615_5 gpc9858 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[24]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[4],stage4_21[12],stage4_20[12],stage4_19[16]}
   );
   gpc615_5 gpc9859 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35]},
      {stage3_20[25]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[5],stage4_21[13],stage4_20[13],stage4_19[17]}
   );
   gpc615_5 gpc9860 (
      {stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40]},
      {stage3_20[26]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[6],stage4_21[14],stage4_20[14],stage4_19[18]}
   );
   gpc615_5 gpc9861 (
      {stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45]},
      {stage3_20[27]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[7],stage4_21[15],stage4_20[15],stage4_19[19]}
   );
   gpc606_5 gpc9862 (
      {stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31], stage3_20[32], stage3_20[33]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[6],stage4_22[8],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc9863 (
      {stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37], stage3_20[38], stage3_20[39]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[7],stage4_22[9],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc9864 (
      {stage3_20[40], stage3_20[41], stage3_20[42], stage3_20[43], stage3_20[44], stage3_20[45]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[8],stage4_22[10],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc9865 (
      {stage3_20[46], stage3_20[47], stage3_20[48], stage3_20[49], stage3_20[50], stage3_20[51]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[9],stage4_22[11],stage4_21[19],stage4_20[19]}
   );
   gpc615_5 gpc9866 (
      {stage3_20[52], stage3_20[53], stage3_20[54], stage3_20[55], stage3_20[56]},
      {stage3_21[36]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[10],stage4_22[12],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc9867 (
      {stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[5],stage4_23[11],stage4_22[13],stage4_21[21]}
   );
   gpc606_5 gpc9868 (
      {stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[6],stage4_23[12],stage4_22[14],stage4_21[22]}
   );
   gpc606_5 gpc9869 (
      {stage3_21[49], stage3_21[50], stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[7],stage4_23[13],stage4_22[15],stage4_21[23]}
   );
   gpc606_5 gpc9870 (
      {stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59], stage3_21[60]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[8],stage4_23[14],stage4_22[16],stage4_21[24]}
   );
   gpc615_5 gpc9871 (
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[9],stage4_23[15],stage4_22[17]}
   );
   gpc615_5 gpc9872 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[10],stage4_23[16],stage4_22[18]}
   );
   gpc615_5 gpc9873 (
      {stage3_22[40], stage3_22[41], stage3_22[42], stage3_22[43], stage3_22[44]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[11],stage4_23[17],stage4_22[19]}
   );
   gpc615_5 gpc9874 (
      {stage3_22[45], stage3_22[46], stage3_22[47], stage3_22[48], stage3_22[49]},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[12],stage4_23[18],stage4_22[20]}
   );
   gpc615_5 gpc9875 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[13],stage4_23[19]}
   );
   gpc615_5 gpc9876 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[14],stage4_23[20]}
   );
   gpc615_5 gpc9877 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[15],stage4_23[21]}
   );
   gpc615_5 gpc9878 (
      {stage3_23[43], stage3_23[44], stage3_23[45], stage3_23[46], stage3_23[47]},
      {stage3_24[27]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[7],stage4_25[11],stage4_24[16],stage4_23[22]}
   );
   gpc615_5 gpc9879 (
      {stage3_23[48], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_24[28]},
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage4_27[4],stage4_26[8],stage4_25[12],stage4_24[17],stage4_23[23]}
   );
   gpc606_5 gpc9880 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[5],stage4_26[9],stage4_25[13]}
   );
   gpc606_5 gpc9881 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[6],stage4_26[10],stage4_25[14]}
   );
   gpc606_5 gpc9882 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46], stage3_25[47]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[7],stage4_26[11],stage4_25[15]}
   );
   gpc606_5 gpc9883 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[3],stage4_28[3],stage4_27[8],stage4_26[12]}
   );
   gpc606_5 gpc9884 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[4],stage4_28[4],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc9885 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[5],stage4_28[5],stage4_27[10],stage4_26[14]}
   );
   gpc606_5 gpc9886 (
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[6],stage4_28[6],stage4_27[11],stage4_26[15]}
   );
   gpc606_5 gpc9887 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage4_30[4],stage4_29[7],stage4_28[7],stage4_27[12],stage4_26[16]}
   );
   gpc606_5 gpc9888 (
      {stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage4_30[5],stage4_29[8],stage4_28[8],stage4_27[13],stage4_26[17]}
   );
   gpc606_5 gpc9889 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40], stage3_26[41]},
      {stage3_28[36], stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41]},
      {stage4_30[6],stage4_29[9],stage4_28[9],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc9890 (
      {stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47]},
      {stage3_28[42], stage3_28[43], stage3_28[44], stage3_28[45], stage3_28[46], stage3_28[47]},
      {stage4_30[7],stage4_29[10],stage4_28[10],stage4_27[15],stage4_26[19]}
   );
   gpc606_5 gpc9891 (
      {stage3_26[48], stage3_26[49], stage3_26[50], stage3_26[51], 1'b0, 1'b0},
      {stage3_28[48], stage3_28[49], stage3_28[50], stage3_28[51], stage3_28[52], stage3_28[53]},
      {stage4_30[8],stage4_29[11],stage4_28[11],stage4_27[16],stage4_26[20]}
   );
   gpc606_5 gpc9892 (
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[9],stage4_29[12],stage4_28[12],stage4_27[17]}
   );
   gpc606_5 gpc9893 (
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[10],stage4_29[13],stage4_28[13],stage4_27[18]}
   );
   gpc606_5 gpc9894 (
      {stage3_27[30], stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[11],stage4_29[14],stage4_28[14],stage4_27[19]}
   );
   gpc606_5 gpc9895 (
      {stage3_27[36], stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[12],stage4_29[15],stage4_28[15],stage4_27[20]}
   );
   gpc1163_5 gpc9896 (
      {stage3_29[24], stage3_29[25], stage3_29[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[4],stage4_30[13],stage4_29[16]}
   );
   gpc1163_5 gpc9897 (
      {stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[5],stage4_30[14],stage4_29[17]}
   );
   gpc1163_5 gpc9898 (
      {stage3_29[30], stage3_29[31], stage3_29[32]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[6],stage4_30[15],stage4_29[18]}
   );
   gpc1163_5 gpc9899 (
      {stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[7],stage4_30[16],stage4_29[19]}
   );
   gpc606_5 gpc9900 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[4],stage4_32[4],stage4_31[8],stage4_30[17],stage4_29[20]}
   );
   gpc606_5 gpc9901 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15]},
      {stage4_33[5],stage4_32[5],stage4_31[9],stage4_30[18],stage4_29[21]}
   );
   gpc606_5 gpc9902 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52], stage3_29[53]},
      {stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21]},
      {stage4_33[6],stage4_32[6],stage4_31[10],stage4_30[19],stage4_29[22]}
   );
   gpc606_5 gpc9903 (
      {stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57], stage3_29[58], 1'b0},
      {stage3_31[22], stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage4_33[7],stage4_32[7],stage4_31[11],stage4_30[20],stage4_29[23]}
   );
   gpc606_5 gpc9904 (
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_32[4], stage3_32[5], stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9]},
      {stage4_34[0],stage4_33[8],stage4_32[8],stage4_31[12],stage4_30[21]}
   );
   gpc606_5 gpc9905 (
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage4_34[1],stage4_33[9],stage4_32[9],stage4_31[13],stage4_30[22]}
   );
   gpc615_5 gpc9906 (
      {stage3_31[28], stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32]},
      {stage3_32[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[10],stage4_32[10],stage4_31[14]}
   );
   gpc615_5 gpc9907 (
      {stage3_31[33], stage3_31[34], stage3_31[35], stage3_31[36], stage3_31[37]},
      {stage3_32[17]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[11],stage4_32[11],stage4_31[15]}
   );
   gpc615_5 gpc9908 (
      {stage3_31[38], stage3_31[39], stage3_31[40], stage3_31[41], 1'b0},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[12],stage4_32[12],stage4_31[16]}
   );
   gpc2116_5 gpc9909 (
      {stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24]},
      {stage3_33[18]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[13],stage4_32[13]}
   );
   gpc2116_5 gpc9910 (
      {stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[19]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc9911 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[20]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc9912 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[21]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[16],stage4_32[16]}
   );
   gpc615_5 gpc9913 (
      {stage3_32[41], stage3_32[42], stage3_32[43], stage3_32[44], stage3_32[45]},
      {stage3_33[22]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[17],stage4_32[17]}
   );
   gpc615_5 gpc9914 (
      {stage3_32[46], stage3_32[47], stage3_32[48], stage3_32[49], stage3_32[50]},
      {stage3_33[23]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[8],stage4_34[10],stage4_33[18],stage4_32[18]}
   );
   gpc215_4 gpc9915 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28]},
      {stage3_34[26]},
      {stage3_35[4], stage3_35[5]},
      {stage4_36[6],stage4_35[9],stage4_34[11],stage4_33[19]}
   );
   gpc606_5 gpc9916 (
      {stage3_33[29], stage3_33[30], stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[7],stage4_35[10],stage4_34[12],stage4_33[20]}
   );
   gpc606_5 gpc9917 (
      {stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38], stage3_33[39], stage3_33[40]},
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage4_37[1],stage4_36[8],stage4_35[11],stage4_34[13],stage4_33[21]}
   );
   gpc606_5 gpc9918 (
      {stage3_33[41], stage3_33[42], stage3_33[43], stage3_33[44], stage3_33[45], stage3_33[46]},
      {stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage4_37[2],stage4_36[9],stage4_35[12],stage4_34[14],stage4_33[22]}
   );
   gpc606_5 gpc9919 (
      {stage3_33[47], stage3_33[48], stage3_33[49], stage3_33[50], stage3_33[51], stage3_33[52]},
      {stage3_35[24], stage3_35[25], stage3_35[26], stage3_35[27], stage3_35[28], stage3_35[29]},
      {stage4_37[3],stage4_36[10],stage4_35[13],stage4_34[15],stage4_33[23]}
   );
   gpc615_5 gpc9920 (
      {stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage3_35[30]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage4_38[0],stage4_37[4],stage4_36[11],stage4_35[14],stage4_34[16]}
   );
   gpc606_5 gpc9921 (
      {stage3_35[31], stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[1],stage4_37[5],stage4_36[12],stage4_35[15]}
   );
   gpc615_5 gpc9922 (
      {stage3_35[37], stage3_35[38], stage3_35[39], stage3_35[40], stage3_35[41]},
      {stage3_36[6]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[2],stage4_37[6],stage4_36[13],stage4_35[16]}
   );
   gpc615_5 gpc9923 (
      {stage3_35[42], stage3_35[43], stage3_35[44], stage3_35[45], stage3_35[46]},
      {stage3_36[7]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[3],stage4_37[7],stage4_36[14],stage4_35[17]}
   );
   gpc615_5 gpc9924 (
      {stage3_35[47], stage3_35[48], stage3_35[49], stage3_35[50], stage3_35[51]},
      {stage3_36[8]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[4],stage4_37[8],stage4_36[15],stage4_35[18]}
   );
   gpc606_5 gpc9925 (
      {stage3_36[9], stage3_36[10], stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[4],stage4_38[5],stage4_37[9],stage4_36[16]}
   );
   gpc606_5 gpc9926 (
      {stage3_36[15], stage3_36[16], stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[5],stage4_38[6],stage4_37[10],stage4_36[17]}
   );
   gpc606_5 gpc9927 (
      {stage3_36[21], stage3_36[22], stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[6],stage4_38[7],stage4_37[11],stage4_36[18]}
   );
   gpc606_5 gpc9928 (
      {stage3_36[27], stage3_36[28], stage3_36[29], stage3_36[30], stage3_36[31], stage3_36[32]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[7],stage4_38[8],stage4_37[12],stage4_36[19]}
   );
   gpc606_5 gpc9929 (
      {stage3_36[33], stage3_36[34], stage3_36[35], stage3_36[36], stage3_36[37], stage3_36[38]},
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28], stage3_38[29]},
      {stage4_40[4],stage4_39[8],stage4_38[9],stage4_37[13],stage4_36[20]}
   );
   gpc606_5 gpc9930 (
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[5],stage4_39[9],stage4_38[10],stage4_37[14]}
   );
   gpc606_5 gpc9931 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], 1'b0},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[6],stage4_39[10],stage4_38[11],stage4_37[15]}
   );
   gpc615_5 gpc9932 (
      {stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33], stage3_38[34]},
      {stage3_39[12]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[2],stage4_40[7],stage4_39[11],stage4_38[12]}
   );
   gpc615_5 gpc9933 (
      {stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38], stage3_38[39]},
      {stage3_39[13]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[3],stage4_40[8],stage4_39[12],stage4_38[13]}
   );
   gpc615_5 gpc9934 (
      {stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43], stage3_38[44]},
      {stage3_39[14]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[4],stage4_40[9],stage4_39[13],stage4_38[14]}
   );
   gpc615_5 gpc9935 (
      {stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48], stage3_38[49]},
      {stage3_39[15]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[5],stage4_40[10],stage4_39[14],stage4_38[15]}
   );
   gpc615_5 gpc9936 (
      {stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53], stage3_38[54]},
      {stage3_39[16]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[6],stage4_40[11],stage4_39[15],stage4_38[16]}
   );
   gpc615_5 gpc9937 (
      {stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58], stage3_38[59]},
      {stage3_39[17]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[7],stage4_40[12],stage4_39[16],stage4_38[17]}
   );
   gpc207_4 gpc9938 (
      {stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22], stage3_39[23], stage3_39[24]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[6],stage4_41[8],stage4_40[13],stage4_39[17]}
   );
   gpc207_4 gpc9939 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[7],stage4_41[9],stage4_40[14],stage4_39[18]}
   );
   gpc207_4 gpc9940 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[8],stage4_41[10],stage4_40[15],stage4_39[19]}
   );
   gpc207_4 gpc9941 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[9],stage4_41[11],stage4_40[16],stage4_39[20]}
   );
   gpc207_4 gpc9942 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[8], stage3_41[9]},
      {stage4_42[10],stage4_41[12],stage4_40[17],stage4_39[21]}
   );
   gpc207_4 gpc9943 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57], stage3_39[58], stage3_39[59]},
      {stage3_41[10], stage3_41[11]},
      {stage4_42[11],stage4_41[13],stage4_40[18],stage4_39[22]}
   );
   gpc606_5 gpc9944 (
      {stage3_41[12], stage3_41[13], stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[12],stage4_41[14]}
   );
   gpc606_5 gpc9945 (
      {stage3_41[18], stage3_41[19], stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[13],stage4_41[15]}
   );
   gpc606_5 gpc9946 (
      {stage3_41[24], stage3_41[25], stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[14],stage4_41[16]}
   );
   gpc606_5 gpc9947 (
      {stage3_41[30], stage3_41[31], stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[15],stage4_41[17]}
   );
   gpc606_5 gpc9948 (
      {stage3_41[36], stage3_41[37], stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41]},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[16],stage4_41[18]}
   );
   gpc606_5 gpc9949 (
      {stage3_41[42], stage3_41[43], stage3_41[44], stage3_41[45], stage3_41[46], stage3_41[47]},
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[17],stage4_41[19]}
   );
   gpc606_5 gpc9950 (
      {stage3_41[48], stage3_41[49], stage3_41[50], stage3_41[51], stage3_41[52], stage3_41[53]},
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage4_45[6],stage4_44[6],stage4_43[6],stage4_42[18],stage4_41[20]}
   );
   gpc207_4 gpc9951 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[7],stage4_44[7],stage4_43[7],stage4_42[19]}
   );
   gpc207_4 gpc9952 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[8],stage4_44[8],stage4_43[8],stage4_42[20]}
   );
   gpc615_5 gpc9953 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18]},
      {stage3_43[42]},
      {stage3_44[4], stage3_44[5], stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[9],stage4_42[21]}
   );
   gpc615_5 gpc9954 (
      {stage3_42[19], stage3_42[20], stage3_42[21], stage3_42[22], stage3_42[23]},
      {stage3_43[43]},
      {stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[10],stage4_42[22]}
   );
   gpc615_5 gpc9955 (
      {stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27], stage3_42[28]},
      {stage3_43[44]},
      {stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21]},
      {stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[11],stage4_42[23]}
   );
   gpc615_5 gpc9956 (
      {stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_43[45]},
      {stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26], stage3_44[27]},
      {stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[12],stage4_42[24]}
   );
   gpc615_5 gpc9957 (
      {stage3_42[34], stage3_42[35], stage3_42[36], stage3_42[37], stage3_42[38]},
      {stage3_43[46]},
      {stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31], stage3_44[32], stage3_44[33]},
      {stage4_46[4],stage4_45[13],stage4_44[13],stage4_43[13],stage4_42[25]}
   );
   gpc615_5 gpc9958 (
      {stage3_42[39], stage3_42[40], stage3_42[41], stage3_42[42], stage3_42[43]},
      {stage3_43[47]},
      {stage3_44[34], stage3_44[35], stage3_44[36], stage3_44[37], stage3_44[38], stage3_44[39]},
      {stage4_46[5],stage4_45[14],stage4_44[14],stage4_43[14],stage4_42[26]}
   );
   gpc615_5 gpc9959 (
      {stage3_42[44], stage3_42[45], stage3_42[46], stage3_42[47], stage3_42[48]},
      {stage3_43[48]},
      {stage3_44[40], stage3_44[41], stage3_44[42], stage3_44[43], stage3_44[44], stage3_44[45]},
      {stage4_46[6],stage4_45[15],stage4_44[15],stage4_43[15],stage4_42[27]}
   );
   gpc615_5 gpc9960 (
      {stage3_42[49], stage3_42[50], stage3_42[51], stage3_42[52], stage3_42[53]},
      {stage3_43[49]},
      {stage3_44[46], stage3_44[47], stage3_44[48], stage3_44[49], stage3_44[50], stage3_44[51]},
      {stage4_46[7],stage4_45[16],stage4_44[16],stage4_43[16],stage4_42[28]}
   );
   gpc615_5 gpc9961 (
      {stage3_43[50], stage3_43[51], stage3_43[52], stage3_43[53], stage3_43[54]},
      {stage3_44[52]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[8],stage4_45[17],stage4_44[17],stage4_43[17]}
   );
   gpc1343_5 gpc9962 (
      {stage3_44[53], stage3_44[54], stage3_44[55]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[1],stage4_46[9],stage4_45[18],stage4_44[18]}
   );
   gpc1343_5 gpc9963 (
      {stage3_44[56], stage3_44[57], stage3_44[58]},
      {stage3_45[10], stage3_45[11], stage3_45[12], stage3_45[13]},
      {stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[1]},
      {stage4_48[1],stage4_47[2],stage4_46[10],stage4_45[19],stage4_44[19]}
   );
   gpc1343_5 gpc9964 (
      {stage3_44[59], stage3_44[60], stage3_44[61]},
      {stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_46[6], stage3_46[7], stage3_46[8]},
      {stage3_47[2]},
      {stage4_48[2],stage4_47[3],stage4_46[11],stage4_45[20],stage4_44[20]}
   );
   gpc623_5 gpc9965 (
      {stage3_44[62], stage3_44[63], stage3_44[64]},
      {stage3_45[18], stage3_45[19]},
      {stage3_46[9], stage3_46[10], stage3_46[11], stage3_46[12], stage3_46[13], stage3_46[14]},
      {stage4_48[3],stage4_47[4],stage4_46[12],stage4_45[21],stage4_44[21]}
   );
   gpc623_5 gpc9966 (
      {stage3_44[65], stage3_44[66], stage3_44[67]},
      {stage3_45[20], stage3_45[21]},
      {stage3_46[15], stage3_46[16], stage3_46[17], stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage4_48[4],stage4_47[5],stage4_46[13],stage4_45[22],stage4_44[22]}
   );
   gpc606_5 gpc9967 (
      {stage3_45[22], stage3_45[23], stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27]},
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8]},
      {stage4_49[0],stage4_48[5],stage4_47[6],stage4_46[14],stage4_45[23]}
   );
   gpc606_5 gpc9968 (
      {stage3_45[28], stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage4_49[1],stage4_48[6],stage4_47[7],stage4_46[15],stage4_45[24]}
   );
   gpc606_5 gpc9969 (
      {stage3_45[34], stage3_45[35], stage3_45[36], stage3_45[37], stage3_45[38], stage3_45[39]},
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage4_49[2],stage4_48[7],stage4_47[8],stage4_46[16],stage4_45[25]}
   );
   gpc615_5 gpc9970 (
      {stage3_46[21], stage3_46[22], stage3_46[23], stage3_46[24], stage3_46[25]},
      {stage3_47[21]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[3],stage4_48[8],stage4_47[9],stage4_46[17]}
   );
   gpc615_5 gpc9971 (
      {stage3_46[26], stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30]},
      {stage3_47[22]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[4],stage4_48[9],stage4_47[10],stage4_46[18]}
   );
   gpc615_5 gpc9972 (
      {stage3_46[31], stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35]},
      {stage3_47[23]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[5],stage4_48[10],stage4_47[11],stage4_46[19]}
   );
   gpc615_5 gpc9973 (
      {stage3_46[36], stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40]},
      {stage3_47[24]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[6],stage4_48[11],stage4_47[12],stage4_46[20]}
   );
   gpc615_5 gpc9974 (
      {stage3_46[41], stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45]},
      {stage3_47[25]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[7],stage4_48[12],stage4_47[13],stage4_46[21]}
   );
   gpc615_5 gpc9975 (
      {stage3_47[26], stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30]},
      {stage3_48[30]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[5],stage4_49[8],stage4_48[13],stage4_47[14]}
   );
   gpc615_5 gpc9976 (
      {stage3_47[31], stage3_47[32], stage3_47[33], stage3_47[34], stage3_47[35]},
      {stage3_48[31]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[6],stage4_49[9],stage4_48[14],stage4_47[15]}
   );
   gpc615_5 gpc9977 (
      {stage3_47[36], stage3_47[37], stage3_47[38], stage3_47[39], stage3_47[40]},
      {stage3_48[32]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[7],stage4_49[10],stage4_48[15],stage4_47[16]}
   );
   gpc615_5 gpc9978 (
      {stage3_47[41], stage3_47[42], stage3_47[43], stage3_47[44], stage3_47[45]},
      {stage3_48[33]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[8],stage4_49[11],stage4_48[16],stage4_47[17]}
   );
   gpc615_5 gpc9979 (
      {stage3_47[46], stage3_47[47], stage3_47[48], stage3_47[49], stage3_47[50]},
      {stage3_48[34]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[9],stage4_49[12],stage4_48[17],stage4_47[18]}
   );
   gpc615_5 gpc9980 (
      {stage3_47[51], stage3_47[52], stage3_47[53], stage3_47[54], stage3_47[55]},
      {stage3_48[35]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[10],stage4_49[13],stage4_48[18],stage4_47[19]}
   );
   gpc615_5 gpc9981 (
      {stage3_47[56], stage3_47[57], stage3_47[58], stage3_47[59], stage3_47[60]},
      {stage3_48[36]},
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage4_51[6],stage4_50[11],stage4_49[14],stage4_48[19],stage4_47[20]}
   );
   gpc615_5 gpc9982 (
      {stage3_47[61], stage3_47[62], stage3_47[63], stage3_47[64], stage3_47[65]},
      {1'b0},
      {stage3_49[42], stage3_49[43], stage3_49[44], stage3_49[45], stage3_49[46], stage3_49[47]},
      {stage4_51[7],stage4_50[12],stage4_49[15],stage4_48[20],stage4_47[21]}
   );
   gpc615_5 gpc9983 (
      {stage3_47[66], stage3_47[67], stage3_47[68], stage3_47[69], stage3_47[70]},
      {1'b0},
      {stage3_49[48], stage3_49[49], stage3_49[50], stage3_49[51], stage3_49[52], stage3_49[53]},
      {stage4_51[8],stage4_50[13],stage4_49[16],stage4_48[21],stage4_47[22]}
   );
   gpc117_4 gpc9984 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[0]},
      {stage3_52[0]},
      {stage4_53[0],stage4_52[0],stage4_51[9],stage4_50[14]}
   );
   gpc117_4 gpc9985 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[1]},
      {stage3_52[1]},
      {stage4_53[1],stage4_52[1],stage4_51[10],stage4_50[15]}
   );
   gpc117_4 gpc9986 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18], stage3_50[19], stage3_50[20]},
      {stage3_51[2]},
      {stage3_52[2]},
      {stage4_53[2],stage4_52[2],stage4_51[11],stage4_50[16]}
   );
   gpc117_4 gpc9987 (
      {stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27]},
      {stage3_51[3]},
      {stage3_52[3]},
      {stage4_53[3],stage4_52[3],stage4_51[12],stage4_50[17]}
   );
   gpc117_4 gpc9988 (
      {stage3_50[28], stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33], stage3_50[34]},
      {stage3_51[4]},
      {stage3_52[4]},
      {stage4_53[4],stage4_52[4],stage4_51[13],stage4_50[18]}
   );
   gpc117_4 gpc9989 (
      {stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38], stage3_50[39], stage3_50[40], stage3_50[41]},
      {stage3_51[5]},
      {stage3_52[5]},
      {stage4_53[5],stage4_52[5],stage4_51[14],stage4_50[19]}
   );
   gpc117_4 gpc9990 (
      {stage3_50[42], stage3_50[43], stage3_50[44], stage3_50[45], stage3_50[46], stage3_50[47], stage3_50[48]},
      {stage3_51[6]},
      {stage3_52[6]},
      {stage4_53[6],stage4_52[6],stage4_51[15],stage4_50[20]}
   );
   gpc117_4 gpc9991 (
      {stage3_50[49], stage3_50[50], stage3_50[51], stage3_50[52], stage3_50[53], stage3_50[54], stage3_50[55]},
      {stage3_51[7]},
      {stage3_52[7]},
      {stage4_53[7],stage4_52[7],stage4_51[16],stage4_50[21]}
   );
   gpc117_4 gpc9992 (
      {stage3_50[56], stage3_50[57], stage3_50[58], stage3_50[59], stage3_50[60], stage3_50[61], stage3_50[62]},
      {stage3_51[8]},
      {stage3_52[8]},
      {stage4_53[8],stage4_52[8],stage4_51[17],stage4_50[22]}
   );
   gpc2135_5 gpc9993 (
      {stage3_51[9], stage3_51[10], stage3_51[11], stage3_51[12], stage3_51[13]},
      {stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[0],stage4_53[9],stage4_52[9],stage4_51[18]}
   );
   gpc2135_5 gpc9994 (
      {stage3_51[14], stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18]},
      {stage3_52[12], stage3_52[13], stage3_52[14]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[1],stage4_53[10],stage4_52[10],stage4_51[19]}
   );
   gpc2135_5 gpc9995 (
      {stage3_51[19], stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23]},
      {stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[2],stage4_53[11],stage4_52[11],stage4_51[20]}
   );
   gpc2135_5 gpc9996 (
      {stage3_51[24], stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28]},
      {stage3_52[18], stage3_52[19], stage3_52[20]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[3],stage4_53[12],stage4_52[12],stage4_51[21]}
   );
   gpc2135_5 gpc9997 (
      {stage3_51[29], stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33]},
      {stage3_52[21], stage3_52[22], stage3_52[23]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[4],stage4_53[13],stage4_52[13],stage4_51[22]}
   );
   gpc2135_5 gpc9998 (
      {stage3_51[34], stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38]},
      {stage3_52[24], stage3_52[25], stage3_52[26]},
      {stage3_53[5]},
      {stage3_54[10], stage3_54[11]},
      {stage4_55[5],stage4_54[5],stage4_53[14],stage4_52[14],stage4_51[23]}
   );
   gpc2135_5 gpc9999 (
      {stage3_51[39], stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43]},
      {stage3_52[27], stage3_52[28], stage3_52[29]},
      {stage3_53[6]},
      {stage3_54[12], stage3_54[13]},
      {stage4_55[6],stage4_54[6],stage4_53[15],stage4_52[15],stage4_51[24]}
   );
   gpc2135_5 gpc10000 (
      {stage3_51[44], stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48]},
      {stage3_52[30], stage3_52[31], stage3_52[32]},
      {stage3_53[7]},
      {stage3_54[14], stage3_54[15]},
      {stage4_55[7],stage4_54[7],stage4_53[16],stage4_52[16],stage4_51[25]}
   );
   gpc2135_5 gpc10001 (
      {stage3_51[49], stage3_51[50], stage3_51[51], stage3_51[52], stage3_51[53]},
      {stage3_52[33], stage3_52[34], stage3_52[35]},
      {stage3_53[8]},
      {stage3_54[16], stage3_54[17]},
      {stage4_55[8],stage4_54[8],stage4_53[17],stage4_52[17],stage4_51[26]}
   );
   gpc606_5 gpc10002 (
      {stage3_52[36], stage3_52[37], stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41]},
      {stage3_54[18], stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage4_56[0],stage4_55[9],stage4_54[9],stage4_53[18],stage4_52[18]}
   );
   gpc606_5 gpc10003 (
      {stage3_52[42], stage3_52[43], stage3_52[44], stage3_52[45], stage3_52[46], stage3_52[47]},
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28], stage3_54[29]},
      {stage4_56[1],stage4_55[10],stage4_54[10],stage4_53[19],stage4_52[19]}
   );
   gpc606_5 gpc10004 (
      {stage3_52[48], stage3_52[49], stage3_52[50], stage3_52[51], stage3_52[52], stage3_52[53]},
      {stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33], stage3_54[34], stage3_54[35]},
      {stage4_56[2],stage4_55[11],stage4_54[11],stage4_53[20],stage4_52[20]}
   );
   gpc1415_5 gpc10005 (
      {stage3_53[9], stage3_53[10], stage3_53[11], stage3_53[12], stage3_53[13]},
      {stage3_54[36]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[3],stage4_55[12],stage4_54[12],stage4_53[21]}
   );
   gpc1415_5 gpc10006 (
      {stage3_53[14], stage3_53[15], stage3_53[16], stage3_53[17], stage3_53[18]},
      {stage3_54[37]},
      {stage3_55[4], stage3_55[5], stage3_55[6], stage3_55[7]},
      {stage3_56[1]},
      {stage4_57[1],stage4_56[4],stage4_55[13],stage4_54[13],stage4_53[22]}
   );
   gpc1415_5 gpc10007 (
      {stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22], stage3_53[23]},
      {stage3_54[38]},
      {stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage3_56[2]},
      {stage4_57[2],stage4_56[5],stage4_55[14],stage4_54[14],stage4_53[23]}
   );
   gpc1415_5 gpc10008 (
      {stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_54[39]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15]},
      {stage3_56[3]},
      {stage4_57[3],stage4_56[6],stage4_55[15],stage4_54[15],stage4_53[24]}
   );
   gpc606_5 gpc10009 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[16], stage3_55[17], stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21]},
      {stage4_57[4],stage4_56[7],stage4_55[16],stage4_54[16],stage4_53[25]}
   );
   gpc606_5 gpc10010 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39], stage3_53[40]},
      {stage3_55[22], stage3_55[23], stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27]},
      {stage4_57[5],stage4_56[8],stage4_55[17],stage4_54[17],stage4_53[26]}
   );
   gpc606_5 gpc10011 (
      {stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44], stage3_53[45], stage3_53[46]},
      {stage3_55[28], stage3_55[29], stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33]},
      {stage4_57[6],stage4_56[9],stage4_55[18],stage4_54[18],stage4_53[27]}
   );
   gpc606_5 gpc10012 (
      {stage3_53[47], stage3_53[48], stage3_53[49], stage3_53[50], stage3_53[51], stage3_53[52]},
      {stage3_55[34], stage3_55[35], stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39]},
      {stage4_57[7],stage4_56[10],stage4_55[19],stage4_54[19],stage4_53[28]}
   );
   gpc207_4 gpc10013 (
      {stage3_54[40], stage3_54[41], stage3_54[42], stage3_54[43], stage3_54[44], stage3_54[45], stage3_54[46]},
      {stage3_56[4], stage3_56[5]},
      {stage4_57[8],stage4_56[11],stage4_55[20],stage4_54[20]}
   );
   gpc207_4 gpc10014 (
      {stage3_54[47], stage3_54[48], stage3_54[49], stage3_54[50], stage3_54[51], stage3_54[52], stage3_54[53]},
      {stage3_56[6], stage3_56[7]},
      {stage4_57[9],stage4_56[12],stage4_55[21],stage4_54[21]}
   );
   gpc606_5 gpc10015 (
      {stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12], stage3_56[13]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[0],stage4_58[0],stage4_57[10],stage4_56[13]}
   );
   gpc606_5 gpc10016 (
      {stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18], stage3_56[19]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[1],stage4_58[1],stage4_57[11],stage4_56[14]}
   );
   gpc606_5 gpc10017 (
      {stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23], stage3_56[24], stage3_56[25]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[2],stage4_58[2],stage4_57[12],stage4_56[15]}
   );
   gpc1163_5 gpc10018 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[3],stage4_59[3],stage4_58[3],stage4_57[13]}
   );
   gpc1163_5 gpc10019 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[4],stage4_59[4],stage4_58[4],stage4_57[14]}
   );
   gpc1163_5 gpc10020 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[5],stage4_59[5],stage4_58[5],stage4_57[15]}
   );
   gpc606_5 gpc10021 (
      {stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7], stage3_59[8]},
      {stage4_61[3],stage4_60[6],stage4_59[6],stage4_58[6],stage4_57[16]}
   );
   gpc606_5 gpc10022 (
      {stage3_57[15], stage3_57[16], stage3_57[17], stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[4],stage4_60[7],stage4_59[7],stage4_58[7],stage4_57[17]}
   );
   gpc606_5 gpc10023 (
      {stage3_57[21], stage3_57[22], stage3_57[23], stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[5],stage4_60[8],stage4_59[8],stage4_58[8],stage4_57[18]}
   );
   gpc606_5 gpc10024 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[6],stage4_60[9],stage4_59[9],stage4_58[9],stage4_57[19]}
   );
   gpc606_5 gpc10025 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[7],stage4_60[10],stage4_59[10],stage4_58[10],stage4_57[20]}
   );
   gpc606_5 gpc10026 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43], stage3_57[44]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[8],stage4_60[11],stage4_59[11],stage4_58[11],stage4_57[21]}
   );
   gpc606_5 gpc10027 (
      {stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48], stage3_57[49], stage3_57[50]},
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43], stage3_59[44]},
      {stage4_61[9],stage4_60[12],stage4_59[12],stage4_58[12],stage4_57[22]}
   );
   gpc1406_5 gpc10028 (
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_60[3], stage3_60[4], stage3_60[5], stage3_60[6]},
      {stage3_61[0]},
      {stage4_62[0],stage4_61[10],stage4_60[13],stage4_59[13],stage4_58[13]}
   );
   gpc606_5 gpc10029 (
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10], stage3_60[11], stage3_60[12]},
      {stage4_62[1],stage4_61[11],stage4_60[14],stage4_59[14],stage4_58[14]}
   );
   gpc1406_5 gpc10030 (
      {stage3_60[13], stage3_60[14], stage3_60[15], stage3_60[16], stage3_60[17], stage3_60[18]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0]},
      {stage4_64[0],stage4_63[0],stage4_62[2],stage4_61[12],stage4_60[15]}
   );
   gpc606_5 gpc10031 (
      {stage3_60[19], stage3_60[20], stage3_60[21], stage3_60[22], stage3_60[23], stage3_60[24]},
      {stage3_62[4], stage3_62[5], stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9]},
      {stage4_64[1],stage4_63[1],stage4_62[3],stage4_61[13],stage4_60[16]}
   );
   gpc606_5 gpc10032 (
      {stage3_60[25], stage3_60[26], stage3_60[27], stage3_60[28], stage3_60[29], stage3_60[30]},
      {stage3_62[10], stage3_62[11], stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15]},
      {stage4_64[2],stage4_63[2],stage4_62[4],stage4_61[14],stage4_60[17]}
   );
   gpc606_5 gpc10033 (
      {stage3_60[31], stage3_60[32], stage3_60[33], stage3_60[34], stage3_60[35], stage3_60[36]},
      {stage3_62[16], stage3_62[17], stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21]},
      {stage4_64[3],stage4_63[3],stage4_62[5],stage4_61[15],stage4_60[18]}
   );
   gpc606_5 gpc10034 (
      {stage3_60[37], stage3_60[38], stage3_60[39], stage3_60[40], stage3_60[41], stage3_60[42]},
      {stage3_62[22], stage3_62[23], stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27]},
      {stage4_64[4],stage4_63[4],stage4_62[6],stage4_61[16],stage4_60[19]}
   );
   gpc606_5 gpc10035 (
      {stage3_60[43], stage3_60[44], stage3_60[45], stage3_60[46], stage3_60[47], stage3_60[48]},
      {stage3_62[28], stage3_62[29], stage3_62[30], stage3_62[31], stage3_62[32], stage3_62[33]},
      {stage4_64[5],stage4_63[5],stage4_62[7],stage4_61[17],stage4_60[20]}
   );
   gpc606_5 gpc10036 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5], stage3_61[6]},
      {stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6]},
      {stage4_65[0],stage4_64[6],stage4_63[6],stage4_62[8],stage4_61[18]}
   );
   gpc606_5 gpc10037 (
      {stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11], stage3_61[12]},
      {stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11], stage3_63[12]},
      {stage4_65[1],stage4_64[7],stage4_63[7],stage4_62[9],stage4_61[19]}
   );
   gpc606_5 gpc10038 (
      {stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17], stage3_61[18]},
      {stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17], stage3_63[18]},
      {stage4_65[2],stage4_64[8],stage4_63[8],stage4_62[10],stage4_61[20]}
   );
   gpc606_5 gpc10039 (
      {stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23], stage3_61[24]},
      {stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23], stage3_63[24]},
      {stage4_65[3],stage4_64[9],stage4_63[9],stage4_62[11],stage4_61[21]}
   );
   gpc606_5 gpc10040 (
      {stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29], stage3_61[30]},
      {stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29], stage3_63[30]},
      {stage4_65[4],stage4_64[10],stage4_63[10],stage4_62[12],stage4_61[22]}
   );
   gpc606_5 gpc10041 (
      {stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35], stage3_61[36]},
      {stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35], stage3_63[36]},
      {stage4_65[5],stage4_64[11],stage4_63[11],stage4_62[13],stage4_61[23]}
   );
   gpc606_5 gpc10042 (
      {stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41], stage3_61[42]},
      {stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41], stage3_63[42]},
      {stage4_65[6],stage4_64[12],stage4_63[12],stage4_62[14],stage4_61[24]}
   );
   gpc606_5 gpc10043 (
      {stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47], stage3_61[48]},
      {stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47], stage3_63[48]},
      {stage4_65[7],stage4_64[13],stage4_63[13],stage4_62[15],stage4_61[25]}
   );
   gpc606_5 gpc10044 (
      {stage3_61[49], stage3_61[50], stage3_61[51], stage3_61[52], stage3_61[53], stage3_61[54]},
      {stage3_63[49], stage3_63[50], stage3_63[51], stage3_63[52], stage3_63[53], stage3_63[54]},
      {stage4_65[8],stage4_64[14],stage4_63[14],stage4_62[16],stage4_61[26]}
   );
   gpc606_5 gpc10045 (
      {stage3_63[55], stage3_63[56], stage3_63[57], stage3_63[58], stage3_63[59], stage3_63[60]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[9],stage4_64[15],stage4_63[15]}
   );
   gpc606_5 gpc10046 (
      {stage3_63[61], stage3_63[62], stage3_63[63], stage3_63[64], stage3_63[65], stage3_63[66]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[1],stage4_65[10],stage4_64[16],stage4_63[16]}
   );
   gpc606_5 gpc10047 (
      {stage3_63[67], stage3_63[68], stage3_63[69], stage3_63[70], stage3_63[71], 1'b0},
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage4_67[2],stage4_66[2],stage4_65[11],stage4_64[17],stage4_63[17]}
   );
   gpc1163_5 gpc10048 (
      {stage3_64[0], stage3_64[1], stage3_64[2]},
      {stage3_65[18], stage3_65[19], stage3_65[20], stage3_65[21], stage3_65[22], stage3_65[23]},
      {stage3_66[0]},
      {stage3_67[0]},
      {stage4_68[0],stage4_67[3],stage4_66[3],stage4_65[12],stage4_64[18]}
   );
   gpc606_5 gpc10049 (
      {stage3_64[3], stage3_64[4], stage3_64[5], stage3_64[6], stage3_64[7], stage3_64[8]},
      {stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5], stage3_66[6]},
      {stage4_68[1],stage4_67[4],stage4_66[4],stage4_65[13],stage4_64[19]}
   );
   gpc606_5 gpc10050 (
      {stage3_64[9], stage3_64[10], stage3_64[11], stage3_64[12], stage3_64[13], stage3_64[14]},
      {stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11], stage3_66[12]},
      {stage4_68[2],stage4_67[5],stage4_66[5],stage4_65[14],stage4_64[20]}
   );
   gpc606_5 gpc10051 (
      {stage3_64[15], stage3_64[16], stage3_64[17], stage3_64[18], stage3_64[19], stage3_64[20]},
      {stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17], stage3_66[18]},
      {stage4_68[3],stage4_67[6],stage4_66[6],stage4_65[15],stage4_64[21]}
   );
   gpc606_5 gpc10052 (
      {stage3_64[21], stage3_64[22], stage3_64[23], stage3_64[24], stage3_64[25], stage3_64[26]},
      {stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23], stage3_66[24]},
      {stage4_68[4],stage4_67[7],stage4_66[7],stage4_65[16],stage4_64[22]}
   );
   gpc606_5 gpc10053 (
      {stage3_64[27], stage3_64[28], stage3_64[29], stage3_64[30], stage3_64[31], stage3_64[32]},
      {stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29], stage3_66[30]},
      {stage4_68[5],stage4_67[8],stage4_66[8],stage4_65[17],stage4_64[23]}
   );
   gpc606_5 gpc10054 (
      {stage3_64[33], stage3_64[34], stage3_64[35], stage3_64[36], stage3_64[37], stage3_64[38]},
      {stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35], stage3_66[36]},
      {stage4_68[6],stage4_67[9],stage4_66[9],stage4_65[18],stage4_64[24]}
   );
   gpc606_5 gpc10055 (
      {stage3_64[39], stage3_64[40], stage3_64[41], stage3_64[42], stage3_64[43], stage3_64[44]},
      {stage3_66[37], stage3_66[38], stage3_66[39], stage3_66[40], stage3_66[41], stage3_66[42]},
      {stage4_68[7],stage4_67[10],stage4_66[10],stage4_65[19],stage4_64[25]}
   );
   gpc606_5 gpc10056 (
      {stage3_64[45], stage3_64[46], stage3_64[47], stage3_64[48], stage3_64[49], stage3_64[50]},
      {stage3_66[43], stage3_66[44], stage3_66[45], stage3_66[46], stage3_66[47], stage3_66[48]},
      {stage4_68[8],stage4_67[11],stage4_66[11],stage4_65[20],stage4_64[26]}
   );
   gpc606_5 gpc10057 (
      {stage3_65[24], stage3_65[25], stage3_65[26], stage3_65[27], stage3_65[28], stage3_65[29]},
      {stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5], stage3_67[6]},
      {stage4_69[0],stage4_68[9],stage4_67[12],stage4_66[12],stage4_65[21]}
   );
   gpc606_5 gpc10058 (
      {stage3_65[30], stage3_65[31], stage3_65[32], 1'b0, 1'b0, 1'b0},
      {stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11], stage3_67[12]},
      {stage4_69[1],stage4_68[10],stage4_67[13],stage4_66[13],stage4_65[22]}
   );
   gpc606_5 gpc10059 (
      {stage3_66[49], stage3_66[50], stage3_66[51], stage3_66[52], stage3_66[53], 1'b0},
      {stage3_68[0], stage3_68[1], stage3_68[2], stage3_68[3], stage3_68[4], 1'b0},
      {stage4_70[0],stage4_69[2],stage4_68[11],stage4_67[14],stage4_66[14]}
   );
   gpc1_1 gpc10060 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc10061 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc10062 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc10063 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc10064 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc10065 (
      {stage3_1[24]},
      {stage4_1[5]}
   );
   gpc1_1 gpc10066 (
      {stage3_1[25]},
      {stage4_1[6]}
   );
   gpc1_1 gpc10067 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc10068 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc10069 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc10070 (
      {stage3_3[39]},
      {stage4_3[9]}
   );
   gpc1_1 gpc10071 (
      {stage3_3[40]},
      {stage4_3[10]}
   );
   gpc1_1 gpc10072 (
      {stage3_3[41]},
      {stage4_3[11]}
   );
   gpc1_1 gpc10073 (
      {stage3_3[42]},
      {stage4_3[12]}
   );
   gpc1_1 gpc10074 (
      {stage3_3[43]},
      {stage4_3[13]}
   );
   gpc1_1 gpc10075 (
      {stage3_3[44]},
      {stage4_3[14]}
   );
   gpc1_1 gpc10076 (
      {stage3_3[45]},
      {stage4_3[15]}
   );
   gpc1_1 gpc10077 (
      {stage3_3[46]},
      {stage4_3[16]}
   );
   gpc1_1 gpc10078 (
      {stage3_3[47]},
      {stage4_3[17]}
   );
   gpc1_1 gpc10079 (
      {stage3_3[48]},
      {stage4_3[18]}
   );
   gpc1_1 gpc10080 (
      {stage3_3[49]},
      {stage4_3[19]}
   );
   gpc1_1 gpc10081 (
      {stage3_3[50]},
      {stage4_3[20]}
   );
   gpc1_1 gpc10082 (
      {stage3_3[51]},
      {stage4_3[21]}
   );
   gpc1_1 gpc10083 (
      {stage3_4[51]},
      {stage4_4[16]}
   );
   gpc1_1 gpc10084 (
      {stage3_4[52]},
      {stage4_4[17]}
   );
   gpc1_1 gpc10085 (
      {stage3_4[53]},
      {stage4_4[18]}
   );
   gpc1_1 gpc10086 (
      {stage3_4[54]},
      {stage4_4[19]}
   );
   gpc1_1 gpc10087 (
      {stage3_4[55]},
      {stage4_4[20]}
   );
   gpc1_1 gpc10088 (
      {stage3_4[56]},
      {stage4_4[21]}
   );
   gpc1_1 gpc10089 (
      {stage3_4[57]},
      {stage4_4[22]}
   );
   gpc1_1 gpc10090 (
      {stage3_4[58]},
      {stage4_4[23]}
   );
   gpc1_1 gpc10091 (
      {stage3_4[59]},
      {stage4_4[24]}
   );
   gpc1_1 gpc10092 (
      {stage3_5[24]},
      {stage4_5[16]}
   );
   gpc1_1 gpc10093 (
      {stage3_5[25]},
      {stage4_5[17]}
   );
   gpc1_1 gpc10094 (
      {stage3_5[26]},
      {stage4_5[18]}
   );
   gpc1_1 gpc10095 (
      {stage3_5[27]},
      {stage4_5[19]}
   );
   gpc1_1 gpc10096 (
      {stage3_5[28]},
      {stage4_5[20]}
   );
   gpc1_1 gpc10097 (
      {stage3_5[29]},
      {stage4_5[21]}
   );
   gpc1_1 gpc10098 (
      {stage3_5[30]},
      {stage4_5[22]}
   );
   gpc1_1 gpc10099 (
      {stage3_5[31]},
      {stage4_5[23]}
   );
   gpc1_1 gpc10100 (
      {stage3_5[32]},
      {stage4_5[24]}
   );
   gpc1_1 gpc10101 (
      {stage3_5[33]},
      {stage4_5[25]}
   );
   gpc1_1 gpc10102 (
      {stage3_5[34]},
      {stage4_5[26]}
   );
   gpc1_1 gpc10103 (
      {stage3_5[35]},
      {stage4_5[27]}
   );
   gpc1_1 gpc10104 (
      {stage3_5[36]},
      {stage4_5[28]}
   );
   gpc1_1 gpc10105 (
      {stage3_5[37]},
      {stage4_5[29]}
   );
   gpc1_1 gpc10106 (
      {stage3_5[38]},
      {stage4_5[30]}
   );
   gpc1_1 gpc10107 (
      {stage3_5[39]},
      {stage4_5[31]}
   );
   gpc1_1 gpc10108 (
      {stage3_5[40]},
      {stage4_5[32]}
   );
   gpc1_1 gpc10109 (
      {stage3_5[41]},
      {stage4_5[33]}
   );
   gpc1_1 gpc10110 (
      {stage3_5[42]},
      {stage4_5[34]}
   );
   gpc1_1 gpc10111 (
      {stage3_5[43]},
      {stage4_5[35]}
   );
   gpc1_1 gpc10112 (
      {stage3_5[44]},
      {stage4_5[36]}
   );
   gpc1_1 gpc10113 (
      {stage3_5[45]},
      {stage4_5[37]}
   );
   gpc1_1 gpc10114 (
      {stage3_5[46]},
      {stage4_5[38]}
   );
   gpc1_1 gpc10115 (
      {stage3_5[47]},
      {stage4_5[39]}
   );
   gpc1_1 gpc10116 (
      {stage3_5[48]},
      {stage4_5[40]}
   );
   gpc1_1 gpc10117 (
      {stage3_5[49]},
      {stage4_5[41]}
   );
   gpc1_1 gpc10118 (
      {stage3_5[50]},
      {stage4_5[42]}
   );
   gpc1_1 gpc10119 (
      {stage3_5[51]},
      {stage4_5[43]}
   );
   gpc1_1 gpc10120 (
      {stage3_5[52]},
      {stage4_5[44]}
   );
   gpc1_1 gpc10121 (
      {stage3_5[53]},
      {stage4_5[45]}
   );
   gpc1_1 gpc10122 (
      {stage3_5[54]},
      {stage4_5[46]}
   );
   gpc1_1 gpc10123 (
      {stage3_6[62]},
      {stage4_6[16]}
   );
   gpc1_1 gpc10124 (
      {stage3_6[63]},
      {stage4_6[17]}
   );
   gpc1_1 gpc10125 (
      {stage3_6[64]},
      {stage4_6[18]}
   );
   gpc1_1 gpc10126 (
      {stage3_6[65]},
      {stage4_6[19]}
   );
   gpc1_1 gpc10127 (
      {stage3_6[66]},
      {stage4_6[20]}
   );
   gpc1_1 gpc10128 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc10129 (
      {stage3_7[36]},
      {stage4_7[21]}
   );
   gpc1_1 gpc10130 (
      {stage3_7[37]},
      {stage4_7[22]}
   );
   gpc1_1 gpc10131 (
      {stage3_7[38]},
      {stage4_7[23]}
   );
   gpc1_1 gpc10132 (
      {stage3_7[39]},
      {stage4_7[24]}
   );
   gpc1_1 gpc10133 (
      {stage3_7[40]},
      {stage4_7[25]}
   );
   gpc1_1 gpc10134 (
      {stage3_7[41]},
      {stage4_7[26]}
   );
   gpc1_1 gpc10135 (
      {stage3_7[42]},
      {stage4_7[27]}
   );
   gpc1_1 gpc10136 (
      {stage3_7[43]},
      {stage4_7[28]}
   );
   gpc1_1 gpc10137 (
      {stage3_7[44]},
      {stage4_7[29]}
   );
   gpc1_1 gpc10138 (
      {stage3_7[45]},
      {stage4_7[30]}
   );
   gpc1_1 gpc10139 (
      {stage3_7[46]},
      {stage4_7[31]}
   );
   gpc1_1 gpc10140 (
      {stage3_7[47]},
      {stage4_7[32]}
   );
   gpc1_1 gpc10141 (
      {stage3_7[48]},
      {stage4_7[33]}
   );
   gpc1_1 gpc10142 (
      {stage3_7[49]},
      {stage4_7[34]}
   );
   gpc1_1 gpc10143 (
      {stage3_7[50]},
      {stage4_7[35]}
   );
   gpc1_1 gpc10144 (
      {stage3_7[51]},
      {stage4_7[36]}
   );
   gpc1_1 gpc10145 (
      {stage3_7[52]},
      {stage4_7[37]}
   );
   gpc1_1 gpc10146 (
      {stage3_7[53]},
      {stage4_7[38]}
   );
   gpc1_1 gpc10147 (
      {stage3_7[54]},
      {stage4_7[39]}
   );
   gpc1_1 gpc10148 (
      {stage3_8[29]},
      {stage4_8[17]}
   );
   gpc1_1 gpc10149 (
      {stage3_8[30]},
      {stage4_8[18]}
   );
   gpc1_1 gpc10150 (
      {stage3_8[31]},
      {stage4_8[19]}
   );
   gpc1_1 gpc10151 (
      {stage3_8[32]},
      {stage4_8[20]}
   );
   gpc1_1 gpc10152 (
      {stage3_8[33]},
      {stage4_8[21]}
   );
   gpc1_1 gpc10153 (
      {stage3_8[34]},
      {stage4_8[22]}
   );
   gpc1_1 gpc10154 (
      {stage3_8[35]},
      {stage4_8[23]}
   );
   gpc1_1 gpc10155 (
      {stage3_8[36]},
      {stage4_8[24]}
   );
   gpc1_1 gpc10156 (
      {stage3_8[37]},
      {stage4_8[25]}
   );
   gpc1_1 gpc10157 (
      {stage3_8[38]},
      {stage4_8[26]}
   );
   gpc1_1 gpc10158 (
      {stage3_8[39]},
      {stage4_8[27]}
   );
   gpc1_1 gpc10159 (
      {stage3_8[40]},
      {stage4_8[28]}
   );
   gpc1_1 gpc10160 (
      {stage3_8[41]},
      {stage4_8[29]}
   );
   gpc1_1 gpc10161 (
      {stage3_8[42]},
      {stage4_8[30]}
   );
   gpc1_1 gpc10162 (
      {stage3_8[43]},
      {stage4_8[31]}
   );
   gpc1_1 gpc10163 (
      {stage3_8[44]},
      {stage4_8[32]}
   );
   gpc1_1 gpc10164 (
      {stage3_8[45]},
      {stage4_8[33]}
   );
   gpc1_1 gpc10165 (
      {stage3_8[46]},
      {stage4_8[34]}
   );
   gpc1_1 gpc10166 (
      {stage3_10[65]},
      {stage4_10[26]}
   );
   gpc1_1 gpc10167 (
      {stage3_10[66]},
      {stage4_10[27]}
   );
   gpc1_1 gpc10168 (
      {stage3_10[67]},
      {stage4_10[28]}
   );
   gpc1_1 gpc10169 (
      {stage3_11[52]},
      {stage4_11[25]}
   );
   gpc1_1 gpc10170 (
      {stage3_11[53]},
      {stage4_11[26]}
   );
   gpc1_1 gpc10171 (
      {stage3_11[54]},
      {stage4_11[27]}
   );
   gpc1_1 gpc10172 (
      {stage3_11[55]},
      {stage4_11[28]}
   );
   gpc1_1 gpc10173 (
      {stage3_11[56]},
      {stage4_11[29]}
   );
   gpc1_1 gpc10174 (
      {stage3_11[57]},
      {stage4_11[30]}
   );
   gpc1_1 gpc10175 (
      {stage3_11[58]},
      {stage4_11[31]}
   );
   gpc1_1 gpc10176 (
      {stage3_11[59]},
      {stage4_11[32]}
   );
   gpc1_1 gpc10177 (
      {stage3_11[60]},
      {stage4_11[33]}
   );
   gpc1_1 gpc10178 (
      {stage3_13[43]},
      {stage4_13[24]}
   );
   gpc1_1 gpc10179 (
      {stage3_13[44]},
      {stage4_13[25]}
   );
   gpc1_1 gpc10180 (
      {stage3_13[45]},
      {stage4_13[26]}
   );
   gpc1_1 gpc10181 (
      {stage3_13[46]},
      {stage4_13[27]}
   );
   gpc1_1 gpc10182 (
      {stage3_14[31]},
      {stage4_14[26]}
   );
   gpc1_1 gpc10183 (
      {stage3_14[32]},
      {stage4_14[27]}
   );
   gpc1_1 gpc10184 (
      {stage3_14[33]},
      {stage4_14[28]}
   );
   gpc1_1 gpc10185 (
      {stage3_14[34]},
      {stage4_14[29]}
   );
   gpc1_1 gpc10186 (
      {stage3_15[45]},
      {stage4_15[17]}
   );
   gpc1_1 gpc10187 (
      {stage3_15[46]},
      {stage4_15[18]}
   );
   gpc1_1 gpc10188 (
      {stage3_15[47]},
      {stage4_15[19]}
   );
   gpc1_1 gpc10189 (
      {stage3_15[48]},
      {stage4_15[20]}
   );
   gpc1_1 gpc10190 (
      {stage3_15[49]},
      {stage4_15[21]}
   );
   gpc1_1 gpc10191 (
      {stage3_15[50]},
      {stage4_15[22]}
   );
   gpc1_1 gpc10192 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc10193 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc10194 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc10195 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc10196 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc10197 (
      {stage3_16[45]},
      {stage4_16[19]}
   );
   gpc1_1 gpc10198 (
      {stage3_16[46]},
      {stage4_16[20]}
   );
   gpc1_1 gpc10199 (
      {stage3_16[47]},
      {stage4_16[21]}
   );
   gpc1_1 gpc10200 (
      {stage3_16[48]},
      {stage4_16[22]}
   );
   gpc1_1 gpc10201 (
      {stage3_16[49]},
      {stage4_16[23]}
   );
   gpc1_1 gpc10202 (
      {stage3_16[50]},
      {stage4_16[24]}
   );
   gpc1_1 gpc10203 (
      {stage3_16[51]},
      {stage4_16[25]}
   );
   gpc1_1 gpc10204 (
      {stage3_16[52]},
      {stage4_16[26]}
   );
   gpc1_1 gpc10205 (
      {stage3_16[53]},
      {stage4_16[27]}
   );
   gpc1_1 gpc10206 (
      {stage3_16[54]},
      {stage4_16[28]}
   );
   gpc1_1 gpc10207 (
      {stage3_16[55]},
      {stage4_16[29]}
   );
   gpc1_1 gpc10208 (
      {stage3_16[56]},
      {stage4_16[30]}
   );
   gpc1_1 gpc10209 (
      {stage3_16[57]},
      {stage4_16[31]}
   );
   gpc1_1 gpc10210 (
      {stage3_16[58]},
      {stage4_16[32]}
   );
   gpc1_1 gpc10211 (
      {stage3_17[36]},
      {stage4_17[15]}
   );
   gpc1_1 gpc10212 (
      {stage3_17[37]},
      {stage4_17[16]}
   );
   gpc1_1 gpc10213 (
      {stage3_17[38]},
      {stage4_17[17]}
   );
   gpc1_1 gpc10214 (
      {stage3_17[39]},
      {stage4_17[18]}
   );
   gpc1_1 gpc10215 (
      {stage3_17[40]},
      {stage4_17[19]}
   );
   gpc1_1 gpc10216 (
      {stage3_17[41]},
      {stage4_17[20]}
   );
   gpc1_1 gpc10217 (
      {stage3_17[42]},
      {stage4_17[21]}
   );
   gpc1_1 gpc10218 (
      {stage3_17[43]},
      {stage4_17[22]}
   );
   gpc1_1 gpc10219 (
      {stage3_18[52]},
      {stage4_18[20]}
   );
   gpc1_1 gpc10220 (
      {stage3_18[53]},
      {stage4_18[21]}
   );
   gpc1_1 gpc10221 (
      {stage3_18[54]},
      {stage4_18[22]}
   );
   gpc1_1 gpc10222 (
      {stage3_18[55]},
      {stage4_18[23]}
   );
   gpc1_1 gpc10223 (
      {stage3_18[56]},
      {stage4_18[24]}
   );
   gpc1_1 gpc10224 (
      {stage3_18[57]},
      {stage4_18[25]}
   );
   gpc1_1 gpc10225 (
      {stage3_18[58]},
      {stage4_18[26]}
   );
   gpc1_1 gpc10226 (
      {stage3_18[59]},
      {stage4_18[27]}
   );
   gpc1_1 gpc10227 (
      {stage3_18[60]},
      {stage4_18[28]}
   );
   gpc1_1 gpc10228 (
      {stage3_18[61]},
      {stage4_18[29]}
   );
   gpc1_1 gpc10229 (
      {stage3_18[62]},
      {stage4_18[30]}
   );
   gpc1_1 gpc10230 (
      {stage3_18[63]},
      {stage4_18[31]}
   );
   gpc1_1 gpc10231 (
      {stage3_20[57]},
      {stage4_20[21]}
   );
   gpc1_1 gpc10232 (
      {stage3_21[61]},
      {stage4_21[25]}
   );
   gpc1_1 gpc10233 (
      {stage3_21[62]},
      {stage4_21[26]}
   );
   gpc1_1 gpc10234 (
      {stage3_24[29]},
      {stage4_24[18]}
   );
   gpc1_1 gpc10235 (
      {stage3_24[30]},
      {stage4_24[19]}
   );
   gpc1_1 gpc10236 (
      {stage3_24[31]},
      {stage4_24[20]}
   );
   gpc1_1 gpc10237 (
      {stage3_24[32]},
      {stage4_24[21]}
   );
   gpc1_1 gpc10238 (
      {stage3_24[33]},
      {stage4_24[22]}
   );
   gpc1_1 gpc10239 (
      {stage3_24[34]},
      {stage4_24[23]}
   );
   gpc1_1 gpc10240 (
      {stage3_25[48]},
      {stage4_25[16]}
   );
   gpc1_1 gpc10241 (
      {stage3_25[49]},
      {stage4_25[17]}
   );
   gpc1_1 gpc10242 (
      {stage3_25[50]},
      {stage4_25[18]}
   );
   gpc1_1 gpc10243 (
      {stage3_25[51]},
      {stage4_25[19]}
   );
   gpc1_1 gpc10244 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc10245 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc10246 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc10247 (
      {stage3_28[57]},
      {stage4_28[19]}
   );
   gpc1_1 gpc10248 (
      {stage3_28[58]},
      {stage4_28[20]}
   );
   gpc1_1 gpc10249 (
      {stage3_28[59]},
      {stage4_28[21]}
   );
   gpc1_1 gpc10250 (
      {stage3_28[60]},
      {stage4_28[22]}
   );
   gpc1_1 gpc10251 (
      {stage3_28[61]},
      {stage4_28[23]}
   );
   gpc1_1 gpc10252 (
      {stage3_28[62]},
      {stage4_28[24]}
   );
   gpc1_1 gpc10253 (
      {stage3_28[63]},
      {stage4_28[25]}
   );
   gpc1_1 gpc10254 (
      {stage3_28[64]},
      {stage4_28[26]}
   );
   gpc1_1 gpc10255 (
      {stage3_28[65]},
      {stage4_28[27]}
   );
   gpc1_1 gpc10256 (
      {stage3_28[66]},
      {stage4_28[28]}
   );
   gpc1_1 gpc10257 (
      {stage3_28[67]},
      {stage4_28[29]}
   );
   gpc1_1 gpc10258 (
      {stage3_28[68]},
      {stage4_28[30]}
   );
   gpc1_1 gpc10259 (
      {stage3_28[69]},
      {stage4_28[31]}
   );
   gpc1_1 gpc10260 (
      {stage3_30[36]},
      {stage4_30[23]}
   );
   gpc1_1 gpc10261 (
      {stage3_30[37]},
      {stage4_30[24]}
   );
   gpc1_1 gpc10262 (
      {stage3_30[38]},
      {stage4_30[25]}
   );
   gpc1_1 gpc10263 (
      {stage3_32[51]},
      {stage4_32[19]}
   );
   gpc1_1 gpc10264 (
      {stage3_32[52]},
      {stage4_32[20]}
   );
   gpc1_1 gpc10265 (
      {stage3_32[53]},
      {stage4_32[21]}
   );
   gpc1_1 gpc10266 (
      {stage3_32[54]},
      {stage4_32[22]}
   );
   gpc1_1 gpc10267 (
      {stage3_32[55]},
      {stage4_32[23]}
   );
   gpc1_1 gpc10268 (
      {stage3_33[53]},
      {stage4_33[24]}
   );
   gpc1_1 gpc10269 (
      {stage3_33[54]},
      {stage4_33[25]}
   );
   gpc1_1 gpc10270 (
      {stage3_33[55]},
      {stage4_33[26]}
   );
   gpc1_1 gpc10271 (
      {stage3_33[56]},
      {stage4_33[27]}
   );
   gpc1_1 gpc10272 (
      {stage3_33[57]},
      {stage4_33[28]}
   );
   gpc1_1 gpc10273 (
      {stage3_33[58]},
      {stage4_33[29]}
   );
   gpc1_1 gpc10274 (
      {stage3_33[59]},
      {stage4_33[30]}
   );
   gpc1_1 gpc10275 (
      {stage3_33[60]},
      {stage4_33[31]}
   );
   gpc1_1 gpc10276 (
      {stage3_33[61]},
      {stage4_33[32]}
   );
   gpc1_1 gpc10277 (
      {stage3_33[62]},
      {stage4_33[33]}
   );
   gpc1_1 gpc10278 (
      {stage3_34[32]},
      {stage4_34[17]}
   );
   gpc1_1 gpc10279 (
      {stage3_34[33]},
      {stage4_34[18]}
   );
   gpc1_1 gpc10280 (
      {stage3_34[34]},
      {stage4_34[19]}
   );
   gpc1_1 gpc10281 (
      {stage3_34[35]},
      {stage4_34[20]}
   );
   gpc1_1 gpc10282 (
      {stage3_34[36]},
      {stage4_34[21]}
   );
   gpc1_1 gpc10283 (
      {stage3_34[37]},
      {stage4_34[22]}
   );
   gpc1_1 gpc10284 (
      {stage3_34[38]},
      {stage4_34[23]}
   );
   gpc1_1 gpc10285 (
      {stage3_34[39]},
      {stage4_34[24]}
   );
   gpc1_1 gpc10286 (
      {stage3_34[40]},
      {stage4_34[25]}
   );
   gpc1_1 gpc10287 (
      {stage3_34[41]},
      {stage4_34[26]}
   );
   gpc1_1 gpc10288 (
      {stage3_34[42]},
      {stage4_34[27]}
   );
   gpc1_1 gpc10289 (
      {stage3_34[43]},
      {stage4_34[28]}
   );
   gpc1_1 gpc10290 (
      {stage3_34[44]},
      {stage4_34[29]}
   );
   gpc1_1 gpc10291 (
      {stage3_35[52]},
      {stage4_35[19]}
   );
   gpc1_1 gpc10292 (
      {stage3_35[53]},
      {stage4_35[20]}
   );
   gpc1_1 gpc10293 (
      {stage3_35[54]},
      {stage4_35[21]}
   );
   gpc1_1 gpc10294 (
      {stage3_35[55]},
      {stage4_35[22]}
   );
   gpc1_1 gpc10295 (
      {stage3_35[56]},
      {stage4_35[23]}
   );
   gpc1_1 gpc10296 (
      {stage3_36[39]},
      {stage4_36[21]}
   );
   gpc1_1 gpc10297 (
      {stage3_36[40]},
      {stage4_36[22]}
   );
   gpc1_1 gpc10298 (
      {stage3_36[41]},
      {stage4_36[23]}
   );
   gpc1_1 gpc10299 (
      {stage3_36[42]},
      {stage4_36[24]}
   );
   gpc1_1 gpc10300 (
      {stage3_36[43]},
      {stage4_36[25]}
   );
   gpc1_1 gpc10301 (
      {stage3_36[44]},
      {stage4_36[26]}
   );
   gpc1_1 gpc10302 (
      {stage3_36[45]},
      {stage4_36[27]}
   );
   gpc1_1 gpc10303 (
      {stage3_36[46]},
      {stage4_36[28]}
   );
   gpc1_1 gpc10304 (
      {stage3_36[47]},
      {stage4_36[29]}
   );
   gpc1_1 gpc10305 (
      {stage3_36[48]},
      {stage4_36[30]}
   );
   gpc1_1 gpc10306 (
      {stage3_36[49]},
      {stage4_36[31]}
   );
   gpc1_1 gpc10307 (
      {stage3_36[50]},
      {stage4_36[32]}
   );
   gpc1_1 gpc10308 (
      {stage3_36[51]},
      {stage4_36[33]}
   );
   gpc1_1 gpc10309 (
      {stage3_36[52]},
      {stage4_36[34]}
   );
   gpc1_1 gpc10310 (
      {stage3_36[53]},
      {stage4_36[35]}
   );
   gpc1_1 gpc10311 (
      {stage3_36[54]},
      {stage4_36[36]}
   );
   gpc1_1 gpc10312 (
      {stage3_36[55]},
      {stage4_36[37]}
   );
   gpc1_1 gpc10313 (
      {stage3_38[60]},
      {stage4_38[18]}
   );
   gpc1_1 gpc10314 (
      {stage3_38[61]},
      {stage4_38[19]}
   );
   gpc1_1 gpc10315 (
      {stage3_38[62]},
      {stage4_38[20]}
   );
   gpc1_1 gpc10316 (
      {stage3_38[63]},
      {stage4_38[21]}
   );
   gpc1_1 gpc10317 (
      {stage3_38[64]},
      {stage4_38[22]}
   );
   gpc1_1 gpc10318 (
      {stage3_38[65]},
      {stage4_38[23]}
   );
   gpc1_1 gpc10319 (
      {stage3_38[66]},
      {stage4_38[24]}
   );
   gpc1_1 gpc10320 (
      {stage3_38[67]},
      {stage4_38[25]}
   );
   gpc1_1 gpc10321 (
      {stage3_38[68]},
      {stage4_38[26]}
   );
   gpc1_1 gpc10322 (
      {stage3_40[36]},
      {stage4_40[19]}
   );
   gpc1_1 gpc10323 (
      {stage3_40[37]},
      {stage4_40[20]}
   );
   gpc1_1 gpc10324 (
      {stage3_40[38]},
      {stage4_40[21]}
   );
   gpc1_1 gpc10325 (
      {stage3_40[39]},
      {stage4_40[22]}
   );
   gpc1_1 gpc10326 (
      {stage3_40[40]},
      {stage4_40[23]}
   );
   gpc1_1 gpc10327 (
      {stage3_40[41]},
      {stage4_40[24]}
   );
   gpc1_1 gpc10328 (
      {stage3_40[42]},
      {stage4_40[25]}
   );
   gpc1_1 gpc10329 (
      {stage3_40[43]},
      {stage4_40[26]}
   );
   gpc1_1 gpc10330 (
      {stage3_40[44]},
      {stage4_40[27]}
   );
   gpc1_1 gpc10331 (
      {stage3_40[45]},
      {stage4_40[28]}
   );
   gpc1_1 gpc10332 (
      {stage3_41[54]},
      {stage4_41[21]}
   );
   gpc1_1 gpc10333 (
      {stage3_41[55]},
      {stage4_41[22]}
   );
   gpc1_1 gpc10334 (
      {stage3_41[56]},
      {stage4_41[23]}
   );
   gpc1_1 gpc10335 (
      {stage3_43[55]},
      {stage4_43[18]}
   );
   gpc1_1 gpc10336 (
      {stage3_43[56]},
      {stage4_43[19]}
   );
   gpc1_1 gpc10337 (
      {stage3_43[57]},
      {stage4_43[20]}
   );
   gpc1_1 gpc10338 (
      {stage3_43[58]},
      {stage4_43[21]}
   );
   gpc1_1 gpc10339 (
      {stage3_43[59]},
      {stage4_43[22]}
   );
   gpc1_1 gpc10340 (
      {stage3_44[68]},
      {stage4_44[23]}
   );
   gpc1_1 gpc10341 (
      {stage3_44[69]},
      {stage4_44[24]}
   );
   gpc1_1 gpc10342 (
      {stage3_44[70]},
      {stage4_44[25]}
   );
   gpc1_1 gpc10343 (
      {stage3_44[71]},
      {stage4_44[26]}
   );
   gpc1_1 gpc10344 (
      {stage3_44[72]},
      {stage4_44[27]}
   );
   gpc1_1 gpc10345 (
      {stage3_44[73]},
      {stage4_44[28]}
   );
   gpc1_1 gpc10346 (
      {stage3_44[74]},
      {stage4_44[29]}
   );
   gpc1_1 gpc10347 (
      {stage3_44[75]},
      {stage4_44[30]}
   );
   gpc1_1 gpc10348 (
      {stage3_44[76]},
      {stage4_44[31]}
   );
   gpc1_1 gpc10349 (
      {stage3_44[77]},
      {stage4_44[32]}
   );
   gpc1_1 gpc10350 (
      {stage3_44[78]},
      {stage4_44[33]}
   );
   gpc1_1 gpc10351 (
      {stage3_44[79]},
      {stage4_44[34]}
   );
   gpc1_1 gpc10352 (
      {stage3_44[80]},
      {stage4_44[35]}
   );
   gpc1_1 gpc10353 (
      {stage3_44[81]},
      {stage4_44[36]}
   );
   gpc1_1 gpc10354 (
      {stage3_44[82]},
      {stage4_44[37]}
   );
   gpc1_1 gpc10355 (
      {stage3_44[83]},
      {stage4_44[38]}
   );
   gpc1_1 gpc10356 (
      {stage3_44[84]},
      {stage4_44[39]}
   );
   gpc1_1 gpc10357 (
      {stage3_46[46]},
      {stage4_46[22]}
   );
   gpc1_1 gpc10358 (
      {stage3_46[47]},
      {stage4_46[23]}
   );
   gpc1_1 gpc10359 (
      {stage3_46[48]},
      {stage4_46[24]}
   );
   gpc1_1 gpc10360 (
      {stage3_47[71]},
      {stage4_47[23]}
   );
   gpc1_1 gpc10361 (
      {stage3_47[72]},
      {stage4_47[24]}
   );
   gpc1_1 gpc10362 (
      {stage3_47[73]},
      {stage4_47[25]}
   );
   gpc1_1 gpc10363 (
      {stage3_49[54]},
      {stage4_49[17]}
   );
   gpc1_1 gpc10364 (
      {stage3_49[55]},
      {stage4_49[18]}
   );
   gpc1_1 gpc10365 (
      {stage3_49[56]},
      {stage4_49[19]}
   );
   gpc1_1 gpc10366 (
      {stage3_49[57]},
      {stage4_49[20]}
   );
   gpc1_1 gpc10367 (
      {stage3_49[58]},
      {stage4_49[21]}
   );
   gpc1_1 gpc10368 (
      {stage3_49[59]},
      {stage4_49[22]}
   );
   gpc1_1 gpc10369 (
      {stage3_49[60]},
      {stage4_49[23]}
   );
   gpc1_1 gpc10370 (
      {stage3_49[61]},
      {stage4_49[24]}
   );
   gpc1_1 gpc10371 (
      {stage3_49[62]},
      {stage4_49[25]}
   );
   gpc1_1 gpc10372 (
      {stage3_49[63]},
      {stage4_49[26]}
   );
   gpc1_1 gpc10373 (
      {stage3_49[64]},
      {stage4_49[27]}
   );
   gpc1_1 gpc10374 (
      {stage3_50[63]},
      {stage4_50[23]}
   );
   gpc1_1 gpc10375 (
      {stage3_52[54]},
      {stage4_52[21]}
   );
   gpc1_1 gpc10376 (
      {stage3_52[55]},
      {stage4_52[22]}
   );
   gpc1_1 gpc10377 (
      {stage3_54[54]},
      {stage4_54[22]}
   );
   gpc1_1 gpc10378 (
      {stage3_54[55]},
      {stage4_54[23]}
   );
   gpc1_1 gpc10379 (
      {stage3_54[56]},
      {stage4_54[24]}
   );
   gpc1_1 gpc10380 (
      {stage3_54[57]},
      {stage4_54[25]}
   );
   gpc1_1 gpc10381 (
      {stage3_54[58]},
      {stage4_54[26]}
   );
   gpc1_1 gpc10382 (
      {stage3_54[59]},
      {stage4_54[27]}
   );
   gpc1_1 gpc10383 (
      {stage3_54[60]},
      {stage4_54[28]}
   );
   gpc1_1 gpc10384 (
      {stage3_54[61]},
      {stage4_54[29]}
   );
   gpc1_1 gpc10385 (
      {stage3_54[62]},
      {stage4_54[30]}
   );
   gpc1_1 gpc10386 (
      {stage3_55[40]},
      {stage4_55[22]}
   );
   gpc1_1 gpc10387 (
      {stage3_55[41]},
      {stage4_55[23]}
   );
   gpc1_1 gpc10388 (
      {stage3_55[42]},
      {stage4_55[24]}
   );
   gpc1_1 gpc10389 (
      {stage3_55[43]},
      {stage4_55[25]}
   );
   gpc1_1 gpc10390 (
      {stage3_55[44]},
      {stage4_55[26]}
   );
   gpc1_1 gpc10391 (
      {stage3_55[45]},
      {stage4_55[27]}
   );
   gpc1_1 gpc10392 (
      {stage3_55[46]},
      {stage4_55[28]}
   );
   gpc1_1 gpc10393 (
      {stage3_56[26]},
      {stage4_56[16]}
   );
   gpc1_1 gpc10394 (
      {stage3_56[27]},
      {stage4_56[17]}
   );
   gpc1_1 gpc10395 (
      {stage3_56[28]},
      {stage4_56[18]}
   );
   gpc1_1 gpc10396 (
      {stage3_56[29]},
      {stage4_56[19]}
   );
   gpc1_1 gpc10397 (
      {stage3_56[30]},
      {stage4_56[20]}
   );
   gpc1_1 gpc10398 (
      {stage3_56[31]},
      {stage4_56[21]}
   );
   gpc1_1 gpc10399 (
      {stage3_56[32]},
      {stage4_56[22]}
   );
   gpc1_1 gpc10400 (
      {stage3_56[33]},
      {stage4_56[23]}
   );
   gpc1_1 gpc10401 (
      {stage3_56[34]},
      {stage4_56[24]}
   );
   gpc1_1 gpc10402 (
      {stage3_56[35]},
      {stage4_56[25]}
   );
   gpc1_1 gpc10403 (
      {stage3_56[36]},
      {stage4_56[26]}
   );
   gpc1_1 gpc10404 (
      {stage3_56[37]},
      {stage4_56[27]}
   );
   gpc1_1 gpc10405 (
      {stage3_56[38]},
      {stage4_56[28]}
   );
   gpc1_1 gpc10406 (
      {stage3_57[51]},
      {stage4_57[23]}
   );
   gpc1_1 gpc10407 (
      {stage3_57[52]},
      {stage4_57[24]}
   );
   gpc1_1 gpc10408 (
      {stage3_58[48]},
      {stage4_58[15]}
   );
   gpc1_1 gpc10409 (
      {stage3_59[45]},
      {stage4_59[15]}
   );
   gpc1_1 gpc10410 (
      {stage3_60[49]},
      {stage4_60[21]}
   );
   gpc1_1 gpc10411 (
      {stage3_60[50]},
      {stage4_60[22]}
   );
   gpc1_1 gpc10412 (
      {stage3_60[51]},
      {stage4_60[23]}
   );
   gpc1_1 gpc10413 (
      {stage3_60[52]},
      {stage4_60[24]}
   );
   gpc1_1 gpc10414 (
      {stage3_61[55]},
      {stage4_61[27]}
   );
   gpc1_1 gpc10415 (
      {stage3_61[56]},
      {stage4_61[28]}
   );
   gpc1_1 gpc10416 (
      {stage3_62[34]},
      {stage4_62[17]}
   );
   gpc1_1 gpc10417 (
      {stage3_62[35]},
      {stage4_62[18]}
   );
   gpc1_1 gpc10418 (
      {stage3_62[36]},
      {stage4_62[19]}
   );
   gpc1_1 gpc10419 (
      {stage3_62[37]},
      {stage4_62[20]}
   );
   gpc1_1 gpc10420 (
      {stage3_62[38]},
      {stage4_62[21]}
   );
   gpc1_1 gpc10421 (
      {stage3_62[39]},
      {stage4_62[22]}
   );
   gpc1_1 gpc10422 (
      {stage3_62[40]},
      {stage4_62[23]}
   );
   gpc1_1 gpc10423 (
      {stage3_67[13]},
      {stage4_67[15]}
   );
   gpc1_1 gpc10424 (
      {stage3_67[14]},
      {stage4_67[16]}
   );
   gpc606_5 gpc10425 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1406_5 gpc10426 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc1163_5 gpc10427 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[4]},
      {stage4_5[1]},
      {stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc606_5 gpc10428 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16], stage4_3[17]},
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage5_7[0],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc606_5 gpc10429 (
      {stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[1],stage5_6[3],stage5_5[4],stage5_4[4]}
   );
   gpc606_5 gpc10430 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[2],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc10431 (
      {stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21], stage4_4[22]},
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17]},
      {stage5_8[2],stage5_7[3],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc606_5 gpc10432 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc10433 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc10434 (
      {stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24], stage4_5[25]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[5],stage5_7[6],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc10435 (
      {stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage4_7[18], stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23]},
      {stage5_9[3],stage5_8[6],stage5_7[7],stage5_6[9],stage5_5[10]}
   );
   gpc606_5 gpc10436 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37]},
      {stage4_7[24], stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29]},
      {stage5_9[4],stage5_8[7],stage5_7[8],stage5_6[10],stage5_5[11]}
   );
   gpc615_5 gpc10437 (
      {stage4_7[30], stage4_7[31], stage4_7[32], stage4_7[33], stage4_7[34]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[5],stage5_8[8],stage5_7[9]}
   );
   gpc615_5 gpc10438 (
      {stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38], stage4_7[39]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[6],stage5_8[9],stage5_7[10]}
   );
   gpc1406_5 gpc10439 (
      {stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[7],stage5_8[10]}
   );
   gpc215_4 gpc10440 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage5_11[3],stage5_10[3],stage5_9[8],stage5_8[11]}
   );
   gpc215_4 gpc10441 (
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[13]},
      {stage4_10[6], stage4_10[7]},
      {stage5_11[4],stage5_10[4],stage5_9[9],stage5_8[12]}
   );
   gpc207_4 gpc10442 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24]},
      {stage4_10[8], stage4_10[9]},
      {stage5_11[5],stage5_10[5],stage5_9[10],stage5_8[13]}
   );
   gpc606_5 gpc10443 (
      {stage4_8[25], stage4_8[26], stage4_8[27], stage4_8[28], stage4_8[29], stage4_8[30]},
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15]},
      {stage5_12[1],stage5_11[6],stage5_10[6],stage5_9[11],stage5_8[14]}
   );
   gpc606_5 gpc10444 (
      {stage4_8[31], stage4_8[32], stage4_8[33], stage4_8[34], 1'b0, 1'b0},
      {stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19], stage4_10[20], stage4_10[21]},
      {stage5_12[2],stage5_11[7],stage5_10[7],stage5_9[12],stage5_8[15]}
   );
   gpc1163_5 gpc10445 (
      {stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[0]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[3],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc10446 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], 1'b0},
      {stage4_11[7]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[1],stage5_12[4],stage5_11[9],stage5_10[9]}
   );
   gpc615_5 gpc10447 (
      {stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12]},
      {stage4_12[7]},
      {stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[5],stage5_11[10]}
   );
   gpc615_5 gpc10448 (
      {stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage4_12[8]},
      {stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[6],stage5_11[11]}
   );
   gpc615_5 gpc10449 (
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22]},
      {stage4_12[9]},
      {stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[7],stage5_11[12]}
   );
   gpc615_5 gpc10450 (
      {stage4_11[23], stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27]},
      {stage4_12[10]},
      {stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[8],stage5_11[13]}
   );
   gpc615_5 gpc10451 (
      {stage4_12[11], stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15]},
      {stage4_13[25]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[9]}
   );
   gpc615_5 gpc10452 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc10453 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc10454 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc10455 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[10]}
   );
   gpc615_5 gpc10456 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc10457 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc10458 (
      {stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc606_5 gpc10459 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7],stage5_17[7]}
   );
   gpc2116_5 gpc10460 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[6]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc2116_5 gpc10461 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[1]},
      {stage4_21[2], stage4_21[3]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc2116_5 gpc10462 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[8]},
      {stage4_20[2]},
      {stage4_21[4], stage4_21[5]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc10463 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[9]},
      {stage4_20[3], stage4_20[4], stage4_20[5], stage4_20[6], stage4_20[7], stage4_20[8]},
      {stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[7],stage5_18[11]}
   );
   gpc615_5 gpc10464 (
      {stage4_18[23], stage4_18[24], stage4_18[25], stage4_18[26], stage4_18[27]},
      {stage4_19[10]},
      {stage4_20[9], stage4_20[10], stage4_20[11], stage4_20[12], stage4_20[13], stage4_20[14]},
      {stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[8],stage5_18[12]}
   );
   gpc615_5 gpc10465 (
      {stage4_18[28], stage4_18[29], stage4_18[30], stage4_18[31], 1'b0},
      {stage4_19[11]},
      {stage4_20[15], stage4_20[16], stage4_20[17], stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[9],stage5_18[13]}
   );
   gpc615_5 gpc10466 (
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16]},
      {stage4_20[21]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[0],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc7_3 gpc10467 (
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[1],stage5_22[7],stage5_21[8]}
   );
   gpc7_3 gpc10468 (
      {stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23], stage4_21[24], stage4_21[25]},
      {stage5_23[2],stage5_22[8],stage5_21[9]}
   );
   gpc1163_5 gpc10469 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[3],stage5_22[9]}
   );
   gpc1163_5 gpc10470 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage4_24[1]},
      {stage4_25[1]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[4],stage5_22[10]}
   );
   gpc1163_5 gpc10471 (
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[2]},
      {stage4_25[2]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[5],stage5_22[11]}
   );
   gpc615_5 gpc10472 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[18]},
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[6],stage5_22[12]}
   );
   gpc615_5 gpc10473 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[19]},
      {stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12], stage4_24[13], stage4_24[14]},
      {stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[7],stage5_22[13]}
   );
   gpc615_5 gpc10474 (
      {stage4_22[19], stage4_22[20], 1'b0, 1'b0, 1'b0},
      {stage4_23[20]},
      {stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18], stage4_24[19], stage4_24[20]},
      {stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[8],stage5_22[14]}
   );
   gpc606_5 gpc10475 (
      {stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[6],stage5_25[6]}
   );
   gpc606_5 gpc10476 (
      {stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12], stage4_25[13], stage4_25[14]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[7],stage5_25[7]}
   );
   gpc207_4 gpc10477 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[8]}
   );
   gpc207_4 gpc10478 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {stage4_28[2], stage4_28[3]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[9]}
   );
   gpc615_5 gpc10479 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_28[4]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4]}
   );
   gpc606_5 gpc10480 (
      {stage4_28[5], stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[5],stage5_28[5]}
   );
   gpc606_5 gpc10481 (
      {stage4_28[11], stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[6],stage5_28[6]}
   );
   gpc606_5 gpc10482 (
      {stage4_28[17], stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[3],stage5_30[3],stage5_29[7],stage5_28[7]}
   );
   gpc606_5 gpc10483 (
      {stage4_28[23], stage4_28[24], stage4_28[25], stage4_28[26], stage4_28[27], stage4_28[28]},
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23]},
      {stage5_32[3],stage5_31[4],stage5_30[4],stage5_29[8],stage5_28[8]}
   );
   gpc207_4 gpc10484 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[4],stage5_31[5],stage5_30[5],stage5_29[9]}
   );
   gpc207_4 gpc10485 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17], stage4_29[18], stage4_29[19]},
      {stage4_31[2], stage4_31[3]},
      {stage5_32[5],stage5_31[6],stage5_30[6],stage5_29[10]}
   );
   gpc615_5 gpc10486 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[0]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[6],stage5_31[7]}
   );
   gpc615_5 gpc10487 (
      {stage4_31[9], stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13]},
      {stage4_32[1]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[1],stage5_33[1],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc10488 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[2],stage5_34[2],stage5_33[2],stage5_32[8]}
   );
   gpc606_5 gpc10489 (
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage5_36[1],stage5_35[3],stage5_34[3],stage5_33[3],stage5_32[9]}
   );
   gpc606_5 gpc10490 (
      {stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17], stage4_32[18], stage4_32[19]},
      {stage4_34[12], stage4_34[13], stage4_34[14], stage4_34[15], stage4_34[16], stage4_34[17]},
      {stage5_36[2],stage5_35[4],stage5_34[4],stage5_33[4],stage5_32[10]}
   );
   gpc606_5 gpc10491 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[3],stage5_35[5],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc10492 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[4],stage5_35[6],stage5_34[6],stage5_33[6]}
   );
   gpc606_5 gpc10493 (
      {stage4_33[24], stage4_33[25], stage4_33[26], stage4_33[27], stage4_33[28], stage4_33[29]},
      {stage4_35[12], stage4_35[13], stage4_35[14], stage4_35[15], stage4_35[16], stage4_35[17]},
      {stage5_37[2],stage5_36[5],stage5_35[7],stage5_34[7],stage5_33[7]}
   );
   gpc606_5 gpc10494 (
      {stage4_33[30], stage4_33[31], stage4_33[32], stage4_33[33], 1'b0, 1'b0},
      {stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21], stage4_35[22], stage4_35[23]},
      {stage5_37[3],stage5_36[6],stage5_35[8],stage5_34[8],stage5_33[8]}
   );
   gpc1163_5 gpc10495 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[4],stage5_36[7]}
   );
   gpc1163_5 gpc10496 (
      {stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage4_38[1]},
      {stage4_39[1]},
      {stage5_40[1],stage5_39[1],stage5_38[1],stage5_37[5],stage5_36[8]}
   );
   gpc1163_5 gpc10497 (
      {stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], 1'b0, 1'b0},
      {stage4_38[2]},
      {stage4_39[2]},
      {stage5_40[2],stage5_39[2],stage5_38[2],stage5_37[6],stage5_36[9]}
   );
   gpc606_5 gpc10498 (
      {stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12], stage4_36[13], stage4_36[14]},
      {stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6], stage4_38[7], stage4_38[8]},
      {stage5_40[3],stage5_39[3],stage5_38[3],stage5_37[7],stage5_36[10]}
   );
   gpc606_5 gpc10499 (
      {stage4_36[15], stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20]},
      {stage4_38[9], stage4_38[10], stage4_38[11], stage4_38[12], stage4_38[13], stage4_38[14]},
      {stage5_40[4],stage5_39[4],stage5_38[4],stage5_37[8],stage5_36[11]}
   );
   gpc606_5 gpc10500 (
      {stage4_36[21], stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26]},
      {stage4_38[15], stage4_38[16], stage4_38[17], stage4_38[18], stage4_38[19], stage4_38[20]},
      {stage5_40[5],stage5_39[5],stage5_38[5],stage5_37[9],stage5_36[12]}
   );
   gpc606_5 gpc10501 (
      {stage4_36[27], stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32]},
      {stage4_38[21], stage4_38[22], stage4_38[23], stage4_38[24], stage4_38[25], stage4_38[26]},
      {stage5_40[6],stage5_39[6],stage5_38[6],stage5_37[10],stage5_36[13]}
   );
   gpc135_4 gpc10502 (
      {stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6], stage4_39[7]},
      {stage4_40[0], stage4_40[1], stage4_40[2]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[7],stage5_39[7]}
   );
   gpc135_4 gpc10503 (
      {stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12]},
      {stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[8],stage5_39[8]}
   );
   gpc135_4 gpc10504 (
      {stage4_39[13], stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17]},
      {stage4_40[6], stage4_40[7], stage4_40[8]},
      {stage4_41[2]},
      {stage5_42[2],stage5_41[2],stage5_40[9],stage5_39[9]}
   );
   gpc615_5 gpc10505 (
      {stage4_39[18], stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22]},
      {stage4_40[9]},
      {stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7], stage4_41[8]},
      {stage5_43[0],stage5_42[3],stage5_41[3],stage5_40[10],stage5_39[10]}
   );
   gpc606_5 gpc10506 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[4],stage5_41[4],stage5_40[11]}
   );
   gpc606_5 gpc10507 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[2],stage5_42[5],stage5_41[5],stage5_40[12]}
   );
   gpc606_5 gpc10508 (
      {stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13], stage4_41[14]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[3],stage5_42[6],stage5_41[6]}
   );
   gpc606_5 gpc10509 (
      {stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19], stage4_41[20]},
      {stage4_43[6], stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage5_45[1],stage5_44[3],stage5_43[4],stage5_42[7],stage5_41[7]}
   );
   gpc606_5 gpc10510 (
      {stage4_41[21], stage4_41[22], stage4_41[23], 1'b0, 1'b0, 1'b0},
      {stage4_43[12], stage4_43[13], stage4_43[14], stage4_43[15], stage4_43[16], stage4_43[17]},
      {stage5_45[2],stage5_44[4],stage5_43[5],stage5_42[8],stage5_41[8]}
   );
   gpc7_3 gpc10511 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17], stage4_42[18]},
      {stage5_44[5],stage5_43[6],stage5_42[9]}
   );
   gpc615_5 gpc10512 (
      {stage4_43[18], stage4_43[19], stage4_43[20], stage4_43[21], stage4_43[22]},
      {stage4_44[0]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[3],stage5_44[6],stage5_43[7]}
   );
   gpc135_4 gpc10513 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[1],stage5_45[4],stage5_44[7]}
   );
   gpc135_4 gpc10514 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[2],stage5_45[5],stage5_44[8]}
   );
   gpc135_4 gpc10515 (
      {stage4_44[11], stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[3],stage5_45[6],stage5_44[9]}
   );
   gpc135_4 gpc10516 (
      {stage4_44[16], stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20]},
      {stage4_45[15], stage4_45[16], stage4_45[17]},
      {stage4_46[3]},
      {stage5_47[4],stage5_46[4],stage5_45[7],stage5_44[10]}
   );
   gpc135_4 gpc10517 (
      {stage4_44[21], stage4_44[22], stage4_44[23], stage4_44[24], stage4_44[25]},
      {stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_46[4]},
      {stage5_47[5],stage5_46[5],stage5_45[8],stage5_44[11]}
   );
   gpc606_5 gpc10518 (
      {stage4_45[21], stage4_45[22], stage4_45[23], stage4_45[24], stage4_45[25], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[6],stage5_46[6],stage5_45[9]}
   );
   gpc2135_5 gpc10519 (
      {stage4_46[5], stage4_46[6], stage4_46[7], stage4_46[8], stage4_46[9]},
      {stage4_47[6], stage4_47[7], stage4_47[8]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[7],stage5_46[7]}
   );
   gpc2135_5 gpc10520 (
      {stage4_46[10], stage4_46[11], stage4_46[12], stage4_46[13], stage4_46[14]},
      {stage4_47[9], stage4_47[10], stage4_47[11]},
      {stage4_48[1]},
      {stage4_49[2], stage4_49[3]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[8],stage5_46[8]}
   );
   gpc2135_5 gpc10521 (
      {stage4_46[15], stage4_46[16], stage4_46[17], stage4_46[18], stage4_46[19]},
      {stage4_47[12], stage4_47[13], stage4_47[14]},
      {stage4_48[2]},
      {stage4_49[4], stage4_49[5]},
      {stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[9],stage5_46[9]}
   );
   gpc615_5 gpc10522 (
      {stage4_46[20], stage4_46[21], stage4_46[22], stage4_46[23], stage4_46[24]},
      {stage4_47[15]},
      {stage4_48[3], stage4_48[4], stage4_48[5], stage4_48[6], stage4_48[7], stage4_48[8]},
      {stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[10],stage5_46[10]}
   );
   gpc615_5 gpc10523 (
      {stage4_47[16], stage4_47[17], stage4_47[18], stage4_47[19], stage4_47[20]},
      {stage4_48[9]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[0],stage5_50[4],stage5_49[5],stage5_48[5],stage5_47[11]}
   );
   gpc615_5 gpc10524 (
      {stage4_47[21], stage4_47[22], stage4_47[23], stage4_47[24], stage4_47[25]},
      {stage4_48[10]},
      {stage4_49[12], stage4_49[13], stage4_49[14], stage4_49[15], stage4_49[16], stage4_49[17]},
      {stage5_51[1],stage5_50[5],stage5_49[6],stage5_48[6],stage5_47[12]}
   );
   gpc7_3 gpc10525 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[6]}
   );
   gpc7_3 gpc10526 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11], stage4_50[12], stage4_50[13]},
      {stage5_52[1],stage5_51[3],stage5_50[7]}
   );
   gpc615_5 gpc10527 (
      {stage4_50[14], stage4_50[15], stage4_50[16], stage4_50[17], stage4_50[18]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[2],stage5_51[4],stage5_50[8]}
   );
   gpc615_5 gpc10528 (
      {stage4_50[19], stage4_50[20], stage4_50[21], stage4_50[22], stage4_50[23]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[3],stage5_51[5],stage5_50[9]}
   );
   gpc117_4 gpc10529 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6], stage4_51[7], stage4_51[8]},
      {stage4_52[12]},
      {stage4_53[0]},
      {stage5_54[2],stage5_53[2],stage5_52[4],stage5_51[6]}
   );
   gpc606_5 gpc10530 (
      {stage4_51[9], stage4_51[10], stage4_51[11], stage4_51[12], stage4_51[13], stage4_51[14]},
      {stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5], stage4_53[6]},
      {stage5_55[0],stage5_54[3],stage5_53[3],stage5_52[5],stage5_51[7]}
   );
   gpc606_5 gpc10531 (
      {stage4_51[15], stage4_51[16], stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20]},
      {stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11], stage4_53[12]},
      {stage5_55[1],stage5_54[4],stage5_53[4],stage5_52[6],stage5_51[8]}
   );
   gpc606_5 gpc10532 (
      {stage4_51[21], stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17], stage4_53[18]},
      {stage5_55[2],stage5_54[5],stage5_53[5],stage5_52[7],stage5_51[9]}
   );
   gpc606_5 gpc10533 (
      {stage4_52[13], stage4_52[14], stage4_52[15], stage4_52[16], stage4_52[17], stage4_52[18]},
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5]},
      {stage5_56[0],stage5_55[3],stage5_54[6],stage5_53[6],stage5_52[8]}
   );
   gpc606_5 gpc10534 (
      {stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23], stage4_53[24]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[1],stage5_55[4],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc10535 (
      {stage4_54[6], stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10]},
      {stage4_55[6]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[1],stage5_56[2],stage5_55[5],stage5_54[8]}
   );
   gpc615_5 gpc10536 (
      {stage4_54[11], stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15]},
      {stage4_55[7]},
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage5_58[1],stage5_57[2],stage5_56[3],stage5_55[6],stage5_54[9]}
   );
   gpc615_5 gpc10537 (
      {stage4_54[16], stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20]},
      {stage4_55[8]},
      {stage4_56[12], stage4_56[13], stage4_56[14], stage4_56[15], stage4_56[16], stage4_56[17]},
      {stage5_58[2],stage5_57[3],stage5_56[4],stage5_55[7],stage5_54[10]}
   );
   gpc615_5 gpc10538 (
      {stage4_54[21], stage4_54[22], stage4_54[23], stage4_54[24], stage4_54[25]},
      {stage4_55[9]},
      {stage4_56[18], stage4_56[19], stage4_56[20], stage4_56[21], stage4_56[22], stage4_56[23]},
      {stage5_58[3],stage5_57[4],stage5_56[5],stage5_55[8],stage5_54[11]}
   );
   gpc606_5 gpc10539 (
      {stage4_55[10], stage4_55[11], stage4_55[12], stage4_55[13], stage4_55[14], stage4_55[15]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage5_59[0],stage5_58[4],stage5_57[5],stage5_56[6],stage5_55[9]}
   );
   gpc606_5 gpc10540 (
      {stage4_55[16], stage4_55[17], stage4_55[18], stage4_55[19], stage4_55[20], stage4_55[21]},
      {stage4_57[6], stage4_57[7], stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11]},
      {stage5_59[1],stage5_58[5],stage5_57[6],stage5_56[7],stage5_55[10]}
   );
   gpc207_4 gpc10541 (
      {stage4_57[12], stage4_57[13], stage4_57[14], stage4_57[15], stage4_57[16], stage4_57[17], stage4_57[18]},
      {stage4_59[0], stage4_59[1]},
      {stage5_60[0],stage5_59[2],stage5_58[6],stage5_57[7]}
   );
   gpc207_4 gpc10542 (
      {stage4_57[19], stage4_57[20], stage4_57[21], stage4_57[22], stage4_57[23], stage4_57[24], 1'b0},
      {stage4_59[2], stage4_59[3]},
      {stage5_60[1],stage5_59[3],stage5_58[7],stage5_57[8]}
   );
   gpc606_5 gpc10543 (
      {stage4_59[4], stage4_59[5], stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[2],stage5_59[4]}
   );
   gpc606_5 gpc10544 (
      {stage4_59[10], stage4_59[11], stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[3],stage5_59[5]}
   );
   gpc606_5 gpc10545 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[2],stage5_61[2],stage5_60[4]}
   );
   gpc606_5 gpc10546 (
      {stage4_60[6], stage4_60[7], stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11]},
      {stage4_62[6], stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage5_64[1],stage5_63[3],stage5_62[3],stage5_61[3],stage5_60[5]}
   );
   gpc606_5 gpc10547 (
      {stage4_60[12], stage4_60[13], stage4_60[14], stage4_60[15], stage4_60[16], stage4_60[17]},
      {stage4_62[12], stage4_62[13], stage4_62[14], stage4_62[15], stage4_62[16], stage4_62[17]},
      {stage5_64[2],stage5_63[4],stage5_62[4],stage5_61[4],stage5_60[6]}
   );
   gpc7_3 gpc10548 (
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17], stage4_61[18]},
      {stage5_63[5],stage5_62[5],stage5_61[5]}
   );
   gpc7_3 gpc10549 (
      {stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22], stage4_61[23], stage4_61[24], stage4_61[25]},
      {stage5_63[6],stage5_62[6],stage5_61[6]}
   );
   gpc606_5 gpc10550 (
      {stage4_62[18], stage4_62[19], stage4_62[20], stage4_62[21], stage4_62[22], stage4_62[23]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[0],stage5_64[3],stage5_63[7],stage5_62[7]}
   );
   gpc606_5 gpc10551 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[4],stage5_63[8]}
   );
   gpc606_5 gpc10552 (
      {stage4_63[6], stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8], stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[5],stage5_63[9]}
   );
   gpc606_5 gpc10553 (
      {stage4_63[12], stage4_63[13], stage4_63[14], stage4_63[15], stage4_63[16], stage4_63[17]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage5_67[2],stage5_66[3],stage5_65[3],stage5_64[6],stage5_63[10]}
   );
   gpc135_4 gpc10554 (
      {stage4_64[6], stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10]},
      {stage4_65[18], stage4_65[19], stage4_65[20]},
      {stage4_66[0]},
      {stage5_67[3],stage5_66[4],stage5_65[4],stage5_64[7]}
   );
   gpc135_4 gpc10555 (
      {stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15]},
      {stage4_65[21], stage4_65[22], 1'b0},
      {stage4_66[1]},
      {stage5_67[4],stage5_66[5],stage5_65[5],stage5_64[8]}
   );
   gpc1163_5 gpc10556 (
      {stage4_66[2], stage4_66[3], stage4_66[4]},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage4_68[0]},
      {stage4_69[0]},
      {stage5_70[0],stage5_69[0],stage5_68[0],stage5_67[5],stage5_66[6]}
   );
   gpc1163_5 gpc10557 (
      {stage4_66[5], stage4_66[6], stage4_66[7]},
      {stage4_67[6], stage4_67[7], stage4_67[8], stage4_67[9], stage4_67[10], stage4_67[11]},
      {stage4_68[1]},
      {stage4_69[1]},
      {stage5_70[1],stage5_69[1],stage5_68[1],stage5_67[6],stage5_66[7]}
   );
   gpc1163_5 gpc10558 (
      {stage4_66[8], stage4_66[9], stage4_66[10]},
      {stage4_67[12], stage4_67[13], stage4_67[14], stage4_67[15], stage4_67[16], 1'b0},
      {stage4_68[2]},
      {stage4_69[2]},
      {stage5_70[2],stage5_69[2],stage5_68[2],stage5_67[7],stage5_66[8]}
   );
   gpc1_1 gpc10559 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc10560 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc10561 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc10562 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc10563 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc10564 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc10565 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc10566 (
      {stage4_3[18]},
      {stage5_3[4]}
   );
   gpc1_1 gpc10567 (
      {stage4_3[19]},
      {stage5_3[5]}
   );
   gpc1_1 gpc10568 (
      {stage4_3[20]},
      {stage5_3[6]}
   );
   gpc1_1 gpc10569 (
      {stage4_3[21]},
      {stage5_3[7]}
   );
   gpc1_1 gpc10570 (
      {stage4_4[23]},
      {stage5_4[7]}
   );
   gpc1_1 gpc10571 (
      {stage4_4[24]},
      {stage5_4[8]}
   );
   gpc1_1 gpc10572 (
      {stage4_5[38]},
      {stage5_5[12]}
   );
   gpc1_1 gpc10573 (
      {stage4_5[39]},
      {stage5_5[13]}
   );
   gpc1_1 gpc10574 (
      {stage4_5[40]},
      {stage5_5[14]}
   );
   gpc1_1 gpc10575 (
      {stage4_5[41]},
      {stage5_5[15]}
   );
   gpc1_1 gpc10576 (
      {stage4_5[42]},
      {stage5_5[16]}
   );
   gpc1_1 gpc10577 (
      {stage4_5[43]},
      {stage5_5[17]}
   );
   gpc1_1 gpc10578 (
      {stage4_5[44]},
      {stage5_5[18]}
   );
   gpc1_1 gpc10579 (
      {stage4_5[45]},
      {stage5_5[19]}
   );
   gpc1_1 gpc10580 (
      {stage4_5[46]},
      {stage5_5[20]}
   );
   gpc1_1 gpc10581 (
      {stage4_6[18]},
      {stage5_6[11]}
   );
   gpc1_1 gpc10582 (
      {stage4_6[19]},
      {stage5_6[12]}
   );
   gpc1_1 gpc10583 (
      {stage4_6[20]},
      {stage5_6[13]}
   );
   gpc1_1 gpc10584 (
      {stage4_11[28]},
      {stage5_11[14]}
   );
   gpc1_1 gpc10585 (
      {stage4_11[29]},
      {stage5_11[15]}
   );
   gpc1_1 gpc10586 (
      {stage4_11[30]},
      {stage5_11[16]}
   );
   gpc1_1 gpc10587 (
      {stage4_11[31]},
      {stage5_11[17]}
   );
   gpc1_1 gpc10588 (
      {stage4_11[32]},
      {stage5_11[18]}
   );
   gpc1_1 gpc10589 (
      {stage4_11[33]},
      {stage5_11[19]}
   );
   gpc1_1 gpc10590 (
      {stage4_12[16]},
      {stage5_12[10]}
   );
   gpc1_1 gpc10591 (
      {stage4_12[17]},
      {stage5_12[11]}
   );
   gpc1_1 gpc10592 (
      {stage4_12[18]},
      {stage5_12[12]}
   );
   gpc1_1 gpc10593 (
      {stage4_12[19]},
      {stage5_12[13]}
   );
   gpc1_1 gpc10594 (
      {stage4_13[26]},
      {stage5_13[7]}
   );
   gpc1_1 gpc10595 (
      {stage4_13[27]},
      {stage5_13[8]}
   );
   gpc1_1 gpc10596 (
      {stage4_14[26]},
      {stage5_14[11]}
   );
   gpc1_1 gpc10597 (
      {stage4_14[27]},
      {stage5_14[12]}
   );
   gpc1_1 gpc10598 (
      {stage4_14[28]},
      {stage5_14[13]}
   );
   gpc1_1 gpc10599 (
      {stage4_14[29]},
      {stage5_14[14]}
   );
   gpc1_1 gpc10600 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc10601 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc10602 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc10603 (
      {stage4_15[22]},
      {stage5_15[15]}
   );
   gpc1_1 gpc10604 (
      {stage4_16[27]},
      {stage5_16[8]}
   );
   gpc1_1 gpc10605 (
      {stage4_16[28]},
      {stage5_16[9]}
   );
   gpc1_1 gpc10606 (
      {stage4_16[29]},
      {stage5_16[10]}
   );
   gpc1_1 gpc10607 (
      {stage4_16[30]},
      {stage5_16[11]}
   );
   gpc1_1 gpc10608 (
      {stage4_16[31]},
      {stage5_16[12]}
   );
   gpc1_1 gpc10609 (
      {stage4_16[32]},
      {stage5_16[13]}
   );
   gpc1_1 gpc10610 (
      {stage4_19[17]},
      {stage5_19[11]}
   );
   gpc1_1 gpc10611 (
      {stage4_19[18]},
      {stage5_19[12]}
   );
   gpc1_1 gpc10612 (
      {stage4_19[19]},
      {stage5_19[13]}
   );
   gpc1_1 gpc10613 (
      {stage4_21[26]},
      {stage5_21[10]}
   );
   gpc1_1 gpc10614 (
      {stage4_23[21]},
      {stage5_23[9]}
   );
   gpc1_1 gpc10615 (
      {stage4_23[22]},
      {stage5_23[10]}
   );
   gpc1_1 gpc10616 (
      {stage4_23[23]},
      {stage5_23[11]}
   );
   gpc1_1 gpc10617 (
      {stage4_24[21]},
      {stage5_24[6]}
   );
   gpc1_1 gpc10618 (
      {stage4_24[22]},
      {stage5_24[7]}
   );
   gpc1_1 gpc10619 (
      {stage4_24[23]},
      {stage5_24[8]}
   );
   gpc1_1 gpc10620 (
      {stage4_25[15]},
      {stage5_25[8]}
   );
   gpc1_1 gpc10621 (
      {stage4_25[16]},
      {stage5_25[9]}
   );
   gpc1_1 gpc10622 (
      {stage4_25[17]},
      {stage5_25[10]}
   );
   gpc1_1 gpc10623 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc10624 (
      {stage4_25[19]},
      {stage5_25[12]}
   );
   gpc1_1 gpc10625 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc10626 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc10627 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc10628 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc10629 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc10630 (
      {stage4_26[19]},
      {stage5_26[15]}
   );
   gpc1_1 gpc10631 (
      {stage4_26[20]},
      {stage5_26[16]}
   );
   gpc1_1 gpc10632 (
      {stage4_27[17]},
      {stage5_27[5]}
   );
   gpc1_1 gpc10633 (
      {stage4_27[18]},
      {stage5_27[6]}
   );
   gpc1_1 gpc10634 (
      {stage4_27[19]},
      {stage5_27[7]}
   );
   gpc1_1 gpc10635 (
      {stage4_27[20]},
      {stage5_27[8]}
   );
   gpc1_1 gpc10636 (
      {stage4_28[29]},
      {stage5_28[9]}
   );
   gpc1_1 gpc10637 (
      {stage4_28[30]},
      {stage5_28[10]}
   );
   gpc1_1 gpc10638 (
      {stage4_28[31]},
      {stage5_28[11]}
   );
   gpc1_1 gpc10639 (
      {stage4_29[20]},
      {stage5_29[11]}
   );
   gpc1_1 gpc10640 (
      {stage4_29[21]},
      {stage5_29[12]}
   );
   gpc1_1 gpc10641 (
      {stage4_29[22]},
      {stage5_29[13]}
   );
   gpc1_1 gpc10642 (
      {stage4_29[23]},
      {stage5_29[14]}
   );
   gpc1_1 gpc10643 (
      {stage4_30[24]},
      {stage5_30[7]}
   );
   gpc1_1 gpc10644 (
      {stage4_30[25]},
      {stage5_30[8]}
   );
   gpc1_1 gpc10645 (
      {stage4_31[14]},
      {stage5_31[9]}
   );
   gpc1_1 gpc10646 (
      {stage4_31[15]},
      {stage5_31[10]}
   );
   gpc1_1 gpc10647 (
      {stage4_31[16]},
      {stage5_31[11]}
   );
   gpc1_1 gpc10648 (
      {stage4_32[20]},
      {stage5_32[11]}
   );
   gpc1_1 gpc10649 (
      {stage4_32[21]},
      {stage5_32[12]}
   );
   gpc1_1 gpc10650 (
      {stage4_32[22]},
      {stage5_32[13]}
   );
   gpc1_1 gpc10651 (
      {stage4_32[23]},
      {stage5_32[14]}
   );
   gpc1_1 gpc10652 (
      {stage4_34[18]},
      {stage5_34[9]}
   );
   gpc1_1 gpc10653 (
      {stage4_34[19]},
      {stage5_34[10]}
   );
   gpc1_1 gpc10654 (
      {stage4_34[20]},
      {stage5_34[11]}
   );
   gpc1_1 gpc10655 (
      {stage4_34[21]},
      {stage5_34[12]}
   );
   gpc1_1 gpc10656 (
      {stage4_34[22]},
      {stage5_34[13]}
   );
   gpc1_1 gpc10657 (
      {stage4_34[23]},
      {stage5_34[14]}
   );
   gpc1_1 gpc10658 (
      {stage4_34[24]},
      {stage5_34[15]}
   );
   gpc1_1 gpc10659 (
      {stage4_34[25]},
      {stage5_34[16]}
   );
   gpc1_1 gpc10660 (
      {stage4_34[26]},
      {stage5_34[17]}
   );
   gpc1_1 gpc10661 (
      {stage4_34[27]},
      {stage5_34[18]}
   );
   gpc1_1 gpc10662 (
      {stage4_34[28]},
      {stage5_34[19]}
   );
   gpc1_1 gpc10663 (
      {stage4_34[29]},
      {stage5_34[20]}
   );
   gpc1_1 gpc10664 (
      {stage4_36[33]},
      {stage5_36[14]}
   );
   gpc1_1 gpc10665 (
      {stage4_36[34]},
      {stage5_36[15]}
   );
   gpc1_1 gpc10666 (
      {stage4_36[35]},
      {stage5_36[16]}
   );
   gpc1_1 gpc10667 (
      {stage4_36[36]},
      {stage5_36[17]}
   );
   gpc1_1 gpc10668 (
      {stage4_36[37]},
      {stage5_36[18]}
   );
   gpc1_1 gpc10669 (
      {stage4_40[22]},
      {stage5_40[13]}
   );
   gpc1_1 gpc10670 (
      {stage4_40[23]},
      {stage5_40[14]}
   );
   gpc1_1 gpc10671 (
      {stage4_40[24]},
      {stage5_40[15]}
   );
   gpc1_1 gpc10672 (
      {stage4_40[25]},
      {stage5_40[16]}
   );
   gpc1_1 gpc10673 (
      {stage4_40[26]},
      {stage5_40[17]}
   );
   gpc1_1 gpc10674 (
      {stage4_40[27]},
      {stage5_40[18]}
   );
   gpc1_1 gpc10675 (
      {stage4_40[28]},
      {stage5_40[19]}
   );
   gpc1_1 gpc10676 (
      {stage4_42[19]},
      {stage5_42[10]}
   );
   gpc1_1 gpc10677 (
      {stage4_42[20]},
      {stage5_42[11]}
   );
   gpc1_1 gpc10678 (
      {stage4_42[21]},
      {stage5_42[12]}
   );
   gpc1_1 gpc10679 (
      {stage4_42[22]},
      {stage5_42[13]}
   );
   gpc1_1 gpc10680 (
      {stage4_42[23]},
      {stage5_42[14]}
   );
   gpc1_1 gpc10681 (
      {stage4_42[24]},
      {stage5_42[15]}
   );
   gpc1_1 gpc10682 (
      {stage4_42[25]},
      {stage5_42[16]}
   );
   gpc1_1 gpc10683 (
      {stage4_42[26]},
      {stage5_42[17]}
   );
   gpc1_1 gpc10684 (
      {stage4_42[27]},
      {stage5_42[18]}
   );
   gpc1_1 gpc10685 (
      {stage4_42[28]},
      {stage5_42[19]}
   );
   gpc1_1 gpc10686 (
      {stage4_44[26]},
      {stage5_44[12]}
   );
   gpc1_1 gpc10687 (
      {stage4_44[27]},
      {stage5_44[13]}
   );
   gpc1_1 gpc10688 (
      {stage4_44[28]},
      {stage5_44[14]}
   );
   gpc1_1 gpc10689 (
      {stage4_44[29]},
      {stage5_44[15]}
   );
   gpc1_1 gpc10690 (
      {stage4_44[30]},
      {stage5_44[16]}
   );
   gpc1_1 gpc10691 (
      {stage4_44[31]},
      {stage5_44[17]}
   );
   gpc1_1 gpc10692 (
      {stage4_44[32]},
      {stage5_44[18]}
   );
   gpc1_1 gpc10693 (
      {stage4_44[33]},
      {stage5_44[19]}
   );
   gpc1_1 gpc10694 (
      {stage4_44[34]},
      {stage5_44[20]}
   );
   gpc1_1 gpc10695 (
      {stage4_44[35]},
      {stage5_44[21]}
   );
   gpc1_1 gpc10696 (
      {stage4_44[36]},
      {stage5_44[22]}
   );
   gpc1_1 gpc10697 (
      {stage4_44[37]},
      {stage5_44[23]}
   );
   gpc1_1 gpc10698 (
      {stage4_44[38]},
      {stage5_44[24]}
   );
   gpc1_1 gpc10699 (
      {stage4_44[39]},
      {stage5_44[25]}
   );
   gpc1_1 gpc10700 (
      {stage4_48[11]},
      {stage5_48[7]}
   );
   gpc1_1 gpc10701 (
      {stage4_48[12]},
      {stage5_48[8]}
   );
   gpc1_1 gpc10702 (
      {stage4_48[13]},
      {stage5_48[9]}
   );
   gpc1_1 gpc10703 (
      {stage4_48[14]},
      {stage5_48[10]}
   );
   gpc1_1 gpc10704 (
      {stage4_48[15]},
      {stage5_48[11]}
   );
   gpc1_1 gpc10705 (
      {stage4_48[16]},
      {stage5_48[12]}
   );
   gpc1_1 gpc10706 (
      {stage4_48[17]},
      {stage5_48[13]}
   );
   gpc1_1 gpc10707 (
      {stage4_48[18]},
      {stage5_48[14]}
   );
   gpc1_1 gpc10708 (
      {stage4_48[19]},
      {stage5_48[15]}
   );
   gpc1_1 gpc10709 (
      {stage4_48[20]},
      {stage5_48[16]}
   );
   gpc1_1 gpc10710 (
      {stage4_48[21]},
      {stage5_48[17]}
   );
   gpc1_1 gpc10711 (
      {stage4_49[18]},
      {stage5_49[7]}
   );
   gpc1_1 gpc10712 (
      {stage4_49[19]},
      {stage5_49[8]}
   );
   gpc1_1 gpc10713 (
      {stage4_49[20]},
      {stage5_49[9]}
   );
   gpc1_1 gpc10714 (
      {stage4_49[21]},
      {stage5_49[10]}
   );
   gpc1_1 gpc10715 (
      {stage4_49[22]},
      {stage5_49[11]}
   );
   gpc1_1 gpc10716 (
      {stage4_49[23]},
      {stage5_49[12]}
   );
   gpc1_1 gpc10717 (
      {stage4_49[24]},
      {stage5_49[13]}
   );
   gpc1_1 gpc10718 (
      {stage4_49[25]},
      {stage5_49[14]}
   );
   gpc1_1 gpc10719 (
      {stage4_49[26]},
      {stage5_49[15]}
   );
   gpc1_1 gpc10720 (
      {stage4_49[27]},
      {stage5_49[16]}
   );
   gpc1_1 gpc10721 (
      {stage4_52[19]},
      {stage5_52[9]}
   );
   gpc1_1 gpc10722 (
      {stage4_52[20]},
      {stage5_52[10]}
   );
   gpc1_1 gpc10723 (
      {stage4_52[21]},
      {stage5_52[11]}
   );
   gpc1_1 gpc10724 (
      {stage4_52[22]},
      {stage5_52[12]}
   );
   gpc1_1 gpc10725 (
      {stage4_53[25]},
      {stage5_53[8]}
   );
   gpc1_1 gpc10726 (
      {stage4_53[26]},
      {stage5_53[9]}
   );
   gpc1_1 gpc10727 (
      {stage4_53[27]},
      {stage5_53[10]}
   );
   gpc1_1 gpc10728 (
      {stage4_53[28]},
      {stage5_53[11]}
   );
   gpc1_1 gpc10729 (
      {stage4_54[26]},
      {stage5_54[12]}
   );
   gpc1_1 gpc10730 (
      {stage4_54[27]},
      {stage5_54[13]}
   );
   gpc1_1 gpc10731 (
      {stage4_54[28]},
      {stage5_54[14]}
   );
   gpc1_1 gpc10732 (
      {stage4_54[29]},
      {stage5_54[15]}
   );
   gpc1_1 gpc10733 (
      {stage4_54[30]},
      {stage5_54[16]}
   );
   gpc1_1 gpc10734 (
      {stage4_55[22]},
      {stage5_55[11]}
   );
   gpc1_1 gpc10735 (
      {stage4_55[23]},
      {stage5_55[12]}
   );
   gpc1_1 gpc10736 (
      {stage4_55[24]},
      {stage5_55[13]}
   );
   gpc1_1 gpc10737 (
      {stage4_55[25]},
      {stage5_55[14]}
   );
   gpc1_1 gpc10738 (
      {stage4_55[26]},
      {stage5_55[15]}
   );
   gpc1_1 gpc10739 (
      {stage4_55[27]},
      {stage5_55[16]}
   );
   gpc1_1 gpc10740 (
      {stage4_55[28]},
      {stage5_55[17]}
   );
   gpc1_1 gpc10741 (
      {stage4_56[24]},
      {stage5_56[8]}
   );
   gpc1_1 gpc10742 (
      {stage4_56[25]},
      {stage5_56[9]}
   );
   gpc1_1 gpc10743 (
      {stage4_56[26]},
      {stage5_56[10]}
   );
   gpc1_1 gpc10744 (
      {stage4_56[27]},
      {stage5_56[11]}
   );
   gpc1_1 gpc10745 (
      {stage4_56[28]},
      {stage5_56[12]}
   );
   gpc1_1 gpc10746 (
      {stage4_58[0]},
      {stage5_58[8]}
   );
   gpc1_1 gpc10747 (
      {stage4_58[1]},
      {stage5_58[9]}
   );
   gpc1_1 gpc10748 (
      {stage4_58[2]},
      {stage5_58[10]}
   );
   gpc1_1 gpc10749 (
      {stage4_58[3]},
      {stage5_58[11]}
   );
   gpc1_1 gpc10750 (
      {stage4_58[4]},
      {stage5_58[12]}
   );
   gpc1_1 gpc10751 (
      {stage4_58[5]},
      {stage5_58[13]}
   );
   gpc1_1 gpc10752 (
      {stage4_58[6]},
      {stage5_58[14]}
   );
   gpc1_1 gpc10753 (
      {stage4_58[7]},
      {stage5_58[15]}
   );
   gpc1_1 gpc10754 (
      {stage4_58[8]},
      {stage5_58[16]}
   );
   gpc1_1 gpc10755 (
      {stage4_58[9]},
      {stage5_58[17]}
   );
   gpc1_1 gpc10756 (
      {stage4_58[10]},
      {stage5_58[18]}
   );
   gpc1_1 gpc10757 (
      {stage4_58[11]},
      {stage5_58[19]}
   );
   gpc1_1 gpc10758 (
      {stage4_58[12]},
      {stage5_58[20]}
   );
   gpc1_1 gpc10759 (
      {stage4_58[13]},
      {stage5_58[21]}
   );
   gpc1_1 gpc10760 (
      {stage4_58[14]},
      {stage5_58[22]}
   );
   gpc1_1 gpc10761 (
      {stage4_58[15]},
      {stage5_58[23]}
   );
   gpc1_1 gpc10762 (
      {stage4_60[18]},
      {stage5_60[7]}
   );
   gpc1_1 gpc10763 (
      {stage4_60[19]},
      {stage5_60[8]}
   );
   gpc1_1 gpc10764 (
      {stage4_60[20]},
      {stage5_60[9]}
   );
   gpc1_1 gpc10765 (
      {stage4_60[21]},
      {stage5_60[10]}
   );
   gpc1_1 gpc10766 (
      {stage4_60[22]},
      {stage5_60[11]}
   );
   gpc1_1 gpc10767 (
      {stage4_60[23]},
      {stage5_60[12]}
   );
   gpc1_1 gpc10768 (
      {stage4_60[24]},
      {stage5_60[13]}
   );
   gpc1_1 gpc10769 (
      {stage4_61[26]},
      {stage5_61[7]}
   );
   gpc1_1 gpc10770 (
      {stage4_61[27]},
      {stage5_61[8]}
   );
   gpc1_1 gpc10771 (
      {stage4_61[28]},
      {stage5_61[9]}
   );
   gpc1_1 gpc10772 (
      {stage4_64[16]},
      {stage5_64[9]}
   );
   gpc1_1 gpc10773 (
      {stage4_64[17]},
      {stage5_64[10]}
   );
   gpc1_1 gpc10774 (
      {stage4_64[18]},
      {stage5_64[11]}
   );
   gpc1_1 gpc10775 (
      {stage4_64[19]},
      {stage5_64[12]}
   );
   gpc1_1 gpc10776 (
      {stage4_64[20]},
      {stage5_64[13]}
   );
   gpc1_1 gpc10777 (
      {stage4_64[21]},
      {stage5_64[14]}
   );
   gpc1_1 gpc10778 (
      {stage4_64[22]},
      {stage5_64[15]}
   );
   gpc1_1 gpc10779 (
      {stage4_64[23]},
      {stage5_64[16]}
   );
   gpc1_1 gpc10780 (
      {stage4_64[24]},
      {stage5_64[17]}
   );
   gpc1_1 gpc10781 (
      {stage4_64[25]},
      {stage5_64[18]}
   );
   gpc1_1 gpc10782 (
      {stage4_64[26]},
      {stage5_64[19]}
   );
   gpc1_1 gpc10783 (
      {stage4_66[11]},
      {stage5_66[9]}
   );
   gpc1_1 gpc10784 (
      {stage4_66[12]},
      {stage5_66[10]}
   );
   gpc1_1 gpc10785 (
      {stage4_66[13]},
      {stage5_66[11]}
   );
   gpc1_1 gpc10786 (
      {stage4_66[14]},
      {stage5_66[12]}
   );
   gpc1_1 gpc10787 (
      {stage4_68[3]},
      {stage5_68[3]}
   );
   gpc1_1 gpc10788 (
      {stage4_68[4]},
      {stage5_68[4]}
   );
   gpc1_1 gpc10789 (
      {stage4_68[5]},
      {stage5_68[5]}
   );
   gpc1_1 gpc10790 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc10791 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc10792 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc10793 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc10794 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc10795 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc10796 (
      {stage4_70[0]},
      {stage5_70[3]}
   );
   gpc615_5 gpc10797 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc207_4 gpc10798 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc10799 (
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc606_5 gpc10800 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], stage5_5[16], stage5_5[17]},
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10], 1'b0},
      {stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc117_4 gpc10801 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {1'b0},
      {stage5_8[0]},
      {stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[4]}
   );
   gpc615_5 gpc10802 (
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12], stage5_6[13]},
      {1'b0},
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[5],stage6_6[5]}
   );
   gpc606_5 gpc10803 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[4],stage6_8[4]}
   );
   gpc606_5 gpc10804 (
      {stage5_8[13], stage5_8[14], stage5_8[15], 1'b0, 1'b0, 1'b0},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], 1'b0, 1'b0},
      {stage6_12[1],stage6_11[1],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc207_4 gpc10805 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5], stage5_9[6]},
      {stage5_11[0], stage5_11[1]},
      {stage6_12[2],stage6_11[2],stage6_10[3],stage6_9[6]}
   );
   gpc606_5 gpc10806 (
      {stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11], stage5_9[12]},
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7]},
      {stage6_13[0],stage6_12[3],stage6_11[3],stage6_10[4],stage6_9[7]}
   );
   gpc1406_5 gpc10807 (
      {stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[4],stage6_11[4]}
   );
   gpc1406_5 gpc10808 (
      {stage5_11[14], stage5_11[15], stage5_11[16], stage5_11[17], stage5_11[18], stage5_11[19]},
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7]},
      {stage5_14[1]},
      {stage6_15[1],stage6_14[1],stage6_13[2],stage6_12[5],stage6_11[5]}
   );
   gpc117_4 gpc10809 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage5_13[8]},
      {stage5_14[2]},
      {stage6_15[2],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc117_4 gpc10810 (
      {stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {1'b0},
      {stage5_14[3]},
      {stage6_15[3],stage6_14[3],stage6_13[4],stage6_12[7]}
   );
   gpc1343_5 gpc10811 (
      {stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[4],stage6_14[4]}
   );
   gpc1343_5 gpc10812 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[5],stage6_14[5]}
   );
   gpc1343_5 gpc10813 (
      {stage5_14[10], stage5_14[11], stage5_14[12]},
      {stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage5_16[6], stage5_16[7], stage5_16[8]},
      {stage5_17[2]},
      {stage6_18[2],stage6_17[2],stage6_16[2],stage6_15[6],stage6_14[6]}
   );
   gpc1343_5 gpc10814 (
      {stage5_14[13], stage5_14[14], 1'b0},
      {stage5_15[12], stage5_15[13], stage5_15[14], stage5_15[15]},
      {stage5_16[9], stage5_16[10], stage5_16[11]},
      {stage5_17[3]},
      {stage6_18[3],stage6_17[3],stage6_16[3],stage6_15[7],stage6_14[7]}
   );
   gpc207_4 gpc10815 (
      {stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7], 1'b0, 1'b0, 1'b0},
      {stage5_19[0], stage5_19[1]},
      {stage6_20[0],stage6_19[0],stage6_18[4],stage6_17[4]}
   );
   gpc7_3 gpc10816 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage6_20[1],stage6_19[1],stage6_18[5]}
   );
   gpc7_3 gpc10817 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13]},
      {stage6_20[2],stage6_19[2],stage6_18[6]}
   );
   gpc2135_5 gpc10818 (
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[3],stage6_19[3]}
   );
   gpc7_3 gpc10819 (
      {stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13]},
      {stage6_21[1],stage6_20[4],stage6_19[4]}
   );
   gpc1415_5 gpc10820 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_21[1]},
      {stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[2],stage6_20[5]}
   );
   gpc207_4 gpc10821 (
      {stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5], stage5_21[6], stage5_21[7], stage5_21[8]},
      {stage5_23[1], stage5_23[2]},
      {stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[3]}
   );
   gpc606_5 gpc10822 (
      {stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[3]}
   );
   gpc606_5 gpc10823 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3]}
   );
   gpc1343_5 gpc10824 (
      {stage5_26[6], stage5_26[7], stage5_26[8]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[2],stage6_26[2]}
   );
   gpc1343_5 gpc10825 (
      {stage5_26[9], stage5_26[10], stage5_26[11]},
      {stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage5_29[1]},
      {stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc10826 (
      {stage5_26[12], stage5_26[13], stage5_26[14], stage5_26[15], stage5_26[16]},
      {stage5_27[8]},
      {stage5_28[6], stage5_28[7], stage5_28[8], stage5_28[9], stage5_28[10], stage5_28[11]},
      {stage6_30[2],stage6_29[2],stage6_28[3],stage6_27[4],stage6_26[4]}
   );
   gpc606_5 gpc10827 (
      {stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6], stage5_29[7]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[3],stage6_29[3]}
   );
   gpc606_5 gpc10828 (
      {stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11], stage5_29[12], stage5_29[13]},
      {stage5_31[6], stage5_31[7], stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11]},
      {stage6_33[1],stage6_32[1],stage6_31[1],stage6_30[4],stage6_29[4]}
   );
   gpc7_3 gpc10829 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage6_32[2],stage6_31[2],stage6_30[5]}
   );
   gpc1415_5 gpc10830 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4]},
      {stage5_33[0]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3]},
      {stage5_35[0]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[2],stage6_32[3]}
   );
   gpc1415_5 gpc10831 (
      {stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage5_33[1]},
      {stage5_34[4], stage5_34[5], stage5_34[6], stage5_34[7]},
      {stage5_35[1]},
      {stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[3],stage6_32[4]}
   );
   gpc606_5 gpc10832 (
      {stage5_32[10], stage5_32[11], stage5_32[12], stage5_32[13], stage5_32[14], 1'b0},
      {stage5_34[8], stage5_34[9], stage5_34[10], stage5_34[11], stage5_34[12], stage5_34[13]},
      {stage6_36[2],stage6_35[2],stage6_34[2],stage6_33[4],stage6_32[5]}
   );
   gpc615_5 gpc10833 (
      {stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_34[14]},
      {stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5], stage5_35[6], stage5_35[7]},
      {stage6_37[0],stage6_36[3],stage6_35[3],stage6_34[3],stage6_33[5]}
   );
   gpc615_5 gpc10834 (
      {stage5_34[15], stage5_34[16], stage5_34[17], stage5_34[18], stage5_34[19]},
      {stage5_35[8]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[4],stage6_35[4],stage6_34[4]}
   );
   gpc2135_5 gpc10835 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10]},
      {stage5_37[0], stage5_37[1], stage5_37[2]},
      {stage5_38[0]},
      {stage5_39[0], stage5_39[1]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[2],stage6_36[5]}
   );
   gpc2135_5 gpc10836 (
      {stage5_36[11], stage5_36[12], stage5_36[13], stage5_36[14], stage5_36[15]},
      {stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage5_38[1]},
      {stage5_39[2], stage5_39[3]},
      {stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[3],stage6_36[6]}
   );
   gpc606_5 gpc10837 (
      {stage5_36[16], stage5_36[17], stage5_36[18], 1'b0, 1'b0, 1'b0},
      {stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5], stage5_38[6], 1'b0},
      {stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[4],stage6_36[7]}
   );
   gpc606_5 gpc10838 (
      {stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10], 1'b0},
      {stage5_39[4], stage5_39[5], stage5_39[6], stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage6_41[0],stage6_40[3],stage6_39[3],stage6_38[4],stage6_37[5]}
   );
   gpc606_5 gpc10839 (
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[1],stage6_40[4]}
   );
   gpc606_5 gpc10840 (
      {stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9], stage5_40[10], stage5_40[11]},
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10], stage5_42[11]},
      {stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[2],stage6_40[5]}
   );
   gpc1325_5 gpc10841 (
      {stage5_40[12], stage5_40[13], stage5_40[14], stage5_40[15], stage5_40[16]},
      {stage5_41[0], stage5_41[1]},
      {stage5_42[12], stage5_42[13], stage5_42[14]},
      {stage5_43[0]},
      {stage6_44[2],stage6_43[2],stage6_42[2],stage6_41[3],stage6_40[6]}
   );
   gpc615_5 gpc10842 (
      {stage5_42[15], stage5_42[16], stage5_42[17], stage5_42[18], stage5_42[19]},
      {stage5_43[1]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[0],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc7_3 gpc10843 (
      {stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5], stage5_43[6], stage5_43[7], 1'b0},
      {stage6_45[1],stage6_44[4],stage6_43[4]}
   );
   gpc7_3 gpc10844 (
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11], stage5_44[12]},
      {stage6_46[1],stage6_45[2],stage6_44[5]}
   );
   gpc7_3 gpc10845 (
      {stage5_44[13], stage5_44[14], stage5_44[15], stage5_44[16], stage5_44[17], stage5_44[18], stage5_44[19]},
      {stage6_46[2],stage6_45[3],stage6_44[6]}
   );
   gpc606_5 gpc10846 (
      {stage5_44[20], stage5_44[21], stage5_44[22], stage5_44[23], stage5_44[24], stage5_44[25]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[3],stage6_45[4],stage6_44[7]}
   );
   gpc606_5 gpc10847 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc10848 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], 1'b0, 1'b0},
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10], stage5_47[11]},
      {stage6_49[1],stage6_48[2],stage6_47[2],stage6_46[5],stage6_45[6]}
   );
   gpc615_5 gpc10849 (
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10]},
      {stage5_47[12]},
      {stage5_48[0], stage5_48[1], stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5]},
      {stage6_50[0],stage6_49[2],stage6_48[3],stage6_47[3],stage6_46[6]}
   );
   gpc606_5 gpc10850 (
      {stage5_48[6], stage5_48[7], stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[1],stage6_49[3],stage6_48[4]}
   );
   gpc606_5 gpc10851 (
      {stage5_48[12], stage5_48[13], stage5_48[14], stage5_48[15], stage5_48[16], stage5_48[17]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], 1'b0, 1'b0},
      {stage6_52[1],stage6_51[1],stage6_50[2],stage6_49[4],stage6_48[5]}
   );
   gpc207_4 gpc10852 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5], stage5_49[6]},
      {stage5_51[0], stage5_51[1]},
      {stage6_52[2],stage6_51[2],stage6_50[3],stage6_49[5]}
   );
   gpc207_4 gpc10853 (
      {stage5_49[7], stage5_49[8], stage5_49[9], stage5_49[10], stage5_49[11], stage5_49[12], stage5_49[13]},
      {stage5_51[2], stage5_51[3]},
      {stage6_52[3],stage6_51[3],stage6_50[4],stage6_49[6]}
   );
   gpc606_5 gpc10854 (
      {stage5_51[4], stage5_51[5], stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[0],stage6_52[4],stage6_51[4]}
   );
   gpc606_5 gpc10855 (
      {stage5_52[0], stage5_52[1], stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5]},
      {stage5_54[0], stage5_54[1], stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5]},
      {stage6_56[0],stage6_55[1],stage6_54[1],stage6_53[1],stage6_52[5]}
   );
   gpc606_5 gpc10856 (
      {stage5_52[6], stage5_52[7], stage5_52[8], stage5_52[9], stage5_52[10], stage5_52[11]},
      {stage5_54[6], stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage6_56[1],stage6_55[2],stage6_54[2],stage6_53[2],stage6_52[6]}
   );
   gpc606_5 gpc10857 (
      {stage5_53[6], stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11]},
      {stage5_55[0], stage5_55[1], stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5]},
      {stage6_57[0],stage6_56[2],stage6_55[3],stage6_54[3],stage6_53[3]}
   );
   gpc1163_5 gpc10858 (
      {stage5_54[12], stage5_54[13], stage5_54[14]},
      {stage5_55[6], stage5_55[7], stage5_55[8], stage5_55[9], stage5_55[10], stage5_55[11]},
      {stage5_56[0]},
      {stage5_57[0]},
      {stage6_58[0],stage6_57[1],stage6_56[3],stage6_55[4],stage6_54[4]}
   );
   gpc1163_5 gpc10859 (
      {stage5_54[15], stage5_54[16], 1'b0},
      {stage5_55[12], stage5_55[13], stage5_55[14], stage5_55[15], stage5_55[16], stage5_55[17]},
      {stage5_56[1]},
      {stage5_57[1]},
      {stage6_58[1],stage6_57[2],stage6_56[4],stage6_55[5],stage6_54[5]}
   );
   gpc606_5 gpc10860 (
      {stage5_56[2], stage5_56[3], stage5_56[4], stage5_56[5], stage5_56[6], stage5_56[7]},
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage6_60[0],stage6_59[0],stage6_58[2],stage6_57[3],stage6_56[5]}
   );
   gpc606_5 gpc10861 (
      {stage5_56[8], stage5_56[9], stage5_56[10], stage5_56[11], stage5_56[12], 1'b0},
      {stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9], stage5_58[10], stage5_58[11]},
      {stage6_60[1],stage6_59[1],stage6_58[3],stage6_57[4],stage6_56[6]}
   );
   gpc606_5 gpc10862 (
      {stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5], stage5_57[6], stage5_57[7]},
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage6_61[0],stage6_60[2],stage6_59[2],stage6_58[4],stage6_57[5]}
   );
   gpc606_5 gpc10863 (
      {stage5_58[12], stage5_58[13], stage5_58[14], stage5_58[15], stage5_58[16], stage5_58[17]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[1],stage6_60[3],stage6_59[3],stage6_58[5]}
   );
   gpc606_5 gpc10864 (
      {stage5_58[18], stage5_58[19], stage5_58[20], stage5_58[21], stage5_58[22], stage5_58[23]},
      {stage5_60[6], stage5_60[7], stage5_60[8], stage5_60[9], stage5_60[10], stage5_60[11]},
      {stage6_62[1],stage6_61[2],stage6_60[4],stage6_59[4],stage6_58[6]}
   );
   gpc1343_5 gpc10865 (
      {stage5_61[0], stage5_61[1], stage5_61[2]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3]},
      {stage5_63[0], stage5_63[1], stage5_63[2]},
      {stage5_64[0]},
      {stage6_65[0],stage6_64[0],stage6_63[0],stage6_62[2],stage6_61[3]}
   );
   gpc1343_5 gpc10866 (
      {stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage5_62[4], stage5_62[5], stage5_62[6], stage5_62[7]},
      {stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage5_64[1]},
      {stage6_65[1],stage6_64[1],stage6_63[1],stage6_62[3],stage6_61[4]}
   );
   gpc606_5 gpc10867 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], 1'b0, 1'b0},
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], 1'b0},
      {stage6_65[2],stage6_64[2],stage6_63[2],stage6_62[4],stage6_61[5]}
   );
   gpc117_4 gpc10868 (
      {stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5], stage5_64[6], stage5_64[7], stage5_64[8]},
      {stage5_65[0]},
      {stage5_66[0]},
      {stage6_67[0],stage6_66[0],stage6_65[3],stage6_64[3]}
   );
   gpc606_5 gpc10869 (
      {stage5_64[9], stage5_64[10], stage5_64[11], stage5_64[12], stage5_64[13], stage5_64[14]},
      {stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], stage5_66[5], stage5_66[6]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[4],stage6_64[4]}
   );
   gpc615_5 gpc10870 (
      {stage5_64[15], stage5_64[16], stage5_64[17], stage5_64[18], stage5_64[19]},
      {stage5_65[1]},
      {stage5_66[7], stage5_66[8], stage5_66[9], stage5_66[10], stage5_66[11], stage5_66[12]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[5],stage6_64[5]}
   );
   gpc2135_5 gpc10871 (
      {stage5_67[0], stage5_67[1], stage5_67[2], stage5_67[3], stage5_67[4]},
      {stage5_68[0], stage5_68[1], stage5_68[2]},
      {stage5_69[0]},
      {stage5_70[0], stage5_70[1]},
      {stage6_71[0],stage6_70[0],stage6_69[0],stage6_68[2],stage6_67[3]}
   );
   gpc2135_5 gpc10872 (
      {stage5_67[5], stage5_67[6], stage5_67[7], 1'b0, 1'b0},
      {stage5_68[3], stage5_68[4], stage5_68[5]},
      {stage5_69[1]},
      {stage5_70[2], stage5_70[3]},
      {stage6_71[1],stage6_70[1],stage6_69[1],stage6_68[3],stage6_67[4]}
   );
   gpc1_1 gpc10873 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc10874 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc10875 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc10876 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc10877 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc10878 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc10879 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc10880 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc10881 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc10882 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc10883 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc10884 (
      {stage5_3[5]},
      {stage6_3[1]}
   );
   gpc1_1 gpc10885 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc10886 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc10887 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc10888 (
      {stage5_5[18]},
      {stage6_5[4]}
   );
   gpc1_1 gpc10889 (
      {stage5_5[19]},
      {stage6_5[5]}
   );
   gpc1_1 gpc10890 (
      {stage5_5[20]},
      {stage6_5[6]}
   );
   gpc1_1 gpc10891 (
      {stage5_16[12]},
      {stage6_16[4]}
   );
   gpc1_1 gpc10892 (
      {stage5_16[13]},
      {stage6_16[5]}
   );
   gpc1_1 gpc10893 (
      {stage5_21[9]},
      {stage6_21[4]}
   );
   gpc1_1 gpc10894 (
      {stage5_21[10]},
      {stage6_21[5]}
   );
   gpc1_1 gpc10895 (
      {stage5_22[6]},
      {stage6_22[3]}
   );
   gpc1_1 gpc10896 (
      {stage5_22[7]},
      {stage6_22[4]}
   );
   gpc1_1 gpc10897 (
      {stage5_22[8]},
      {stage6_22[5]}
   );
   gpc1_1 gpc10898 (
      {stage5_22[9]},
      {stage6_22[6]}
   );
   gpc1_1 gpc10899 (
      {stage5_22[10]},
      {stage6_22[7]}
   );
   gpc1_1 gpc10900 (
      {stage5_22[11]},
      {stage6_22[8]}
   );
   gpc1_1 gpc10901 (
      {stage5_22[12]},
      {stage6_22[9]}
   );
   gpc1_1 gpc10902 (
      {stage5_22[13]},
      {stage6_22[10]}
   );
   gpc1_1 gpc10903 (
      {stage5_22[14]},
      {stage6_22[11]}
   );
   gpc1_1 gpc10904 (
      {stage5_23[9]},
      {stage6_23[4]}
   );
   gpc1_1 gpc10905 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc10906 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc10907 (
      {stage5_24[6]},
      {stage6_24[4]}
   );
   gpc1_1 gpc10908 (
      {stage5_24[7]},
      {stage6_24[5]}
   );
   gpc1_1 gpc10909 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc10910 (
      {stage5_25[6]},
      {stage6_25[2]}
   );
   gpc1_1 gpc10911 (
      {stage5_25[7]},
      {stage6_25[3]}
   );
   gpc1_1 gpc10912 (
      {stage5_25[8]},
      {stage6_25[4]}
   );
   gpc1_1 gpc10913 (
      {stage5_25[9]},
      {stage6_25[5]}
   );
   gpc1_1 gpc10914 (
      {stage5_25[10]},
      {stage6_25[6]}
   );
   gpc1_1 gpc10915 (
      {stage5_25[11]},
      {stage6_25[7]}
   );
   gpc1_1 gpc10916 (
      {stage5_25[12]},
      {stage6_25[8]}
   );
   gpc1_1 gpc10917 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc10918 (
      {stage5_30[7]},
      {stage6_30[6]}
   );
   gpc1_1 gpc10919 (
      {stage5_30[8]},
      {stage6_30[7]}
   );
   gpc1_1 gpc10920 (
      {stage5_33[7]},
      {stage6_33[6]}
   );
   gpc1_1 gpc10921 (
      {stage5_33[8]},
      {stage6_33[7]}
   );
   gpc1_1 gpc10922 (
      {stage5_34[20]},
      {stage6_34[5]}
   );
   gpc1_1 gpc10923 (
      {stage5_39[10]},
      {stage6_39[4]}
   );
   gpc1_1 gpc10924 (
      {stage5_40[17]},
      {stage6_40[7]}
   );
   gpc1_1 gpc10925 (
      {stage5_40[18]},
      {stage6_40[8]}
   );
   gpc1_1 gpc10926 (
      {stage5_40[19]},
      {stage6_40[9]}
   );
   gpc1_1 gpc10927 (
      {stage5_41[2]},
      {stage6_41[4]}
   );
   gpc1_1 gpc10928 (
      {stage5_41[3]},
      {stage6_41[5]}
   );
   gpc1_1 gpc10929 (
      {stage5_41[4]},
      {stage6_41[6]}
   );
   gpc1_1 gpc10930 (
      {stage5_41[5]},
      {stage6_41[7]}
   );
   gpc1_1 gpc10931 (
      {stage5_41[6]},
      {stage6_41[8]}
   );
   gpc1_1 gpc10932 (
      {stage5_41[7]},
      {stage6_41[9]}
   );
   gpc1_1 gpc10933 (
      {stage5_41[8]},
      {stage6_41[10]}
   );
   gpc1_1 gpc10934 (
      {stage5_49[14]},
      {stage6_49[7]}
   );
   gpc1_1 gpc10935 (
      {stage5_49[15]},
      {stage6_49[8]}
   );
   gpc1_1 gpc10936 (
      {stage5_49[16]},
      {stage6_49[9]}
   );
   gpc1_1 gpc10937 (
      {stage5_52[12]},
      {stage6_52[7]}
   );
   gpc1_1 gpc10938 (
      {stage5_57[8]},
      {stage6_57[6]}
   );
   gpc1_1 gpc10939 (
      {stage5_60[12]},
      {stage6_60[5]}
   );
   gpc1_1 gpc10940 (
      {stage5_60[13]},
      {stage6_60[6]}
   );
   gpc1_1 gpc10941 (
      {stage5_65[2]},
      {stage6_65[6]}
   );
   gpc1_1 gpc10942 (
      {stage5_65[3]},
      {stage6_65[7]}
   );
   gpc1_1 gpc10943 (
      {stage5_65[4]},
      {stage6_65[8]}
   );
   gpc1_1 gpc10944 (
      {stage5_65[5]},
      {stage6_65[9]}
   );
   gpc1_1 gpc10945 (
      {stage5_68[6]},
      {stage6_68[4]}
   );
   gpc1_1 gpc10946 (
      {stage5_68[7]},
      {stage6_68[5]}
   );
   gpc1_1 gpc10947 (
      {stage5_68[8]},
      {stage6_68[6]}
   );
   gpc1_1 gpc10948 (
      {stage5_68[9]},
      {stage6_68[7]}
   );
   gpc1_1 gpc10949 (
      {stage5_68[10]},
      {stage6_68[8]}
   );
   gpc1_1 gpc10950 (
      {stage5_68[11]},
      {stage6_68[9]}
   );
   gpc1_1 gpc10951 (
      {stage5_69[2]},
      {stage6_69[2]}
   );
   gpc135_4 gpc10952 (
      {stage6_4[0], stage6_4[1], stage6_4[2], 1'b0, 1'b0},
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc615_5 gpc10953 (
      {stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_7[0]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1],stage7_6[1]}
   );
   gpc15_3 gpc10954 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc623_5 gpc10955 (
      {stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[2]}
   );
   gpc23_3 gpc10956 (
      {stage6_11[2], stage6_11[3], stage6_11[4]},
      {stage6_12[6], stage6_12[7]},
      {stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc117_4 gpc10957 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage6_15[0]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1]}
   );
   gpc7_3 gpc10958 (
      {stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5], stage6_15[6], stage6_15[7]},
      {stage7_17[1],stage7_16[1],stage7_15[1]}
   );
   gpc15_3 gpc10959 (
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4]},
      {stage6_18[0]},
      {stage7_19[0],stage7_18[0],stage7_17[2]}
   );
   gpc606_5 gpc10960 (
      {stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5], stage6_18[6]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[1],stage7_18[1]}
   );
   gpc1163_5 gpc10961 (
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_23[0]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1]}
   );
   gpc1163_5 gpc10962 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[6], stage6_22[7], stage6_22[8], stage6_22[9], stage6_22[10], stage6_22[11]},
      {stage6_23[1]},
      {stage6_24[1]},
      {stage7_25[1],stage7_24[1],stage7_23[1],stage7_22[2],stage7_21[2]}
   );
   gpc15_3 gpc10963 (
      {stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5], stage6_24[6]},
      {stage6_25[0]},
      {stage7_26[0],stage7_25[2],stage7_24[2]}
   );
   gpc606_5 gpc10964 (
      {stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5], stage6_25[6]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], 1'b0},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[3]}
   );
   gpc606_5 gpc10965 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], 1'b0, 1'b0},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[1]}
   );
   gpc1406_5 gpc10966 (
      {stage6_29[0], stage6_29[1], stage6_29[2], stage6_29[3], stage6_29[4], stage6_29[5]},
      {stage6_31[0], stage6_31[1], stage6_31[2], 1'b0},
      {stage6_32[0]},
      {stage7_33[0],stage7_32[1],stage7_31[1],stage7_30[1],stage7_29[2]}
   );
   gpc135_4 gpc10967 (
      {stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage6_33[0], stage6_33[1], stage6_33[2]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[1],stage7_32[2]}
   );
   gpc15_3 gpc10968 (
      {stage6_33[3], stage6_33[4], stage6_33[5], stage6_33[6], stage6_33[7]},
      {stage6_34[1]},
      {stage7_35[1],stage7_34[1],stage7_33[2]}
   );
   gpc117_4 gpc10969 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage6_37[0]},
      {stage6_38[0]},
      {stage7_39[0],stage7_38[0],stage7_37[0],stage7_36[0]}
   );
   gpc15_3 gpc10970 (
      {stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_38[1]},
      {stage7_39[1],stage7_38[1],stage7_37[1]}
   );
   gpc3_2 gpc10971 (
      {stage6_38[2], stage6_38[3], stage6_38[4]},
      {stage7_39[2],stage7_38[2]}
   );
   gpc2135_5 gpc10972 (
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], stage6_39[4]},
      {stage6_40[0], stage6_40[1], stage6_40[2]},
      {stage6_41[0]},
      {stage6_42[0], stage6_42[1]},
      {stage7_43[0],stage7_42[0],stage7_41[0],stage7_40[0],stage7_39[3]}
   );
   gpc207_4 gpc10973 (
      {stage6_40[3], stage6_40[4], stage6_40[5], stage6_40[6], stage6_40[7], stage6_40[8], stage6_40[9]},
      {stage6_42[2], stage6_42[3]},
      {stage7_43[1],stage7_42[1],stage7_41[1],stage7_40[1]}
   );
   gpc7_3 gpc10974 (
      {stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4], stage6_41[5], stage6_41[6], stage6_41[7]},
      {stage7_43[2],stage7_42[2],stage7_41[2]}
   );
   gpc215_4 gpc10975 (
      {stage6_43[0], stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4]},
      {stage6_44[0]},
      {stage6_45[0], stage6_45[1]},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[3]}
   );
   gpc207_4 gpc10976 (
      {stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], stage6_44[5], stage6_44[6], stage6_44[7]},
      {stage6_46[0], stage6_46[1]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1]}
   );
   gpc615_5 gpc10977 (
      {stage6_47[0], stage6_47[1], stage6_47[2], stage6_47[3], 1'b0},
      {stage6_48[0]},
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage7_51[0],stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1]}
   );
   gpc7_3 gpc10978 (
      {stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5], 1'b0, 1'b0},
      {stage7_50[1],stage7_49[1],stage7_48[1]}
   );
   gpc615_5 gpc10979 (
      {stage6_50[0], stage6_50[1], stage6_50[2], stage6_50[3], stage6_50[4]},
      {stage6_51[0]},
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4], stage6_52[5]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[2]}
   );
   gpc1343_5 gpc10980 (
      {stage6_52[6], stage6_52[7], 1'b0},
      {stage6_53[0], stage6_53[1], stage6_53[2], stage6_53[3]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc15_3 gpc10981 (
      {stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4], stage6_55[5]},
      {stage6_56[0]},
      {stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1423_5 gpc10982 (
      {stage6_56[1], stage6_56[2], stage6_56[3]},
      {stage6_57[0], stage6_57[1]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3]},
      {stage6_59[0]},
      {stage7_60[0],stage7_59[0],stage7_58[0],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc10983 (
      {stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5], stage6_57[6]},
      {stage6_58[4], stage6_58[5], stage6_58[6]},
      {stage6_59[1]},
      {stage7_60[1],stage7_59[1],stage7_58[1],stage7_57[2]}
   );
   gpc606_5 gpc10984 (
      {stage6_59[2], stage6_59[3], stage6_59[4], 1'b0, 1'b0, 1'b0},
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4], stage6_61[5]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[2],stage7_59[2]}
   );
   gpc606_5 gpc10985 (
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3], stage6_60[4], stage6_60[5]},
      {stage6_62[0], stage6_62[1], stage6_62[2], stage6_62[3], stage6_62[4], 1'b0},
      {stage7_64[0],stage7_63[1],stage7_62[1],stage7_61[1],stage7_60[3]}
   );
   gpc3_2 gpc10986 (
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage7_65[0],stage7_64[1]}
   );
   gpc3_2 gpc10987 (
      {stage6_64[3], stage6_64[4], stage6_64[5]},
      {stage7_65[1],stage7_64[2]}
   );
   gpc1163_5 gpc10988 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[0]}
   );
   gpc117_4 gpc10989 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc1_1 gpc10990 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc10991 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc10992 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc10993 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc10994 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc10995 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc10996 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc10997 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc10998 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc10999 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc11000 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc11001 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc11002 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc11003 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc11004 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc11005 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc11006 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc11007 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc11008 (
      {stage6_5[6]},
      {stage7_5[4]}
   );
   gpc1_1 gpc11009 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc11010 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc11011 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc11012 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc11013 (
      {stage6_7[5]},
      {stage7_7[6]}
   );
   gpc1_1 gpc11014 (
      {stage6_9[5]},
      {stage7_9[2]}
   );
   gpc1_1 gpc11015 (
      {stage6_9[6]},
      {stage7_9[3]}
   );
   gpc1_1 gpc11016 (
      {stage6_9[7]},
      {stage7_9[4]}
   );
   gpc1_1 gpc11017 (
      {stage6_10[4]},
      {stage7_10[3]}
   );
   gpc1_1 gpc11018 (
      {stage6_11[5]},
      {stage7_11[3]}
   );
   gpc1_1 gpc11019 (
      {stage6_13[0]},
      {stage7_13[2]}
   );
   gpc1_1 gpc11020 (
      {stage6_13[1]},
      {stage7_13[3]}
   );
   gpc1_1 gpc11021 (
      {stage6_13[2]},
      {stage7_13[4]}
   );
   gpc1_1 gpc11022 (
      {stage6_13[3]},
      {stage7_13[5]}
   );
   gpc1_1 gpc11023 (
      {stage6_13[4]},
      {stage7_13[6]}
   );
   gpc1_1 gpc11024 (
      {stage6_14[7]},
      {stage7_14[2]}
   );
   gpc1_1 gpc11025 (
      {stage6_16[1]},
      {stage7_16[2]}
   );
   gpc1_1 gpc11026 (
      {stage6_16[2]},
      {stage7_16[3]}
   );
   gpc1_1 gpc11027 (
      {stage6_16[3]},
      {stage7_16[4]}
   );
   gpc1_1 gpc11028 (
      {stage6_16[4]},
      {stage7_16[5]}
   );
   gpc1_1 gpc11029 (
      {stage6_16[5]},
      {stage7_16[6]}
   );
   gpc1_1 gpc11030 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc11031 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc11032 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc11033 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc11034 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc11035 (
      {stage6_23[2]},
      {stage7_23[2]}
   );
   gpc1_1 gpc11036 (
      {stage6_23[3]},
      {stage7_23[3]}
   );
   gpc1_1 gpc11037 (
      {stage6_23[4]},
      {stage7_23[4]}
   );
   gpc1_1 gpc11038 (
      {stage6_23[5]},
      {stage7_23[5]}
   );
   gpc1_1 gpc11039 (
      {stage6_23[6]},
      {stage7_23[6]}
   );
   gpc1_1 gpc11040 (
      {stage6_25[7]},
      {stage7_25[4]}
   );
   gpc1_1 gpc11041 (
      {stage6_25[8]},
      {stage7_25[5]}
   );
   gpc1_1 gpc11042 (
      {stage6_26[0]},
      {stage7_26[2]}
   );
   gpc1_1 gpc11043 (
      {stage6_26[1]},
      {stage7_26[3]}
   );
   gpc1_1 gpc11044 (
      {stage6_26[2]},
      {stage7_26[4]}
   );
   gpc1_1 gpc11045 (
      {stage6_26[3]},
      {stage7_26[5]}
   );
   gpc1_1 gpc11046 (
      {stage6_26[4]},
      {stage7_26[6]}
   );
   gpc1_1 gpc11047 (
      {stage6_30[6]},
      {stage7_30[2]}
   );
   gpc1_1 gpc11048 (
      {stage6_30[7]},
      {stage7_30[3]}
   );
   gpc1_1 gpc11049 (
      {stage6_34[2]},
      {stage7_34[2]}
   );
   gpc1_1 gpc11050 (
      {stage6_34[3]},
      {stage7_34[3]}
   );
   gpc1_1 gpc11051 (
      {stage6_34[4]},
      {stage7_34[4]}
   );
   gpc1_1 gpc11052 (
      {stage6_34[5]},
      {stage7_34[5]}
   );
   gpc1_1 gpc11053 (
      {stage6_35[0]},
      {stage7_35[2]}
   );
   gpc1_1 gpc11054 (
      {stage6_35[1]},
      {stage7_35[3]}
   );
   gpc1_1 gpc11055 (
      {stage6_35[2]},
      {stage7_35[4]}
   );
   gpc1_1 gpc11056 (
      {stage6_35[3]},
      {stage7_35[5]}
   );
   gpc1_1 gpc11057 (
      {stage6_35[4]},
      {stage7_35[6]}
   );
   gpc1_1 gpc11058 (
      {stage6_36[7]},
      {stage7_36[1]}
   );
   gpc1_1 gpc11059 (
      {stage6_41[8]},
      {stage7_41[3]}
   );
   gpc1_1 gpc11060 (
      {stage6_41[9]},
      {stage7_41[4]}
   );
   gpc1_1 gpc11061 (
      {stage6_41[10]},
      {stage7_41[5]}
   );
   gpc1_1 gpc11062 (
      {stage6_45[2]},
      {stage7_45[2]}
   );
   gpc1_1 gpc11063 (
      {stage6_45[3]},
      {stage7_45[3]}
   );
   gpc1_1 gpc11064 (
      {stage6_45[4]},
      {stage7_45[4]}
   );
   gpc1_1 gpc11065 (
      {stage6_45[5]},
      {stage7_45[5]}
   );
   gpc1_1 gpc11066 (
      {stage6_45[6]},
      {stage7_45[6]}
   );
   gpc1_1 gpc11067 (
      {stage6_46[2]},
      {stage7_46[2]}
   );
   gpc1_1 gpc11068 (
      {stage6_46[3]},
      {stage7_46[3]}
   );
   gpc1_1 gpc11069 (
      {stage6_46[4]},
      {stage7_46[4]}
   );
   gpc1_1 gpc11070 (
      {stage6_46[5]},
      {stage7_46[5]}
   );
   gpc1_1 gpc11071 (
      {stage6_46[6]},
      {stage7_46[6]}
   );
   gpc1_1 gpc11072 (
      {stage6_49[6]},
      {stage7_49[2]}
   );
   gpc1_1 gpc11073 (
      {stage6_49[7]},
      {stage7_49[3]}
   );
   gpc1_1 gpc11074 (
      {stage6_49[8]},
      {stage7_49[4]}
   );
   gpc1_1 gpc11075 (
      {stage6_49[9]},
      {stage7_49[5]}
   );
   gpc1_1 gpc11076 (
      {stage6_51[1]},
      {stage7_51[2]}
   );
   gpc1_1 gpc11077 (
      {stage6_51[2]},
      {stage7_51[3]}
   );
   gpc1_1 gpc11078 (
      {stage6_51[3]},
      {stage7_51[4]}
   );
   gpc1_1 gpc11079 (
      {stage6_51[4]},
      {stage7_51[5]}
   );
   gpc1_1 gpc11080 (
      {stage6_54[3]},
      {stage7_54[2]}
   );
   gpc1_1 gpc11081 (
      {stage6_54[4]},
      {stage7_54[3]}
   );
   gpc1_1 gpc11082 (
      {stage6_54[5]},
      {stage7_54[4]}
   );
   gpc1_1 gpc11083 (
      {stage6_56[4]},
      {stage7_56[3]}
   );
   gpc1_1 gpc11084 (
      {stage6_56[5]},
      {stage7_56[4]}
   );
   gpc1_1 gpc11085 (
      {stage6_56[6]},
      {stage7_56[5]}
   );
   gpc1_1 gpc11086 (
      {stage6_60[6]},
      {stage7_60[4]}
   );
   gpc1_1 gpc11087 (
      {stage6_63[0]},
      {stage7_63[2]}
   );
   gpc1_1 gpc11088 (
      {stage6_63[1]},
      {stage7_63[3]}
   );
   gpc1_1 gpc11089 (
      {stage6_63[2]},
      {stage7_63[4]}
   );
   gpc1_1 gpc11090 (
      {stage6_65[0]},
      {stage7_65[2]}
   );
   gpc1_1 gpc11091 (
      {stage6_65[1]},
      {stage7_65[3]}
   );
   gpc1_1 gpc11092 (
      {stage6_65[2]},
      {stage7_65[4]}
   );
   gpc1_1 gpc11093 (
      {stage6_65[3]},
      {stage7_65[5]}
   );
   gpc1_1 gpc11094 (
      {stage6_65[4]},
      {stage7_65[6]}
   );
   gpc1_1 gpc11095 (
      {stage6_65[5]},
      {stage7_65[7]}
   );
   gpc1_1 gpc11096 (
      {stage6_65[6]},
      {stage7_65[8]}
   );
   gpc1_1 gpc11097 (
      {stage6_65[7]},
      {stage7_65[9]}
   );
   gpc1_1 gpc11098 (
      {stage6_65[8]},
      {stage7_65[10]}
   );
   gpc1_1 gpc11099 (
      {stage6_65[9]},
      {stage7_65[11]}
   );
   gpc1_1 gpc11100 (
      {stage6_68[8]},
      {stage7_68[2]}
   );
   gpc1_1 gpc11101 (
      {stage6_68[9]},
      {stage7_68[3]}
   );
   gpc1_1 gpc11102 (
      {stage6_69[2]},
      {stage7_69[2]}
   );
   gpc1_1 gpc11103 (
      {stage6_70[1]},
      {stage7_70[2]}
   );
   gpc1_1 gpc11104 (
      {stage6_71[0]},
      {stage7_71[1]}
   );
   gpc1_1 gpc11105 (
      {stage6_71[1]},
      {stage7_71[2]}
   );
   gpc615_5 gpc11106 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], 1'b0, 1'b0, 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1415_5 gpc11107 (
      {stage7_3[0], stage7_3[1], stage7_3[2], stage7_3[3], 1'b0},
      {stage7_4[0]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc7_3 gpc11108 (
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5], stage7_7[6]},
      {stage8_9[0],stage8_8[0],stage8_7[1]}
   );
   gpc1415_5 gpc11109 (
      {stage7_9[0], stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4]},
      {stage7_10[0]},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc3_2 gpc11110 (
      {stage7_10[1], stage7_10[2], stage7_10[3]},
      {stage8_11[1],stage8_10[1]}
   );
   gpc7_3 gpc11111 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], stage7_13[6]},
      {stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc623_5 gpc11112 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[0], stage7_15[1]},
      {stage7_16[0], stage7_16[1], stage7_16[2], stage7_16[3], stage7_16[4], stage7_16[5]},
      {stage8_18[0],stage8_17[0],stage8_16[0],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc11113 (
      {stage7_17[0], stage7_17[1], stage7_17[2]},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc2223_5 gpc11114 (
      {stage7_21[0], stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1]},
      {stage7_23[0], stage7_23[1]},
      {stage7_24[0], stage7_24[1]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1]}
   );
   gpc615_5 gpc11115 (
      {stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[2]},
      {stage7_25[0], stage7_25[1], stage7_25[2], stage7_25[3], stage7_25[4], stage7_25[5]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc117_4 gpc11116 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], stage7_26[6]},
      {stage7_27[0]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[0],stage8_27[1],stage8_26[1]}
   );
   gpc15_3 gpc11117 (
      {stage7_29[0], stage7_29[1], stage7_29[2], 1'b0, 1'b0},
      {stage7_30[0]},
      {stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc2223_5 gpc11118 (
      {stage7_30[1], stage7_30[2], stage7_30[3]},
      {stage7_31[0], stage7_31[1]},
      {stage7_32[0], stage7_32[1]},
      {stage7_33[0], stage7_33[1]},
      {stage8_34[0],stage8_33[0],stage8_32[0],stage8_31[1],stage8_30[1]}
   );
   gpc207_4 gpc11119 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc207_4 gpc11120 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], stage7_35[6]},
      {stage7_37[0], stage7_37[1]},
      {stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc3_2 gpc11121 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage8_39[0],stage8_38[1]}
   );
   gpc2116_5 gpc11122 (
      {stage7_39[0], stage7_39[1], stage7_39[2], stage7_39[3], 1'b0, 1'b0},
      {stage7_40[0]},
      {stage7_41[0]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[0],stage8_39[1]}
   );
   gpc1415_5 gpc11123 (
      {stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4], stage7_41[5]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc207_4 gpc11124 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4], stage7_45[5], stage7_45[6]},
      {stage7_47[0], stage7_47[1]},
      {stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc11125 (
      {stage7_46[0], stage7_46[1], stage7_46[2], stage7_46[3], stage7_46[4], stage7_46[5], stage7_46[6]},
      {stage7_48[0], stage7_48[1]},
      {stage8_49[0],stage8_48[1],stage8_47[1],stage8_46[1]}
   );
   gpc207_4 gpc11126 (
      {stage7_49[0], stage7_49[1], stage7_49[2], stage7_49[3], stage7_49[4], stage7_49[5], 1'b0},
      {stage7_51[0], stage7_51[1]},
      {stage8_52[0],stage8_51[0],stage8_50[0],stage8_49[1]}
   );
   gpc1343_5 gpc11127 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage7_51[2], stage7_51[3], stage7_51[4], stage7_51[5]},
      {stage7_52[0], stage7_52[1], 1'b0},
      {stage7_53[0]},
      {stage8_54[0],stage8_53[0],stage8_52[1],stage8_51[1],stage8_50[1]}
   );
   gpc1415_5 gpc11128 (
      {stage7_54[0], stage7_54[1], stage7_54[2], stage7_54[3], stage7_54[4]},
      {stage7_55[0]},
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3]},
      {stage7_57[0]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[0],stage8_54[1]}
   );
   gpc2223_5 gpc11129 (
      {stage7_56[4], stage7_56[5], 1'b0},
      {stage7_57[1], stage7_57[2]},
      {stage7_58[0], stage7_58[1]},
      {stage7_59[0], stage7_59[1]},
      {stage8_60[0],stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc215_4 gpc11130 (
      {stage7_60[0], stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4]},
      {stage7_61[0]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[0],stage8_61[0],stage8_60[1]}
   );
   gpc606_5 gpc11131 (
      {stage7_63[0], stage7_63[1], stage7_63[2], stage7_63[3], stage7_63[4], 1'b0},
      {stage7_65[0], stage7_65[1], stage7_65[2], stage7_65[3], stage7_65[4], stage7_65[5]},
      {stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[0],stage8_63[1]}
   );
   gpc1163_5 gpc11132 (
      {stage7_64[0], stage7_64[1], stage7_64[2]},
      {stage7_65[6], stage7_65[7], stage7_65[8], stage7_65[9], stage7_65[10], stage7_65[11]},
      {stage7_66[0]},
      {stage7_67[0]},
      {stage8_68[0],stage8_67[1],stage8_66[1],stage8_65[1],stage8_64[1]}
   );
   gpc606_5 gpc11133 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], 1'b0, 1'b0},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc11134 (
      {stage7_69[0], stage7_69[1], stage7_69[2], 1'b0, 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], stage7_71[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc11135 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc11136 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc11137 (
      {stage7_5[4]},
      {stage8_5[1]}
   );
   gpc1_1 gpc11138 (
      {stage7_6[1]},
      {stage8_6[1]}
   );
   gpc1_1 gpc11139 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc11140 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc11141 (
      {stage7_16[6]},
      {stage8_16[1]}
   );
   gpc1_1 gpc11142 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc11143 (
      {stage7_20[0]},
      {stage8_20[1]}
   );
   gpc1_1 gpc11144 (
      {stage7_22[2]},
      {stage8_22[1]}
   );
   gpc1_1 gpc11145 (
      {stage7_28[1]},
      {stage8_28[1]}
   );
   gpc1_1 gpc11146 (
      {stage7_32[2]},
      {stage8_32[1]}
   );
   gpc1_1 gpc11147 (
      {stage7_33[2]},
      {stage8_33[1]}
   );
   gpc1_1 gpc11148 (
      {stage7_40[1]},
      {stage8_40[1]}
   );
   gpc1_1 gpc11149 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc11150 (
      {stage7_53[1]},
      {stage8_53[1]}
   );
   gpc1_1 gpc11151 (
      {stage7_55[1]},
      {stage8_55[1]}
   );
   gpc1_1 gpc11152 (
      {stage7_59[2]},
      {stage8_59[1]}
   );
   gpc1_1 gpc11153 (
      {stage7_61[1]},
      {stage8_61[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor_CLA512_64 compressor_CLA512_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485] + src32[486] + src32[487] + src32[488] + src32[489] + src32[490] + src32[491] + src32[492] + src32[493] + src32[494] + src32[495] + src32[496] + src32[497] + src32[498] + src32[499] + src32[500] + src32[501] + src32[502] + src32[503] + src32[504] + src32[505] + src32[506] + src32[507] + src32[508] + src32[509] + src32[510] + src32[511])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485] + src33[486] + src33[487] + src33[488] + src33[489] + src33[490] + src33[491] + src33[492] + src33[493] + src33[494] + src33[495] + src33[496] + src33[497] + src33[498] + src33[499] + src33[500] + src33[501] + src33[502] + src33[503] + src33[504] + src33[505] + src33[506] + src33[507] + src33[508] + src33[509] + src33[510] + src33[511])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485] + src34[486] + src34[487] + src34[488] + src34[489] + src34[490] + src34[491] + src34[492] + src34[493] + src34[494] + src34[495] + src34[496] + src34[497] + src34[498] + src34[499] + src34[500] + src34[501] + src34[502] + src34[503] + src34[504] + src34[505] + src34[506] + src34[507] + src34[508] + src34[509] + src34[510] + src34[511])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485] + src35[486] + src35[487] + src35[488] + src35[489] + src35[490] + src35[491] + src35[492] + src35[493] + src35[494] + src35[495] + src35[496] + src35[497] + src35[498] + src35[499] + src35[500] + src35[501] + src35[502] + src35[503] + src35[504] + src35[505] + src35[506] + src35[507] + src35[508] + src35[509] + src35[510] + src35[511])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485] + src36[486] + src36[487] + src36[488] + src36[489] + src36[490] + src36[491] + src36[492] + src36[493] + src36[494] + src36[495] + src36[496] + src36[497] + src36[498] + src36[499] + src36[500] + src36[501] + src36[502] + src36[503] + src36[504] + src36[505] + src36[506] + src36[507] + src36[508] + src36[509] + src36[510] + src36[511])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485] + src37[486] + src37[487] + src37[488] + src37[489] + src37[490] + src37[491] + src37[492] + src37[493] + src37[494] + src37[495] + src37[496] + src37[497] + src37[498] + src37[499] + src37[500] + src37[501] + src37[502] + src37[503] + src37[504] + src37[505] + src37[506] + src37[507] + src37[508] + src37[509] + src37[510] + src37[511])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485] + src38[486] + src38[487] + src38[488] + src38[489] + src38[490] + src38[491] + src38[492] + src38[493] + src38[494] + src38[495] + src38[496] + src38[497] + src38[498] + src38[499] + src38[500] + src38[501] + src38[502] + src38[503] + src38[504] + src38[505] + src38[506] + src38[507] + src38[508] + src38[509] + src38[510] + src38[511])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485] + src39[486] + src39[487] + src39[488] + src39[489] + src39[490] + src39[491] + src39[492] + src39[493] + src39[494] + src39[495] + src39[496] + src39[497] + src39[498] + src39[499] + src39[500] + src39[501] + src39[502] + src39[503] + src39[504] + src39[505] + src39[506] + src39[507] + src39[508] + src39[509] + src39[510] + src39[511])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485] + src40[486] + src40[487] + src40[488] + src40[489] + src40[490] + src40[491] + src40[492] + src40[493] + src40[494] + src40[495] + src40[496] + src40[497] + src40[498] + src40[499] + src40[500] + src40[501] + src40[502] + src40[503] + src40[504] + src40[505] + src40[506] + src40[507] + src40[508] + src40[509] + src40[510] + src40[511])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485] + src41[486] + src41[487] + src41[488] + src41[489] + src41[490] + src41[491] + src41[492] + src41[493] + src41[494] + src41[495] + src41[496] + src41[497] + src41[498] + src41[499] + src41[500] + src41[501] + src41[502] + src41[503] + src41[504] + src41[505] + src41[506] + src41[507] + src41[508] + src41[509] + src41[510] + src41[511])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485] + src42[486] + src42[487] + src42[488] + src42[489] + src42[490] + src42[491] + src42[492] + src42[493] + src42[494] + src42[495] + src42[496] + src42[497] + src42[498] + src42[499] + src42[500] + src42[501] + src42[502] + src42[503] + src42[504] + src42[505] + src42[506] + src42[507] + src42[508] + src42[509] + src42[510] + src42[511])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485] + src43[486] + src43[487] + src43[488] + src43[489] + src43[490] + src43[491] + src43[492] + src43[493] + src43[494] + src43[495] + src43[496] + src43[497] + src43[498] + src43[499] + src43[500] + src43[501] + src43[502] + src43[503] + src43[504] + src43[505] + src43[506] + src43[507] + src43[508] + src43[509] + src43[510] + src43[511])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485] + src44[486] + src44[487] + src44[488] + src44[489] + src44[490] + src44[491] + src44[492] + src44[493] + src44[494] + src44[495] + src44[496] + src44[497] + src44[498] + src44[499] + src44[500] + src44[501] + src44[502] + src44[503] + src44[504] + src44[505] + src44[506] + src44[507] + src44[508] + src44[509] + src44[510] + src44[511])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485] + src45[486] + src45[487] + src45[488] + src45[489] + src45[490] + src45[491] + src45[492] + src45[493] + src45[494] + src45[495] + src45[496] + src45[497] + src45[498] + src45[499] + src45[500] + src45[501] + src45[502] + src45[503] + src45[504] + src45[505] + src45[506] + src45[507] + src45[508] + src45[509] + src45[510] + src45[511])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485] + src46[486] + src46[487] + src46[488] + src46[489] + src46[490] + src46[491] + src46[492] + src46[493] + src46[494] + src46[495] + src46[496] + src46[497] + src46[498] + src46[499] + src46[500] + src46[501] + src46[502] + src46[503] + src46[504] + src46[505] + src46[506] + src46[507] + src46[508] + src46[509] + src46[510] + src46[511])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485] + src47[486] + src47[487] + src47[488] + src47[489] + src47[490] + src47[491] + src47[492] + src47[493] + src47[494] + src47[495] + src47[496] + src47[497] + src47[498] + src47[499] + src47[500] + src47[501] + src47[502] + src47[503] + src47[504] + src47[505] + src47[506] + src47[507] + src47[508] + src47[509] + src47[510] + src47[511])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485] + src48[486] + src48[487] + src48[488] + src48[489] + src48[490] + src48[491] + src48[492] + src48[493] + src48[494] + src48[495] + src48[496] + src48[497] + src48[498] + src48[499] + src48[500] + src48[501] + src48[502] + src48[503] + src48[504] + src48[505] + src48[506] + src48[507] + src48[508] + src48[509] + src48[510] + src48[511])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485] + src49[486] + src49[487] + src49[488] + src49[489] + src49[490] + src49[491] + src49[492] + src49[493] + src49[494] + src49[495] + src49[496] + src49[497] + src49[498] + src49[499] + src49[500] + src49[501] + src49[502] + src49[503] + src49[504] + src49[505] + src49[506] + src49[507] + src49[508] + src49[509] + src49[510] + src49[511])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485] + src50[486] + src50[487] + src50[488] + src50[489] + src50[490] + src50[491] + src50[492] + src50[493] + src50[494] + src50[495] + src50[496] + src50[497] + src50[498] + src50[499] + src50[500] + src50[501] + src50[502] + src50[503] + src50[504] + src50[505] + src50[506] + src50[507] + src50[508] + src50[509] + src50[510] + src50[511])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485] + src51[486] + src51[487] + src51[488] + src51[489] + src51[490] + src51[491] + src51[492] + src51[493] + src51[494] + src51[495] + src51[496] + src51[497] + src51[498] + src51[499] + src51[500] + src51[501] + src51[502] + src51[503] + src51[504] + src51[505] + src51[506] + src51[507] + src51[508] + src51[509] + src51[510] + src51[511])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485] + src52[486] + src52[487] + src52[488] + src52[489] + src52[490] + src52[491] + src52[492] + src52[493] + src52[494] + src52[495] + src52[496] + src52[497] + src52[498] + src52[499] + src52[500] + src52[501] + src52[502] + src52[503] + src52[504] + src52[505] + src52[506] + src52[507] + src52[508] + src52[509] + src52[510] + src52[511])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485] + src53[486] + src53[487] + src53[488] + src53[489] + src53[490] + src53[491] + src53[492] + src53[493] + src53[494] + src53[495] + src53[496] + src53[497] + src53[498] + src53[499] + src53[500] + src53[501] + src53[502] + src53[503] + src53[504] + src53[505] + src53[506] + src53[507] + src53[508] + src53[509] + src53[510] + src53[511])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485] + src54[486] + src54[487] + src54[488] + src54[489] + src54[490] + src54[491] + src54[492] + src54[493] + src54[494] + src54[495] + src54[496] + src54[497] + src54[498] + src54[499] + src54[500] + src54[501] + src54[502] + src54[503] + src54[504] + src54[505] + src54[506] + src54[507] + src54[508] + src54[509] + src54[510] + src54[511])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485] + src55[486] + src55[487] + src55[488] + src55[489] + src55[490] + src55[491] + src55[492] + src55[493] + src55[494] + src55[495] + src55[496] + src55[497] + src55[498] + src55[499] + src55[500] + src55[501] + src55[502] + src55[503] + src55[504] + src55[505] + src55[506] + src55[507] + src55[508] + src55[509] + src55[510] + src55[511])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485] + src56[486] + src56[487] + src56[488] + src56[489] + src56[490] + src56[491] + src56[492] + src56[493] + src56[494] + src56[495] + src56[496] + src56[497] + src56[498] + src56[499] + src56[500] + src56[501] + src56[502] + src56[503] + src56[504] + src56[505] + src56[506] + src56[507] + src56[508] + src56[509] + src56[510] + src56[511])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485] + src57[486] + src57[487] + src57[488] + src57[489] + src57[490] + src57[491] + src57[492] + src57[493] + src57[494] + src57[495] + src57[496] + src57[497] + src57[498] + src57[499] + src57[500] + src57[501] + src57[502] + src57[503] + src57[504] + src57[505] + src57[506] + src57[507] + src57[508] + src57[509] + src57[510] + src57[511])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485] + src58[486] + src58[487] + src58[488] + src58[489] + src58[490] + src58[491] + src58[492] + src58[493] + src58[494] + src58[495] + src58[496] + src58[497] + src58[498] + src58[499] + src58[500] + src58[501] + src58[502] + src58[503] + src58[504] + src58[505] + src58[506] + src58[507] + src58[508] + src58[509] + src58[510] + src58[511])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485] + src59[486] + src59[487] + src59[488] + src59[489] + src59[490] + src59[491] + src59[492] + src59[493] + src59[494] + src59[495] + src59[496] + src59[497] + src59[498] + src59[499] + src59[500] + src59[501] + src59[502] + src59[503] + src59[504] + src59[505] + src59[506] + src59[507] + src59[508] + src59[509] + src59[510] + src59[511])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485] + src60[486] + src60[487] + src60[488] + src60[489] + src60[490] + src60[491] + src60[492] + src60[493] + src60[494] + src60[495] + src60[496] + src60[497] + src60[498] + src60[499] + src60[500] + src60[501] + src60[502] + src60[503] + src60[504] + src60[505] + src60[506] + src60[507] + src60[508] + src60[509] + src60[510] + src60[511])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485] + src61[486] + src61[487] + src61[488] + src61[489] + src61[490] + src61[491] + src61[492] + src61[493] + src61[494] + src61[495] + src61[496] + src61[497] + src61[498] + src61[499] + src61[500] + src61[501] + src61[502] + src61[503] + src61[504] + src61[505] + src61[506] + src61[507] + src61[508] + src61[509] + src61[510] + src61[511])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485] + src62[486] + src62[487] + src62[488] + src62[489] + src62[490] + src62[491] + src62[492] + src62[493] + src62[494] + src62[495] + src62[496] + src62[497] + src62[498] + src62[499] + src62[500] + src62[501] + src62[502] + src62[503] + src62[504] + src62[505] + src62[506] + src62[507] + src62[508] + src62[509] + src62[510] + src62[511])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485] + src63[486] + src63[487] + src63[488] + src63[489] + src63[490] + src63[491] + src63[492] + src63[493] + src63[494] + src63[495] + src63[496] + src63[497] + src63[498] + src63[499] + src63[500] + src63[501] + src63[502] + src63[503] + src63[504] + src63[505] + src63[506] + src63[507] + src63[508] + src63[509] + src63[510] + src63[511])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hab68f38290d2df7a12e1b3a198b67d2d0458b9ad4de4d97b603ef4797d82a0aad185b512eac6b258dcb8d9cb418526908ab6d6c581d9236c63b2cf6ad17abe3a4f89505e250d024bbcb8eebaba293800ec51e089cbced0eb157d7f83368abb34113a9b9f744f7e54c5a264cc47889763e2e52cce8a9ca1b52fd81eeaaa7a8778b613b8ed800cda3de1340ac866a6611f51aca791c7a1b159dc0cd2846401773f675841e17a14fd0245422bbe8979f4e5a8eebb74eb48637d26d496e25ddaa2a23065a270728303bcf0a863abb7b457ee40238caad84619577e44f29b686fe5106bf74bd6468d9d9129dfc8e1225514cb96afd5501c630111f9dd17509f84bcdaa7b5645f77765b6e791b90ee2084bb8e69cb089abe10654d8afecb446015599e5dc10c40a852fbb8a9596934b69c010c73acae3915bd617d42a8717666f9b7fed0567ac3163a2c53652c13268c0de9a2b5b60d3d38e725c427936f08bdfb503ffdd29109513e3a3e45c4733efc31255bbfafcb38da7be77a0a9536709f5dded2c8d9bc321b186808a671157bbf858127099d1b1862706a42820d8e616b4da17b39d3a078eb032700cc0a0d2eef8081dd5c2c065b348d1045b1d813fb8241e5344ec3b9d8d1c0f78f6ebfa02b290aa96c0b4d582419fea160e065ddbf323bb61799029ae74a88f4176cd5a93cf6facd32c8d019613356ec59bc23ef30e8b1b388a46a239c22916e66aec42381dbbf28cbaaebb7917900d37301b2a8e845c9bc38bb06c4a9dcb02dd3fd60f0b4e622e4482e1aa0f897f88b3a4f5abde83d0175ceee170db0eaf042a257bd36236096c48028298aa24f1ea168c74797f80d2d4bbe8d34d13caa21f4d01a2004a56ffc7d9c40e5421d4dc8e1da4a2d5a63ea3c2fb08047cdc3423bc9eb8f35fa3f0aff0875a99784531b41ba956f40ac88f5810a967f972ce537d94d04788f233fa44f88cd2802397491618a8a115f287b64ebb80063d441e6f8369f6a37f0ba1ef86252bc75a3dc76fa107578f3ed2a0ec18968b41fa4ba3f1a839ccf41c8e6a919960c0ee788d75f5ff5181d9fb0caa5fe51dfcaee1736c7050d3ced89fd4d88464b30d0cb0e46cb10721944c8e3da54de59da32213169acda2883b3c58368ada21c9e0015bb3d193e7a431a7c0983da8ccb20a0f4a7f94b39232d350e75509745997b2d502dd9f2913e524f180e63f9c1642c66614fee38469b2109cc52e133b4887dd62cb8cb1f730ab8fdfb178b2a69ff2269350d7ec313998b385116cf011f91cd4df279b7d80dcd62184b134d24b14cc371c7f6e8b3203c1af2e4b4f18ecaa0d5e09dbc3bd50fe70fabe114e8f841215f565976609de77217cc1bee8c0f136824c7d4f6234e4349160bd87a9162595a731d312f1be4d57e78281b4e97528315e89c86dcbcd22fe3fc7880640dddf9d1df400848cfed42532507276799598c9a5ad588caf1166a206bd3ebb92817d53b469b3c332da63311bc3192cdcab4c5f642c6a9f78260157063924d6378d6bacfa78bacc894fcb0f96a299668e4fc718055b95ed7666c041340c9626183946eede2968ab0d8ae265127226310aad30d0b0d5b0de435cfbdb8d91e177e7ed98942c6cc2ff4ccedbaf1a543338011761c96b17557ac71c5ee5a173ca4b1a809edccea4ac02b9f4e440326d105f8a4daa57a823f8c854cb1021b71bab3788f2b23887ef8bc982a6e9fbf21c8e616b932ddcdb9ce42b2c6f1d5b6321a63cda994cfe5ac61ea43f6ab178ca8be3349d32eef41fe87fbbd35e0d91c8bb08c72317e5e1cc987489fe28987241b19bc7be61720bc8a76237d8d70fddc405f1e10853ae8039dc7b58220754095a562342cad1ede35d4ec18be6835473747795306a661912c9d2189080e853e43078c6ca95342f0a9e28362a2369f743ffef22a60bbb4306ddd0377110857c96e1e58d6e89dc3dcfd018414b154f597ed38e84950a082431a3f85b2592aaccd240e9743934cc4863ebcb46f0611db1826f29bc1c13a38bb1179c9cb1e01dd62d8c59a02cc1a1ddf70afb08e1b2ce925aaee210248738d73e3a0b4c9fdcccb77f1d12aa2063a40b8fc0cd859cd0ec866716710266020e1c0bee0cc7769b8600b83176090e4670b1104f81eece2d6131ac0125ab0f94a3b3ee74105c9c99c2512080765b29334db5959a720ec93c67e08921a8d91b02356de390ef49732e2fea5c575b73e1843be0dff4c178b3bfcbd86302d1f8a01d2f838db38c30cddc52855efed50e25c724ae366471aaec698a5dbecd319c24469b650a2ad51bdfa5546689c822f6977802280decb1535d4a051e8d37c93c9ba1e77fdc3b42d00270c0875faf8aae3fc5a186241f32435b780a2c02678f06e34398a013f5567c401496ba63f8bda18e300c5b2f47c884ddd75566b0687e082b2d56b84870f3a3d16a1d649c85e110b437eafae7b13a0f86fbd2193d93f4ba7dcb3b0659bc0d5338cac23d8c76da4bea6e2baaccb4dc1b142138c1f0e172863b748720115c188583fcb199306abf616d267031b1ad49695754af271320bb5cd51c44c0ef77ed7e900ec0c1023f1537bcdfb33f361ea2b1bf4e86893d343d29752c52a9b6817151e4de37789b69960983fc327164ac70eb4781113b258adac06ddf8fe29578bd82778aa8ffa618c022cf568d19ba74d77a3ad21b258be256de85a50cc87bd1c628fb962cf84f8095c87f8b2fe126344f630100be96e291fa5fdb3aa1f4fbf4f81925d90747c9d7185751fc053f47d4cad9123cebecb83f0d7dfdbebbb7d5d35f3c36552a2acc991761c3208d22b46a6f669ae66bf3d307de85ab09b3abc016ba0bab62b4f540e60ec43fc0f4a7cfe3083f46c82a7b5c14ba1ae8b201461dddeea4a23a4229a36e8005fcae6ca852b201217215de643760d1b62346ad8745f652edc63e22c3d0c32186c9767cdd4bc5d3f568b6e357ebb7eb256c4aa630613db1ed66ca16cf188902c7592407a58038beff44f382d06ec8103607f3bd033724ab00591985aceb3cf4667cb8f35dbb15c33fc30b385a63d9cd4b4045bd03cbc095194a4070bfad58c6239ddbc29c3f119026e19ed3feda1959589f87309a2ed21049c2eb494d797286b3968af3b95893236db81cbf22e8ffb6bf6f26610735439b384f5d8b78859a1311069dab52ad32d128d454475b7e29805164d599a47bae817e7b5fd1b9d51f45250a1a683a3fe4a241264b768ea9329331739d989bd55526e7c4910ba8b81af1857afce07ae02ddd4962ad71b7d0c6dd5cbb67fa4e2f85dbd35ff24ca18ed0fad3e283ac1f7a20a4b69b2265c9a79ce5856f24c37a781bdc44ecc996dfb63d42fe9be589fc0725a3899f6eafcdb1aa82244d4ca605c70550b02bdb4240980d53f91334859c2de87568a8b4dc508caa3011a020ba6b20add0184002de2bdff820fd272a5d763d5f88b956fcafb6d9538efeacbb2cce41e2e401923a36bfae0e1f71d48ec7cef365a9c07779503fc78506b1a38d93972d529c5fe7ad70f031fdea2c8a9b878d417e0a5a438471797bfd378c4c43662f00728e59523de6faa0ddc6c6a5b9e8f075d053bcdc3615676b37c80f39fce559832c04e9d7ce6a9becc0bbbb672dfe29e318820cdc2888cbabc6af916c9bb8fd30613507341c294f7b359a4cd79a4d4c1387adb85d7b63df3e87665000c184e9b9e06c0384525b7f92663745a9009bb45e13aa7b4dbf200409babd16362433a2570d6c5cb6f5cfc3cd7f4e75676bde45ac0d55e4fb53eae155bf7d6c6f509cacc582f657a0c82097ec908b8455558ca5836d69291b9ce67f5c0619a9fb6a5d5d659da6069b3ef647ca89467e17eaeef43abb8b62a44723142258db85c3650440ad274e2ebff055786b167a87ef3933a0fdfd5d45f38b6c78706d4868f963309a070faad78975a5d4d1d4e69026427b76c515a055493ee021673d2f8ab8f671efb0e3687dfc22b626e3e1bbb00e235b40178d45c48987cb9c908f7b21f6e1cb221ff97385d7c27a3eda93c1a07a1c310f76378ec02016b075651eb0cd8c73d3ab9e58cd0917b131d9194e87ac8f571de1915c3b4304eb88519077318014e0e298f54508e9b041b755df13d5f7b777575b77f472ac41d1056ae75362dbbd9fd6e6e20b38b824a5090419c5914bf316a5af3382303a0f3c5a57f97ad2e1ae6c3f82054673e85ec4431f1ac1bcdd41aeb339ed23d19e6794673ba3937c32e412098da2120f2daf1541fbae375fca8e46a602eb7bde19c22114914bc46fef13fb387fe3bb895fe4284319e9136f96d6f1d6481535f232bfdb98d908d6ae0f4174509df90ccc1c99ad22cf93ba7ddf1d50f4c25170141256ab6f1ad65658a97e71264958d70adf5c3cb041a06680f104866de08abc088146fa47750636a15b21a7606e27821573ebafcd0c9916bd2759af686fb4558c86ef37dc0ff657264c3ab6ee4f0f8acee45e64e68e9c0526e018e012faac143203323f7c0f040740d0f7ad403c9a7cc5b56c5a144ec289f8be15d334296575548dd43f7cbb3cc2b9b5dd6d8b5641727fea8548f0249bc69058d2e1daf7fb234ad9fd3222552ef7f131c70587d559b2a0b3962ec89392b29453d6ec8d19d024581e8e7204c9fd36914e13e54ee387a3cb4bae7900830e40ef2ef4cfd53347049454b9c265bd34daea5b1e8ba218576e2776fccfbef3a3dcff259409d5bfc765d0895962bf677788a81cd6eda106755a0e52b34e72b48a55f3040b0fb7b36a195c287c67aa3250ea4f3652dee1ab34fbff26bde4887c026f36013d32d04e525fd909f7dea91bbdf408153f780abe8a61c53c15ec3156dcc266a7ae2a35565bbd197ec803bde9f34402c99a82315a041182956d8a88c3085b22f12dc850c83ee9614a3bc88ec1e87ad7e4d6f5e06ab5300244f1bd208ae532d93f03d7a09cbaf9bbaf8e611e96cc9d16dc595861e9bd32cd6fca8215785b04021a77770dd0ee157ad1da3349957f236cbe8bd26ada477f43e311158d010f86cdf749ad358016e5f3aa15973ae92ac2e2c23bde7a2b1806233a2fb7d2b2d74cd4b15eb4665bb44bda2993766816c8ec677b9bc184c33307ea310652c0dd5023d5ece2d70c6026a28df8d28787fab2b4adcdf54bc9dd2f7f0acc9c6a741e55b0a6495d12c7e9b708d73325d65ab895120298d132967242bd7a2a0b191b337285fa95a5d6fe2221768912ce2e8bdaa9d6d4382a315b3d5a52727177c9a6c8acdca3fdea47c5e19a6f499d3d7c167da34a4973325a6e52b81a7a913eff440810ad60c60b9fda3413198bd87022c79ea08297a634ff9fd267a882d914436116390278de5c7b52d8f652b786cf492c102fc6d4d6ad0b57915619348d65f172e062d9aa3c2946badfb88d09ba8182d6900ab0337a789c47b8ad1b6e4ec34ddfca1d4a14c0999a726bbcc287cecaefebc4e5cfd42ce8da457bee68929e103f5a42489947fd5a5181092be9fea6861677db38878be9f81e5be822ec944dfc7626fb548c23e88e4934f511453f60fd279285d16ca780af7e722d5a0059bbc5e96bd2eb0e4ee12d7e4fa8e1cbd02f4df948f8d0bf813e7a33c9066fcc38c90ccf71c18fdbf75af840917f87623450a1b1588ea40874e5b9afe191f079be535f29b33741a3b96c8a1295b69988b36ab7b715c7acd79594bbdde0114a0307a6c8e63beac5b4eef53ff0d7df85010bc5719e4d2207149f637449a6a1f08cb174379986fcc9bdf2e93115efb382f5b8c7944b746d02392a07ff426a0204a14ed;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4d68c7c05320361ebcbd44d526c70e896485c44c4ce1a71b2b64ea14a10c8f50f316436424c84a0847c7c8130a73bdc3de4f17cde746d41c809f3c0fc2430847089f1e3fd6e9c4f81e38eb558de8fecaf25a8420001dece1ed5ecdfd7d23000067cd8d4d9d498277b9169571749b12998ffb823820b852c87d0bf54146d74d64534d625c7da56dfaeeb4444d01e7618ffa623857458abb38ee56ae4cdc0ae19c3781cf3bb39db5aaa7cf7126960df7ef5ea278c84e1dee6cbd469d5dba7e725ca9303e5321f3c57536e42b2a7c0270b044269654427411a8d6d242e41200360e0ffdd98d94ca78dc1a09055e56c1397d6ede00e7244c84d052047a9ffbde53fd811cb873c3907a913e8b5861928f45a5b1d4d4ee1d84e5ef06ece64efe87907da877687cd78b07b6aa77c15fbf08e4af0ac3bc0e165963bd5504e9cafacaf831a9a164fc58dae72368d16b61fd1d3fd0b38f799a5a4a2126a466098c4fa0355ba9e7228012b9dd512a1f83af80f44bd0830f2714c0fba593f9032618da2a0ec5d202c974dc0b2c50c2514fcc2ca67ec8d48f48bfc5a879d211b5857e76922a5e66b68c89c262d0393c0a9d5e349a552eba160bd436e149743c693285fbd32d08d5239ba7fbc2394eeea0c19d8311369d5af85238fef0cc4cf070036847c411bdfd0136ed23bd04294e0af9a81680f68741613de95a511c16ea641b87678b5f3b3720e33985d2bbd77cabb2bb11336508921da685c27e86bf1ccb66cb3e58aa89d5afa072a231578edbf54280010eb7b419607fc3319c77d083752cbe1c14495922a04297245f4954ae87a9c96049cb5d528e3258eec38139e63e123a34476916b97eb2090bb2000496951bbf707d4521f4fccde8d8ce553c17b9d9e41204842d57ca9751b2ad96d7bd8a36d88e333678f92ded10ec5c242f5ecb2482d9b19c070af6f81bcbd5a771d5fdfb2e25be916a3c75e0a2332cabcbb211ded8fbd1ead27523c76f4afe0fe38e13cea79cd6ecf47a843a20a6c13a1357aad9fba402337d7a0da9b56a2649ba8946d81b44952768cd9b894f8ae928f441830919c67c93cc7cdad441bbc6d0d8d2d3ceff0ea06eef7fd552a51925efe6a94175bfe5f4cecc4b3c625c56efdbd50b6b6392e906355f3fdac7f600e47203cfa72b4c61aea88bb92b258292db05c5614165d1a36536f630b0cfb07e0d1f9790d49b660f645adc5ba001dd7fd810a2cf151fb5c478df49f91e5f72e5df1816368f669f1ab6279234d8db423fdd4112c2236b4bc446e9f76afb707c0b5ff79bed5f2d5f14c430f921bcee4ce46e0fe43eccbfc63eb41a623a94d2454a77e489229e3cbe445ed8055f01a78769e53dc3600284bc39f50d33fea1c332b09676929e2d24c59e61f57e9e2901b53c8229c7abb72c94a9aa2ebe23c4a6c43910363baf99873a647fcddad4ec127270b968071f679d1cca8d86f3ca46fb0f7cb9b60f29220295c7dce5323e9914f8b634b636ba977353a6ebc8361063d6740741a9addff826f352c0a9e5f051886fb467b5fd93cca41dcf45368ebd62109b7dc8541b7c5743711d2e41dc33400e59fc1df63cb60bf30d30b1ca5d9c42da5cbf49d44eac28e816a6eb487042bc9e486c26a3e76fee3a663f850358df63e44c7ce0c123208b805f28e55d2fdf65a8372d3c1b328e4d32dacdcc2e29aaa35f8b1c5b5895bf5c50207ee21febdfe80216730f548d43d597991f87ee57b7de10101c7f353a3c5bfc59cf03a6b03c259a745e02d30d6647297846b457897170f48045d04229038e7a6f063a5f838165f3b3dcd669709e927b13eb8b9aabc806e41bb3e567d44119a4f14ea985496dd283fe57140fb29328db6699bba20d997c336cc643eddf13e24e52a3f30b5c7fccc833973f9f2844bc185b77ff4c5ed96743f68653eed2c0d78510907ab7d3c9d9f37724f5a32ff45697f026eed8e44bdd0b96029f6b46e869c3e2f8a12b0939517b8e4153f6040b4c87978e079ac6b8f0f40128996ee4c6af2399fcf18e55e8d3cdd99cc14e65c92da2f1a2088999717d30e28e100dd86d6821df7f01054ffbe268c453adb66126b82aa689a601f57d393ee36207681eacfc47500d5e4b28de56d1ddc0831ee05f3914677a907e179e4fe8f597051f4baa18530d01232c006b1d34d53e2cf7ba159a1d7d54cc9a25d44e5aaf1f6f10322e3acc5abf2d66cb4fb0205a50b35bc6ea00be81144940d6a7cec4e18ed6630969900909bb8e4139ca843e4ccd15b85cdc9d97a72d5a46d3532b335fe99d1ce61672955e3cb088f4f4938df9a5224fd019b97dfebc8c07fda8573a97eba2e0fdfab4aa5f3e102ae1e68bfc96359155ffa8518564c9bedfa93834e497c4c3bbff0740a14f711c40faff1294cfc78ab59acec89d1e1e4877dd57e5a1f664667b625dc94a398189a826b12039e3d410aa2b9fe874d672f2a68f2054422810bb97bde7a90cb7cdd06d4bb5813a1294a39f8624a269740c36e130c85bb1798c156994592517d0fbb24e3b42ab86bfaaa9afe5abc90920323653e292006bfb001bf107d5c1700a77fdfed228da86de9993cfd5bca28bc143635a8ced58719ce1e6c49410cdc9f7ce96eb06abe70effcfc321c602052c184c3efcf6224d58221b6c555cef232130169758e1372cf223d6348f2790e87401f74eb8669afa8148ed835aec2b530f2ab865aed271e630d6649e38da996353031c145c0c38e58386afbade1f847be01ddc61ea6e93ad94952f9d630a6f3f8c9bab566d3276b2db6bceb542b116ea41a94eebd5bdf08c3ac7956fc1cca58cdddeca1197869baeeb797f32fae9b952fb99975bc0887671d9fcd25c0914b422ab34bb800a3c383388b0e9a31855819c4b8be80a6c1bf05977760ad9dec3d2da5a8e5e1f51dd4644f95f111174269869b48510f69634b7d722872b9110023e48c04ce659c4d135d21ee92bde11182d11aea70d155a64704267f8444d89fcf655ebfbdafe08aab99c9b1a133be285032ea9c2f044fd75c833a61b6675a724376066facbb303800d9dedd60de56ed1b88d0085a91edfe3dae6d8635ef2fd1eff1e2e267c761a805b2473087160ad106718037b27bd596db58557ba5f4389659a3e0692234614946416af035b2a7c25699dcb10c1f91dff1e1f22136adf57c2c4d6ff12e928874bbd337b9b2795de5bbd01b1a123d4b85f3ea72ffc799e11dec253f0332b7cbd074c79c8f765cdbb512795b684cf2fd499eadad4a453a7af3a5c94d9621d873d727cacb8f2661b96c6af5224446ade1d81ca715419d9874c7c3b8b8f07bf1fd4e1b3b4d56bbc2f5989e0d158eba24e5f070e51068e1c6e094126b6537a69d1ac1fa34adb52aceea554bafd62bd34726a965623edfbfc4908e3382b764925cd4d4c96902db203ff873b0ac5cdcb316aebf8985d663df6d73ba2cecffcfb63706d418dcd74bc80fd1c26f47a70d293ee957b0c11b088d04290a3b1ad56d4d8e883f89e90f12d26eef2a507b547a11a4466e8deb6b704b064c0e78f3031ac6f23eb03ed0dfcd12d4395340c864f6c1c9dda696f549df356b1dbd2517e234119b8ffe5a0337a0ba596cc412479aa49779271489cd8e40761651c00ddc1708c5de1f0cb14a5c91a57821fe8d70fd53388260bcefead5a98c5249fccdde7923e2aee633c7b02ce1f26987c603bc2f14a301fd2b91a7bf905bb38a15f33d31630eec4f637cf0751c93f8271246437675c61c1eecd252c3e883f614609d4dc316762a26e50b63f4dbcdd89e920a50a5b8ad34d35c163aa54ecf5d57f13fd7deb65d9a81c6c2ed3d75e2dc2ff34a54413c10de9db6f5833f5c97ef1afbdfa90d394caf33e9befb01d2526015460aff6a152ec0c780a2e6759dae38bf3d3af1061a03f3c3a4790a6be6827996ef65fc618493dac0a9cbb313031b21ae6965d93e4d1dd4c401ba357af48d7147eddf407b6cce9dc35203f0f64a64f5ce537d4a10a193dd506e6618477e05216a7a6cdd445405b7ed2e49730e40b24f82fc77ec3bf6158831c87eeaa74a50c321636e9580b274e3df267abf49bff3d8c96087f6dcf7755a338964bb7808998e413636677db31a0d8c939c15b49f3baf3420897a2a2ac34a912db2547274970e56ac92f65d55b7464ca1710aa7189031099a303a13e916c681d9fdd45402115ba2e3049c96ea1e5cd7a1661e17325bf0204c4fb0c707d27a0e849f2689aabf265f8057c53812e8e483efe99fd5e50ed501960184a927f0281eee4fa86f4baeeffe1f4f15e761df3cf35e419569a2bd0bd42ff513c1fb86505ac7a17165552ad591f84f58bd4585f09841655155f8a2044fd6d02f83ded5b632842f219a71722aef3c09b9643389f29bf81c1a121f5e9c3c043b99d3d9f5182d5cca099480f9f90d4139418447b8c7f6ae79e934c2427bba5da73b4fb3fd338b86b2e05bb8e61ca3b4749ef473d0dbe7cb82eb30b93b1683b121a017850ecc0b9e95dbd29b5a4e81ab0b1ee67b660f595f828a1552806b857f9649a2ca1ca32ceaca72c76a541fd4cecf03df54752fca0fd0f95d6948091d80876fd63c15a5f600f77dff90309d100a3967bff4a64db064736d574c0d4a737325d6e3779a60e63d8ab996c3c6915beeaace400034cb4ca1456536345302fdaff96e933037de6df70e5db8447f935bb59b0b1233505aa7a0ecf87cc6ec6649c2f824d6764c7572993280e464e87d1309c2d30a0feb915ccd4098da194a6b4856f72666a16f84affd6789d00cfd90c7ab6ef32571644f4fb99bde4b645c153a7d0d207973811241f05368d3df87b86bb010e1d80c52faec316c07f1a66d2bb560ca2da70b3ab82e1667894cb939ea7a365860de114548373ce4eba76391fa0410cd609d77c1fa4fdc7cecfa20def43a899b4381226bcf1e2a98696d194029cbeccadfc032b73cfd81c6d1f8175fdcb8430bfe095d70723dada692c18746acef4dbe0bd629ad356f50507118b692a1efae75a0680a39016a4f69be3879225c9d9b5401e232a6cdad861ce2377baeb154bf186945af4241cd2f5cf238837564695073a2d3daf4948ddfad80cc20274f4bd72ffd795a3f983c0d981cabcfd60d0304361a35ad38e61a4b3e40da0fbb2dd98768c24ce6c3e6cc4734423f25bc3978b89fcdf217bb0e6b603c9b379be0f4c5e7756b08faeded4db6657ccf233af349c00785756e646fd28a8ba6feedff71beb77ee004d68a21725e5617632a96c3e7ac03bdcb40818c3fc3685ef5f9ef51a54aa66a1b78dab7e90ee0ce50cd381905be6b8107d812ad448c4afdb53f805e70b25b84059490ab15dc3f123a853d25f9469e6e0dfc21698f3855d55e5aa1b9650e1dff2c392b0540d9880a189cacb83db667effc605e39f98110ba0c94df4e069076e4aa00ead68bfd85eca98c190ee303d3d0eb25194e32e32b05f6131a758a7fd141cc952d245e330ecb6a3db855310c9a43bac61d4e4194cf40d4564b04203c77279c852c374e6cef6c5d431d90941595c1d2928df97067224f5ada0f1fe472176d8f42f84e510bc427962b9e29aaf44e6f37a34534d68920ef01730fd516ef996959e874cc5001e7d67d4df7facc536883b0421d0e778e580a2ba6251c35a5f776126b31fc5b09e4c108ca8f545dc0a61430ec21d6a96d26a904fe448b67515b91e8b5408f3ddb02b5ecc38a4f8633a8c841f8613aee38060aed27395f56321aefe77408cb55f446862a8cd483677b2ebe4b5683e689ddec8a6409100e88f8eb8a10ccef9ce87ad;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h932c8f579041bf774442b296f225a919c3aeae3991b8499edab30f6737fd8e8929d7e42e1ba232b4e1ecfa72e71b803f48c6bea017de305034225a76c0a96457f1c27ce64b2f2903266fd52dd4ee42390194ee7638634491a5efdfdaebe68ecc6dcd152b4ac4615d593c9b33cbb62776c886b559f13ef0a9904fc363a7476a96f27fc0960de7e58017b46d33cc227ac048c85a69a31d7e9a80f0fa44379571cebe5f33deaf79140e8de2e17cb64ca3d9148af2db2cdaac590da8440958073809a9832dc96a77d1e076fef3f56dc9476560aa041ca38e14e57de73a565d5f3d94e9ae11aed1943f51ffc476c5b36a9c6a3ee54991808db9dc8cf126c822b596dcee3a896e57b50d917ddaefed7928beee4f4fe6c2e14fc60b913cecc1249ca0aedd91aed53490314ae138a29b7e02d6cb91d3f33fa45311ffa525e0142a35bb3a0e37a0ba5e58b8e4bd0756178dad596a26c2906becbfc3cbbbb1188c55586f7d86f7feda51bffe94c26624eb3f0fe06bbab0303e5299833d60d3e5ffa06ebc936a220f7925934291f4f80b6db12fd077ac7fd28d87f96c2e71da22e14bfb0af4f0e5964e8d28bc4be2374eda0ff9cabb96b64455db4b1107aec83a7424e845f7648d17ba674db94de37807abf706b16e50db5bd6a72b3e227c7ead53902bd4eb5612981fd8f01fc7d8b5a5920fd980882972269a89472f04c3d709e9d755a8a37ed9507002771e2fffcf58b638a57088e95f414dc8546d69ecd314a13c741012a97baa9c6c581e116fd2175009c329fdc52133895050aeb030ae01ce3c4f2ec4fd77f327e4489e07484068d3790631e7257a06ee4f4129ed034a0e1bdac35c71bdf835e4f331d81db5b9efaaf3d41ef530fbd52d6ed7e9ca9db902ef66e8aec66084c3fea1f69088e5cc4bd0bbabb223b185760ade369920348c9f964a41306fce52e722ff79c26146a093c0052e2f6de0ec6d4bcc966295ad5d5760ad56ef4a8d3e94d3b4c629e5feb68c4d628cdbdb0881a53703fc7955cb53fce54405c1c2c0016a67e2ae098978946b27b21f8329ed18c3cef99c3ba7a1bc0d18d11bafb6bcb020c218b32225c7d074f93d74c1fc359ab5428bb0616c2c343a9ac97ef2b9113ecdb46ba4001b159607a3c5061a309ee98d37850d00be6b95e4b30f2dbde0dd18e028dd5650329dd8363655a839b9d29f081f472290adb863b8be8722c2d4e9570ecc7fa3a5eb817ef8e13b53d4efb93202e1c1ac0963cd1dc5c1de5408fbea4000f608bd16b5de7a113d02457d93722a138bbe2fed93c37d7343fe1506c0cba562de5377fd9f12a2f947c08e19b98b437c63b1c8789c475b6df3b3be4900d50988b98ddbb7a60e90bd0ed18dafb58683574dc0a8a080676f98d8371a69ea03ffac56ade053788683adb9af4ef28e4a6c819252b104c2a41c23b66756ebca7d0b55b3f1631825ed23e072ecca43ba5af565f69b712a8b9faf6eaaa5189fa005643ff6d217285476d086be508bce7ea4d59a36b7647fd1b59c8f8d30ffe3cea25c09a2894524d9d7b732c2cab11304d88944c851d6d7e812473885b10b3e5ffe99ac4f95cae5fa3d82b38db9c494f77ac24bf2b94f8d6284db3b84ee6a3a20866ceb17e4f05e310528c70f62400921a6817d73ea675c0d69bc000624d33f5ff325f8c995eae2a1711ce39381e00ccfff4a94b2bdcd52d25a38e42a691066cfeebcd1353977388612e99002868c44821988c0c67a20b2604a31d1b14f4ad9a9c47bbbdbb406da59fe406664e55eba1c0ab0c931c060f2462bcd33fca390388baf6a6e99b214871308415fe8f998d18ff401d41e416039236f409976a8031c3caf4ff261ffc9f655a76ce88c53bfc80778cecebca6e44530570d808a201289510e280ebc0dda25a828c1286233d8a25421fd29aa20e2c370729bf2256d953677c1a8baf208eb4587b597ce0a258adde6d00f793bb48b4769c9c799434f0331c252940fe2b0c2d3f2f0a326ffe45d9d69c3433ed911809819eff2a7f14fe66017416c9db66fd7f9fd684a191985fad459146f4f904c577727bee663cf89a9c420289c1d590350a5ecb6c709a6b0d2d83728c28b6cbf86a54afc3252aa2016a1d3e4900c33ffc4139fad6c87754ee75b51d87de7fd05905359522973eaed8dc6c52ad8748bf63d19155b22581b7bf505a0c8bdc9d313e4bf17ccd335fc86876f0bd40f9ae0d11d4598224093a6578df5b607615927a823df31654aa61bbfe33f83aea09760db6b236752a5f2765c6c020a6a071d7eba448a1bbce6f601dcd9965fe43c060e6fc6b1c83ce4e3af91661aa374d6c91ff82a197565fbc921d0c77e14b326b3f91383610b2022089d76ca5b9127a1f294882b364241209c7f26ecb18e26c630383071995ed5c9bea45227053352f3ba7eab46ace37d0e7eb335f9111e28761b27db1daf8ae3e090779e6e96c28aaa1be2e926de876f1ef4b099c728c69279b478a7bf87ce71880198c6d01e0f6b3f0d75a38fdb694bf2a0ab6e6d2be1990d1c5af9b757015700649a13ca323033714c8992bad2895e86a10cbd89772e9e3280c875b6a584fa2673c2fc8c5ee75e5cc281804e76787eff821a0bf128c65af50d8fcc9d6992b5a915802bb8043d51788773fe8689ad7994bb920b39f88d98134af6883cb6919e78c363ddfd19d900b0adbae3652583c58b641a3d8ebd5c144fa99fb6adbd32412b4be2534e152686d81f17dd879226e56edd24536c8f5cdd7ef07491b0255683a4ae7cea64df1c537ba1b21bc244118ded801357df249da53b51f6a1522c648dc5feeb57ff72a4d48f4b23bfc23bce945011668df5f82a5ecc8e6874e1fa5862f66d1f3939063ab7f58aa59cef17613f9ded3cc4a02d05cb02bd38205fb68818fde430cec593601c897ec7ed0bdb609b48267843cb6e002a2ef62b62338155724d53f0a47bd3ac981de12a7658c2fa8aca5541d91e2b16d93d34f2f2775c80c62f6e521f437a495bfadbf5a53edf7425e1e8c6a6f81b115bfded9d3aaab8d03f4a1ffec76eb3002141065d0009e0392fc8983c8eb961ef8a7f04f83022df3bd1a95afb908d310fe730558e549437374e2444c619e2522e0967f7e0f5ebf4bc7a31bf024032477cee3a76cfcc33dd80f539de36bc8fca66bda17ca737b8f96d3ea73fa529ee460c0b2368d27d9954c7b6c75ab6f280d570d3455605625834804ecaa82f708a5173d8a91f838d978062fd83c12a12cd00214168e99ba7abdaf42f680f98fcd6cdb037c5439ab4dfb99435c2428ab814d72dfe975225bbfbdb60dd11b86763043c08f1cee8de5c65275d22199ed9ac95a8ae2a636b46fe1a277d542ac0135e4750ff22ff6191fd7f43cea64122d081dedcaae40acbef5b92b529a250412b844252ef13e04e7bbb5ecd5d6cc01eada3238cc64616cdd325f49c42a23daf65638aeb57c29eda63b7ef3c170dffd702902d19585a1ce19b67ac16422b0d6c847607e3434243f6a9b19e59da3cb3c5a45a2e42255c815dec3853343bda1ef10df9660164268c31aca75581c7d916d2f65337da4fa73c9790b78f632d22d95b0e5b089dac2ca34311134a4a9d1ac1801ed168a148737b44876486999896f7483e0e74cff0f34dd093997c798f43512b9fd67479058146e3880f4d2b7662a96f6c0ea169f4defda8102672659564b2b3449a484d83dd73ae389c22e79baac62222cd19f7bd20c02b55a8a0ed69edc837a299da58ce9c380ebbe15110cdc173aa0ff34167d3b0e0199fa514c112f225aed4a6678709f6b83e1269a612c790ae672d6798aeb0387259d1fc5ab4cadd06520ed9f0b4e9c51d9cb868b74f27e9a60fffef582673dd50623371aea099f69dde5dd0f2c08d6b05cb8c7316d8c8b39510fe5237e8791aa82a1acb9f9e5e537f0276a2c540bd0c1844093c28d270772d620696e7b2b8c0e8064a45c36cfd34b5afa19bd6db4bc0c2319c70a26ec63fe226120b000580a78f0fb212d4dd57558e095c52bde7e4326c2c57bab2c96612f4e9e03e7f08f7aa0c34205af1001571f89d8d9949cae3a88b0475f58f48206eb47c18eba30f354c9c3af08743ffb028a36113d5b9a0c28821548655b8fad2a907f94acbf5da2606c354e4740c6b33bc0f8a2ee255c3e3ecaff23c7f9d4e9d06f18ef7bf597b21f20376e15e38ee7f96d1eb3a30fe25801f088dc5205d0b7e8eb758a72111b65ea7477467007157a06bde57a65d7578acbfe6358f4754bcbecbd35f2d28d588ce0806d5302636e82598681e12e2b6b267993631d4af8f0bdce2f08c4a18bbc4b998f3a709cdb658c457b3bd7fcab6bbdef14bda525b06fd02849fc6342f08461ddba802bed4be536149629795fadb8bc089d99803f18f6491640990503e4877f822095287b861d43de4cc827e56a1162d115a0bc5a28d7339ba219b8a5c907f27963c6d13eb1d9613cf086ac2a5182301faa257ba0ea23c8b35a0a7247a337c894cf2d2df2de5317eb671cb0f80ee0fb3dffbf9bb9aee62ee20731f0e095d17b8e4adfcef4412d195a62680a28f26f3f3062ea08855a04892b58bc01244e43ef1e365fd3909721b649f449308329fb5af82a16fc3ce665092b7aa3ac6e03ca92d08507f06bf3f37e43099c955f3e34d7a4f6c2829b7b5d405dc80a3a3ccd937ec68e35b2408ba5718a6cea4fbcb5a4db8d685416d34976cb8139a403c4ff99ff338242e0f041a7308183319c04d0c070789914016483517f7ee2e83d21c9f0e1bf882a9021e5fd243b0ec80539f509e9c6852f80bc12672529d599b0846ce76a867428be932d0684d3abb8fa1d6f025db27222160451ea55c8cbe93423b8ceef11fd523df51f8c95e574d4d4b66f834fdb27939f60b89d23c0771bf8d563fa6d3a65f89274599404fd2f2078c55db9a6883507a6a344fec95365fb4dde4112afa5c3cef59187f1a4fc609516dfd2dcad1108d8a0913f00187009f4ac95ea86da08d13cdbc76a076df94daa6d0e1f8c7398ac22bd9c5bbe9b88abce0c72c99e6f4e539bfbc4ee7848ca18aa735c34cd60f4de86aeb0d3ab46c4f6f817ca855406f0b66f4d47ffaba058ba7b58439cd204921ad74d8e05d12797189164a33ad1626e7d54a748fb1c237e238ad767c1971af0f4db5101a07cadd0bcebbc58c24d6ca17830188f01f8be635f7947e7f6db3ac7fecec17c843a873a244de1912eabacbf798dbde4f530f27f2fb4b883fdec1639c6b00ba63bbbd7ae0012abf2f1b685115074346b32766d517c3625e86d3481af1d87ccf688a412e031b43df4da8bbc173976d979c44a8fb10ef60552310431aeeba071561d00da016acb5f464ef2b2ae21943831246f251f5d4c383bebdf0aa4ba1f9a55c5413a315df8944f0e89d2f2cac3726a7a3436fea20e2a8a15c6bd5cab66b2505e5c20d3108fd9a4d2b02c104d4a99f001794aed8927329c0cdf6a1ace0e710f80cd6d35e2c8817c2da0963bb7ee059cc73c8d6690575d29be7377db9e364ab0abd6e47c21f678f014b4f91618382922617aa31b4579d8f481603df87c66d3abca08237ce0deee1ffa5ade9a0c7a8fa9d97e46c4b43c4e456a6a508cb59b87b60222b85f126625d4adce8b58c7a9113006c145f621171d723fc6d2f5447d2d8cad76eee072d0932207368d7467085d83105337e0bbbdde4fcbdacbe4d5dd5eb831025bac2518ed412bba2715c011ff73d7efc9ddfa80fb11e2767d8f11c9298a417ff92fe90331e7badb45a5db1198692922ffa7c88a252835d563d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha59cb5907be8190dc74fa73c1a71044d9d2ac4dd7e8d456363c80e775425b65a62e879c170e889b8c3fc6077d788a7925c1167c1bc92c5a8fa5d9c9fdfe947fccfe6028504c28085bd4d666d5489cd7e7c7c4bd3343dd61665ba5fb66bec70f3171183b20e3bb89fe76b139ee5d1ab59cf9b01cab98d03048b6a5a127afe11c9b799961aa4a53a5ebdd8924f4947faf36d4b4259fcc98e5b3646701edca9adff643f52292a67ed788eff6338371bd836a2cd134d3cfb80fe18f3dae84cbd7b8711f86bb4ef756d354176eaeefbd8b3fe114d3274cb2c45018df59c7fc02a69693783d3e2175fb97dd4622f9f1367c71399b810063242279bb8c2386497c73008475d513ad6cbccc7690ca5660c9bce16eeabc297eff5ecd3b9008dab3a7608b0601ea2c98f749a7d95ccbf31181c63cdcdfa05347065fa771a767d58027e638c261eadf34ec17f249bd090b098b1a89ffafa8aff8c6d156e156aaaab3d49f22ba8cbfd7e98b21c376128bf00cdd333d7a09a40cdbbaff1e8fec8086901100fc651e8458fa538fd6a9db44fc0c926dfdbc57fea029c8c547fe027bb2165c231b020afb53df7e97d9cd0e8e9fe4b1d2617d006915b6f51b22f99ff467f4c5b623ba9862c5033ac6ccd8ea0d6e8d021e5d0ef6475c8a1c0da6a96cc3b2b1331d9e71a1f309319184646cb4362c273f11a0d93d667066d944e9106c4dd8f85442c26f5752b8e96827dcbf081c2e47fc875c9ba2473234084cf83efa92379e4c25c096ddbea1275f5a6196d860076b9d9b619cbaaca2dbe3789f11872a05fadc9eba92d89f2d0023ebcb29645dfb9120699692315f202871415ff74f733cb7f466228dcc467189970a29a7ae294dc516f55fb550ba381eb75013265973cc5a7b521f8f640f9fa2f752c334c7ce12af79e91be6fb029a7196fedfef6cc8bd21a1f9c7c76b39852ade59191ccdf5de38dd1682706484896c6304f25a5d7bf540b5608ce6bfada382e9e697bc10714854c8c783c17d6f212bfe11ec7f773a565bb338128c09beb42a1355be27fcc342c2e5dfcac343e3af6bd6d53df5b6dc5c05f7a8471bff52d88d8bf2b7c9acbbe06d7d9175196af559b3b770da122d8847e78ce33cd54e803ba4113cadc9d9514ed2e56746665c429794d9b3709980a0ff91ef814120344c284610eccdefbf28af76063a7266b2a1532f01eb2ea3ef06b1a6793a1fdc997d565a5dc72cfd69f68f10dadb3606362564c6e35b0a8cd63a9cae8753265fb5358f5b406fce508755535fcb7092029f82331311d1a46acbc263a87406a3200351e82ad3df39f6d8277f30ce045b25ef789ee28daafa475925d047c58daf7db5f140c9b5a790d8870bfde3155231b5af7c94381fb1b5dd142bccb3c9a8ee6f7266ffa4a47d8991b2ee64e10c328514575cb514611403c10058b9a12415f3983c4680b82a390fad091509729263ba5656b1033aa25f779e1120324423abaf8c8a053ee57e493df6f362649516c823b20b4f92282e4cd9e3038bc17f9de98deb4a8e1da56310c9ae6647f57510d8ad859aaab7ced22f15b3c372384117ca9e0fc5f64c0d89aed733aadce6232c5f4477c39095b41a002de63cb047d520116309374d11536ee8b380a5c823d974e9197c81ddbca41e8b7f80501ec9b3c5266c3c408580fbd6b29e77d3f152a2e6bcaee751df9324aafb35a703b48a1b95117a45b5af1a53351848d04cc260480b93269e48b9b96a4db956b772ecf78663c5364cff93f52fcbd0e1287be9a79a22486eac2777610096d0ef68fb116beb13bd76c16a852d1fa1e1652fbbe5e3ea1d0039d8b9b66558ee901e7df83adff5a0465c969db87e7ec9cd3d3f07aea978a7a3981224afc84f79cfb9b07f9a67f37104532a839998b7734246c951356f3f408ab440199949e718994026d6642229ace7bbb839378f0cbb56b7de1805a2e3613435c89fb1bef29146583400efa499c3e80ce3b81f2d3c1d26b22d0b2eec1f25e683bdc4c57fc3cbbdf2ddf21d16100135ed16c20d2b90d9249bb94a531d00e119936b8fd803650a9a64cba1abc9ca8c73c8c1ba8bbcd883768f7d312cde677e8f6f4729f9e7829eb2da0b5356fcdd9458b0851577e23a665f39c591f6257d12c189c6e4caaceaf1c2be672ac6f681863ab6dfaa1a5a274e5e285ee13404be6f4193d0954338d2792fee339f317b32dd680bc244ba2a285b3f60856725d60479e2d6ddae1e92b6758e1ced1714439c5488b0036f9516acd1785ac69fa476f3d308063b9dcff941a2fa48075e878e9079d20266cb7f10f6fdbc201002c9e3118cbd2c3b7cb45c010cf9471382116c8fd4c925874825e633fcc6a6239d0f78df617b3aa2ba0f2d78c119a8d867bc3904741683908d63176ecf2f001d02b6790eb1423d1aa78457c62cf6ff27f5d2a35c75e80062087bd45f500c5c0ea78ba0bffe6d68d72c0e39b5fe94005b9a563afcf904b8a86896228a1334aa611f6f9fc9855fbbdcdaaa673ebda3aa4bb13e6f90107e18149079ca0f320ece3f24b50073d462d43e2def78f1802fa66f1565858606b114c761458143418cadf51ee25bae27ef1e161402f8e4ecfa3a4ee47fa0a54ea90ea9690d81cf59b7093eaf2c9d513feade552061e53f87e92c80f0ef52e071b73349c70260021d6488cb71109cdaffd952b34f499b0c94741532cc7f76f1c20a0451125d5c7acbbf35de0d57e26cf2b94a28a1d83e621b61a8e3954225004a591d36ae434f787957372fe6c772fe8176e06e33a53859ff6b420081e311299d412802703bcaa169e97addbec84ea2fca2978ac68056fe7c523ea68609b0dff27983a4ecf728e1924ca2835560da5075bd65210d3fab9a3ab44cf1c65506f60b6f35ae9c60c439c727a15be21c168bda15d91648be9ae73232810195468f3403b13603eabdbd07ffd44b5ddb4b89a14fbd99d35e19496856082ba94f48d7348f6807d2848f92876f7d1ec6a1ef95a631ac6c791cc0123b2f4b223debfd8e45961b17cb8a240600ae4155c8ae11e17822e3d83690000b414e19f309c70e1d1e1f56657eff1100db0c0d4cdecb9aff166bc8d3faabfff19f459f133b4bc029d5bf9d6c704ce6739ad9d68db6368292bd7437736ff3b9ec4f862879645882a1ea88bd772fbd4f0e263b0b03dfd3005eddfe272906b2422d560f59df5c72d52522b174eae083078125baebb3d1a58abde2724f621b0958d772daddf0bc4b1c47df6f002c4fc7509c2b788ceb0e7508c0ab506e3c20c68b79bbdef4f7bdcfa146e3c0493a79b9b9a8baff3bed2966d74e3304d2cb42e95ce88ba1be29a5260f0244e26d71049c041e241eccb069a4c1732fdcd32122b3207b84d0488f76110b8fc93cbbfe5ef6a81d92bfb80ede10a85f801ca2b27ad116c2d7e02dcd5b1bcf813561ac27b5fe69e3f4242618bfd13a16b79d8108e0be09fe02272bfbe133df5c7b1c527b83de9bdfed0cb48d75df261bf3203fd01533f395d373394d1283222137439b27beabfbc4daf1ca3082e9ed42ff0759df7b44d0d1fde3f7a25b81b7186de136af4f55918e7e380abc77c82c892f3f7763427fe2942f20ef73662a060b2cb703cb8ecf04c2ba77737f411f385609595877d006938cf3eafc68a67ee66734a17d52af0c70499bc3f43e49249ceedbf14fd4e772acf7157cd1e46d7d9c06f1e2f032a907569b322068092a65e2f00a50f36b97a5d9448f74e80130a3cfe3efeb1c7204dfcd4225753ee948f59e2176ab1f302bbb6980c7434371bd3840aac76ec4d8b272647a70e2fa159883f608c556fbaea8b1ee3fd4e28082485e6db3e66b8a446ff3311324fa3d118b38d53694cedc19871bbe26903cb72dd61a1e1ceb1288f8a4957e83668bd6bf3908a0e7555bdde3aa5fa95aa2a06713eabda7a6644c45c45c1b1b954aa930d508f59c30f2dbbcd0913e29f438dd43f5e0560a9913bf9d119f876e14e99caab40e47a811e401024431f942bd68ae7d7a05bc3933dcfc709bcc7ec5a5650de43ea3c8776d0b828238b711374351a11518b9c1d49b254fb9a946f224a744d4d15a09005a10851b0b655435784ce741a12bedd6e615b1ab4a02d98333eec96e4aa486fee8f4a2e1578dd198e489f60a1e9f85169e87d6478a962924117adc1c189a2781d2c413b7fd27f60c946afb10dc9403a9791ee80937a2e9481a4113f3dc37447b290893c5096e2a6d9393828756ccd5e004126cc3f2fe2cdbcc2e6bd9231ea8dd5a8d09a17b8e90e69df2ef78db2e917fe26fe8af62711c26f90d33b58ce27c8f1b4444456d4f29b17a860a123c8bbe21a32f56579e7b43524920caeac015c73d8a935b51d5b6833699bd09693bf42639901a6e4fa3a43fb924e5349daa4efb564aa1e4735f7b2a559099c3ef9a30766854706c453124174e3604770da2452604a82acfd08ad5514881489ab0e6948ecae7fb7dbdc578da94578b48257c58ca6226d65b5639975823e9d7531ac85fb5ab5d1aaab4cdc807ddca11a3dcb496dba37d88698c1a87c7cd6539d121ecc9a00b7da823cc3628817c748d8e94c37fba7e4ee1c65f7de992b383640b129cb5e42d1f50b94df6702c9f0f3366548e22821d9a0a5abb7034c9f4b9f3ebc90d14f4abe8ee635fc82d66cfd0b4afedb9cb6ed963e476fb941dd2d40c155219b511191cdbb019d13b315e6bedc4283e07403e5b1241d1042793c070e1b9f9ece632b0325706bff5f81945a69aa594369c9c15ea9b6d5e51854fd04b7e937d9edf91a30c4aceb48ec29dc73e8f9c380813cbc8835e51e5a6dacbaddb5635e79b220e7f40909d6d703eb223a91dab817685f4002db9f1584a8152c4bda88a2056168e0559b93651e74328dce30109e3cacfc80ca35a24a31a15ef16d4fb73eeaccabe59cef25a917a6dc34e0e284b39e11030b256071b4631e23c4092b30a7a5c30d329e85c547d15e1a60c409c377ff9de0d5b4cb1c72d80f1625fbed6306e75bfaaab57849c9763d54162be25a318579a46df0a6e45133cb7d8798b53ca4a2aeff8d949bd745b1ef8a8f8ea3cd7dbe31a4b4a0809d3cfeda6b7c47420e9f83ac6aa98dffb2e1379fc641f1eaaf4b5275a5c4b3d290662b79d29a364fa709152004c5d682de92b86f917978871aadce3e4a7869d02ea3b908bb1725aa161b6bea05cb65f9f5bfd18df53f4c249dbcd80d660df5f7b61a28c5344871b791695c20bfe77f43020bede23b9c8c83f0b3726a25dba425db90bb67d66b418446d9f03487b2e69e952feeaeb86282863e336067a23695613d9658316751c1f745d6728ecfee97fc8384671096015f126d115eabbec345f5a1d8e38fbbf758884d8cdd08c4967e44a36200102e78e700503cf7d6607a5ef1d76931673fc65d0eec95ed86754065454d6d5cf8f076384b57fa9cd05358fa56ed386038c9bae10da63efd9e9cafb75d8dd68ee0f75381d470638e316551794e035255de71a5dde97f5b6ff7725fab42956f4a3ec76e1c24e835c9172e1e23601fa11ede5536c3cde13cf2b1bb30043437d612b9c4820409ece6edfdebb5042f940402964585535444afb67e5cd0c42e6733704e5d0d0ab764a2500c412b42a235459aa4dd3938cb6c801e0f8524de5c5551e70f7b9684e17361b98f81e9dcdfed6116d868776ed008e88f90fed5713943e97402a776993a4306bdfcbcb63078449c26258f39b670a51bfb1ade92d923c65cfaa758d8fccc5bcc5343d693e9dc025d06c2027c6b537eb2264231d79a61543f1e23c775;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha3203795f9974884ff24d4423942199076940b70999e39550dc671afb2ec0a59092337c1664b0a08571bba6a648fc0088c69ebfbaeb5079ed6c7d5ce132a9bfe6b39875a62da41d0735e46addf03c18c66e6a751bd478f3d4f25b5fd641f1b245d4cd43f506d7aaac601f55f9fe74441bd72223cbb93ee41a5ca0601001d780393ab5a28cb57dacde94a1a3693fbb1e3708f7a2799b3dcd6f0b954fd2a854083733fd4070beb9d4b9b9e0deb0aca9d93fe0a1895ddd53863f913084f81d04a4421ab2cfca7a5eaeba3131b629dcd96cb9a50acb34550412e323e76f8025f6153277d45dcc59791734d5a8379cec29fed4144ca07c34c8ac1083b76851adccab58f41c2d082db2a947bb8f484b9712430e856e63ba43dd80ea0274c5ecf4cfcef8c4883bde98140ddc1302780cb832561b66d077890b0cb3fadcb55e7c5970de63ce9ebf7d117d0f29429175e272cc48adc614b4bc90f5bbaa9a9e1bea5baa796116b856c87befd00cf3c4d97947dd2e6630be6c39d2faeae1e8be6e3cfeb5ec6c22e3a20f44f6a6e2abd519ba0dd2da77df10d47fc2fa7db481bc26c7acf6ba7bd1c06da767167253669d5ca1f8e322a03ce82a0c612bcd691f696f8536a972e40a52fc4847e2789de95a232e82b6622d28e921bca9f6ba943619d9116fdead84cb510628f98b6dcdb170f6aea771cb540954def3e1dc330c44766829f5a9d5c33ff32a42ba2c6dc5877b12fa07fcf1d4fbf35b65861c2958f55bb8c0d99f7d32dde195f8984554d497428b954eed9e036716b031c26b99eb8e319126d5ae940f4ca132afac68b8d4a4c9d25d71fd11d96550cde808e394ec5aaabfaf3cf6315d0b4979cdd2fcc412d9e58e1eed5ee3259779d1d1204e8f83c87e28286eacb36dd12f37a37f8f5a30061ae6744b3635ba1ee138c33a8c90702fa64bda98d3b7458736bf2a010afdb193e3b4b77606eadbf9358ce1fa4fd173b256d2f89bc7165ba6464199cb795fd1f48142b48e8cb272d59d0c4fee8c6d09ac0b26cfcd05c2c70e5fa076aff46b7ebbeb35289d34ffe0fc1a420d0d23a5444de6decb73f1ed9447f1da7d340213cc4491b4bf09c8f526a71c2d51da5e508920c77f6420acb7f5e6ca26eeed12109d9d20caf730d1d9fd8142677dfe35ca6a36136039cf117de75945d76f6748c519b53245cad0e7020192a2903c20b16608dbaec7b2447aa481b14b9113a33dbc600c4035bb0cdd708d14aa138c34e04bdc5fff3f4b4daf77e6227a09b7b64c3f22935dc1fe6cc47a83601a18a9137dd956f4844e27d2af84de9e16d0564323c7cc7ffd7ba11596ba22949df3e888e98442370ff3a10be5a7287af74ae7ae5245dc5314d8db9066048737c29463a97dee5a1e0991f0fc6c59c3a2b4eb7346a00c77f756091062e51a44f74ea6e23ba48c11d8adfc3f73367ba686ce298fbbde33c34ba7b27bcebd995a6dafc834df5e986b069cdb2936631ba9e86ae0b4b3e2a2afd198cf8226f130969125d44ded7ab242794299de62e5ef0c929ac1c7f1daaee1ef398f2b88f1f8c386124bd898b51d3cf158bca7ee9d6276e03fdb826bce5749a4b600a3da3ae8d202143fd9d0cb856f23bb5787796a29de78b0511caca0779f3d2dcffee6345b891898c013c006dd68aa9583676aa832d3e77ab649c81194601253021965867fe8822fa2f4e6ad1ec53d75464c863b7effb3def68a0930e306665636a2938a7a00e0a4af6190751d32bf2953da88d48e9010f58a693eab68bf7ba10cc691b00767bbfe58fcdd0bcf1743bcf7a0c0a292522cff96faaa8aa7950f346501128bddc8e1805645199b2db04edc2848d219b16217e85fc58824d07dd86ffcea51d42aa4b2a55a14fac2d48a819de31407c2ccfc3b6cc29edc480df1d79b1de7a5a91406ad0742d3a7329635cd1a997b26c235a9312734850b5a559fcacb721750b841032a11d20fe23596795c207c72d723945ea191ed46e5b4f08cdfd8c6904fed2d5a87cdd9f761a7d0f754940ea6368fc49cd2df84a08f60b1957a4d2d7b51bed64d0f45a761587b003bc518ed4cf959db51efaafbd7778c0641f6eba57e507193ceac99bade28c5eff689ba37633719199136e81f2f27855c3e7894de26b128a8a42442521dcff76780bc1a864c156dc6df4eb1c11374eea12bae85ac87c34c2964f98763b866a41049800cb47aec9e188f3860acb5e83fdeac4b901110b4036d08f43d5de3986ab4369b5ea25904e74d42b1eda3e032b92f49e0bc7be2bab2357757e34488a901da8ab171d4b178def8b054a28f35a0885dcd344b5089f44d8e84682c44c83a9b43f794bfa96cf71215ef929ca0dfb43433992da8a1291ba8ef13611620ee62e5a7a8a24c08ed2f031d06585047b03c7042b6acde2dac02d1cd9343b70f6e1d468ebb312717ee1f26c761c5fb866f205f3892a605b985c623e8023f213dd967acf771dd36842ebbe5e3b346bf957be3d40edfdeb417734ee802d0881e598330adcaf529351af63fd392b40b240682bedb8aa17bb71089375c20246f659694f01a1823ae6fb0d84cebcdb900e5bdf736b47fbd64ecddb24e998265f34661d73996b9346a1bb65ea0be87dc317577591047444068c683f77f2e766816690842e15abe148eaf18369f0d302b50609cecfc4d4cf095bbd21fc8f22db79bc7288e4dbd50e7290cbc40f701922e82f1109028f2f53d7038b22c54089f462edb35df13966803c57bc5df9b0b91fc7d1d313e37926196bd047ada83c5ef063aaa7a67469dbef6a3e7272c021fb85e76975e6d179e9eac2562cef3c234f7f8e343fb30462d9e6260d99d1b9c558b1c4c7a5b05dfe97fb3d7a9bd80687142164b108701e6044b477e974141b1a237ff06691301c572ad49ad01d5edfcd29ba9a81a1bb43598185f90f1643b004f56927ef7bd97f1329da3ac97cb1f035ec263c1d9ca5d278da15929938a0fa2373ce791351dd94fa3c957965ecd13747753274291e6f4e570ecf0d81d8b85d3332b94c8df7efe401daf4546347d0c154d2417e0a8a036ad0b14c0889e08ef9bcc145075d63b88e0d19fc249337e783f185fc460d9b7ae2b34abe5e144a6cb4af3502bbce84a2a13be1c4531501466301cf4d984e68eafdca4c23bdd618161ea2cdffb44fa891883a27ca13b47e83ad30c8788d230ece5988a53efa8bb3d0ace44bc2b8046babe87f8af61095363150cd13f0ca2d1a53b8c73d8c0b8c2c197253537d0fdd795366c6643187fafd19d2bc618b8235e7a824e2aabfa3c38d5a2e82a6e24f9f884cabb8b0c090e616b5273e703d755bd1248525434a01717cb0b860b4f767aaec7f3dafbc5111f33cd95e2f3a4bbacbe87d0c2241582480cba163894a58b02d7fd6db03e83a3ba0b61dcd5fdbdffa27ca9344db2d472586f56f812a844d893f521291ada971496af55f79b8f85aa478974c349008df353453bfe36d9c56d004fcae11e51e6112798c2b77591d0cd3c48d9b7861007978c511938cfaa3b284b3fffa8453b52048f310cf684f2b362a87322c2e156d4b42a5b266e68f174af71342a9895721d0a4e15e304e10e56eedf1d802457cdcfb0760d4a0b354f17d2041c9fd957a68b89dbb61aae4b0c926627909bdfd33011f49c9603ecfe0b56dacc264a6a833d36dffc0b350a463f627bd2b1e94e9281c98a886bf3b900dddd90205b0495b56db79dd678c20b7d74ba9b1bdb95c41bbe1905ff21f563bbff25bd284d7d0312b7a70a2e2ec9814b38e66b5f94f7f01b847392cdaf8d966908ad63e9c9c7b9c155738a885695c2bdb549144913f2153baf224bce75a92fc9b066b40cfa4f529114d237baf1d2f6c9efbfaecbc347fa4e2ebb81a03b40076e660ea46e2f7a8c97d9ba635677faab964828acedc6047838c250003a7aec09fd3a1fba179f7ebc71843a104ecbf1bdece1a09846eec732c87d8b1edb0c70d6f302a8ab42a561eff3a3642cfac16eb53a753492a7c7026c3a1c130c798cf4147b32561d2b870b09192fd4cee931aadeee2d2e7a36c61a92893389228b3471ef056807c6af7819044168004291c4e8b05f6d7256083a2d5ec08878b788e3d46b142d8310e37c93ad58ae89701961a0b12741988543a64a33d5dd5938fb55a978b51f92396451d9c7d067082c8fc9fbb8d9eeb0751fbe8697510dcbf9f4a0008abe18743b8d2f6c2722ce28a5307656dd128b86d02e9b0f13843e219eaa1ca83e3f7d29f5d3bb3b45811a2725953d9a1bd0603475090a3bd742ca56320c464270f62cedf4562c09675f180f1993304e852a0ada4fbec83d3faa0189b0f856547681ee7cd56d89ef016185fc0a60218945f94166b3b2215535f19b95ccb59e488c0154fe8522a506cf35258d7b96920eebbddfb146d2eb07d39771b8a27e8ad947a9c0c6c24d5b2b48393dc260e730dfc03a3aaf39dff83f1dd7be2cc5cf31e7f62386152e7f1e8ccf4944cfbd8c0ea59d05212ce0621b595ac867303b9ba1990c6724e676ff60c602fb34094e7ee944f08869bd5ce2cba8f68c69735fbc9baf18990936abbebdd3263664a094e2f4b9632a0571f85b215b0718f4f149bddaf126fda97abfe67cac72fc230a04462c1fcac7053c40f4c65b7131c80181caed082c8a6c0f5d5303ac6324b7a0b7828454755c4e581fa045e4d95ecb6ce2d502a907042c487a1067709f7f30cbf9ca9fd93cd43de79fde8d2b603edb3948baaabd00671c50bbe46b875ba1f0b89fc7e10ed1115d7392a92e8f00f0a38f7aa0ebecc7ccb883ac85801fbe04ce0b295db1928994bc404a9672651fbd2a757a552dcca7032125c204801d35e9d0546c58e618385523df38b02a97d490f3e8516802b226a511e2a926ceafa4e7ae8468bedc91a8418d8dbadd989690a6714b917e38edf378cf7e894d2dd40a1ea1d008e50851946a51eb2f67121546908467280f21a073f2d4f1748444ffa0d077a5daebec3e007d6e779a64401a9fb7c4812f262966d11812fcadf0672806b4a3bc540ab7e66fd184cce6d46f0999c44771b16b7113dbcd132f70cb1c2027c7620fc371e54afd32b0e1316edfbdb39df1772db1b74e3afc2171216edfdb5c1428bb959ec6efff9e9c9f14ae84ec23b7ff5303f7cf7e83ff2f0885150c266d09ded843adc827637e4646ecadee35f0ed57ba2df440dca4fa228cd231d934f3e2dd14d157fb011bf30871deace29ff9ce3ccdebd4159bdb6625c826b90a1877a8cf8f179e3a3860bc6da723a3b32b340e53a406eae792e17470133b133b03e51dfc3c33dfe05d5acfb0ab9d561048cb7c376e68236e9451e6476a07bf343bbe7ae0396f1c30f0f4d63465c1de6f620a19bee9e16c1078b1ce099e5dec2c68dbbb7a311e72b69c5a5090b3a0a90b6f552f5845be63d6de08708ee2274207aca6afac9066aa2bf61052e7f8f6be96cc260e12d3ef0b175957187146d437d8b87bc052bee2090ace6df306a0e9ad1b6313dce029c10dc40d8e778a932ede4441c41fa38ddd31e98c654590100618eafb55ff50ad1b0307821cec525575faaacd4640c89eb3f48df5d25ea23a042d8e25874a2c25da00974e82f9a20f26ef6dc577656593ec6230cf10831c4c73e41068104ad076cd261aceb91c6deb24a9e883a2ad30845b51cb5c7b30f3c2c90593fb0d115924a5053d8fc5a3d03b1bf19ecf326fb803e529dfb75fcfbed9ec48ab3536fd64dd9f849d39ef69aa0462739ec1c7c6d7ab4b58f9bb5d5e3396f0bfd6685dfe487012e3a9fe64f286be0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h45e1de8ee144e50f1806aaa1b0235654e605d45baa0f79097ce2274fc25947b8a369362bff06f836ba6a5f13d218e535dc19d3986d737ba66adb76344adc4b7814495c8b7d47bb967b419118508cdf654fd140ceec1390d762f73e1df7c976c16c09a26740bcf43fb9f9a34599f19ae68b03cff784220ba6c702ea9a3227ee3e137d31646f95d7b34ffb5acf6fbb2d69f508253bf2b2f896565920f48d45b48682d33bebed0fa20337990ff4bab8c509e9d2a6740534cb35bac47eb82311b5dfcfcbe2c5d284666e8eda548554ccf1331b55a744bdd141e346863d43077daefaef47f5b417b6d222be424a05ac8ecce6b861ee2c80a5e0baed3752cbd72d7b954d2cf68ec730c91fc5bc98c1758bcdadcc84ee92a6db18bde7c7f653469bd996e39fe9f975041b9addb0805ffd67e8b0c980b0a72e60a6b1ebfe201ac1081dadac77c374171d422afae4eb91e3fb848cc8a9c8e9a0e6a8b6c60faa04d1a274e3aa7a706e8b72deb027a5b5f68d9d1233154f5451d5a96d4b2b32a2ec7606a0ae57679eeaaf11fab33a7642a597822397a74e247ae14665e6c0c572466385f602d7b46850e26364a478b402018259c30513ec84adf0158f779d714d2ea1d4301039bd77cbdf5c5aa3d5abd632c78b18f6a6a429ccfc6885923f3e1d6c63ed7fe05a6c3eff1403f99f4364166d3f8ea317e5433d10daddc88066b4690adb59d41f253d2b694ea1e395788e0245154d79747e2eeef3f58e4c9325fbeb88c9a14a3ebcfcf8ae0790507d6f1cd51d1de8c3c8ab4d1eb4720d42bead98e44fdb0c2222653006b1719fa3ceb4e1d9a135b564b8fa3a6618b53fc25dff941abf7e59779fec406b7601ca5c2562aaa105c68e29fb8da305da8787cf08d1cd0e341b84917151bd1252a18b54e3e60c8a6545452173c044c265c853e327dd66d6ccf68425071f471ff717730a57a82681cc8a8794815e62b1ce2f2b2e7a8cd89e4947d251c4433d9459c1db031aacf2df4cd6ae5e63454db5b2458080af378cd137a865d281e233288c07750db93ac01ce02587c4106c55a157f28a1186ad1f1bd9064a0f690fd9913423863b661c6216021f325d33802018fc1dd46b2176a2d548016f6d786ad14ea4c3c557ab216b9f297c0a3516162b734a6b7d5b65138a60c411b69fcfe4ac8a3fcad5aa8ba56b468c72227aaab9a83a1a68a31b3ece4eabcda2477d1b4a533b781685cc59a700be43aacfa3232475bf312747896c48f6d37b1c85031d951500f826e5834219eb327a82122c2966443dc9b1cd2c4c9bd2062ee35d58e680d3b8a6caefcf3b965b4190e09b010a42a8a2c090d672d16e7af9ec8a1eff69d1482808797a1b8b9d76ba66212a259fdb5085b4a709c786cd17aa73c36f3af57a548f6e67b63eccc47c5ed69d2ec8466dd353620e5c3b7679e1a4246316fd7888c6b53794ef5def086b28604d5d6589a87e890d0787e1adaa60392e3850491e4553fe3d5340680776e0921c83c31f0df66b7a4cf3e9795c4997e51ff4d808120c74d1ca433fb00a90dd76b5834545d4fa915e83a28c101f0ad64cf6a1819b6b335c33f66e33a3f6325e1b3f23525ac5cf11eaae2168f66d46cb76c2bcee2e6e7397fe8951f60bed385cb5a06473b871fa27015639e9717303d55d73aa8f1d61098a2b3ce04524712b7382b87d080bef26ed041bfe4fdcf98863d714442d263b61ea7787675e6d1060c4edadbdc5a56275e1e8c758e5730ab996391b23fb5ae149e93c1143116086c05c0472c32e355338720c846080a7687ece6e399b440aed12ae4810a43bfa38de82c7551c9a5f94afc85b023a1b36c4fbe14d54f7881533e1eaeb45a9de58624294040529a6fb106a5c262c84a7785f9a02f03c7a86ae941c6b3723423e9042f5e2ca999f6803c290f9e8ff6e180ce89d6c8e578536750a2f3d8fa8659abc3b4911dac373af40039295cd9f54773a3a8dc53a25486978e87d2c13c19ef2cf2651d336ed8218e1ceb4c22305d6d08da748a8bd453bc9f7702d424fd1738ac4e6f93ae5190f8369a5ca9b2a5a3d1c96dba4cb76c9a7ffe742f624f4dc2deffceb55733535646c480d7e90791a37d3cfed4dcdf14ba89f7143945e347e6a8ad14a8bcda360ce7e6a45c65ce357f869f206c59c728de66ecba369bd2b2adb5a19eff281f83085c52291d14bb73322e17d02074ca7f1359c23d97d53fd1782852255bcd5b9a974b54fe4d6fde60092fb18626156a048ff50b9025d45fd69fdd0320cc56bac7b644cf357030d0bd35b898cdcb413e4aa26e4cd26dde2375f8c07122aa3ec2f71ba00cb8ef972d0be1a273540259354dca7cdb45d8afcb71ff6a5fb2731594383cab7b514862acd3846546341793cff9fce0e50697eea435dd7283536da02d3cd02d93da387e9051a4d957ccbbd116439160ff59f5de2bd5d34777ad503507bde9de389966fdced522a08e202b6fbcc30d7b9260d07345e43e3786686afd1eb46213e77de57941b779b4417cbd139aec79bd207d71bafcdafba6735071c8a61e05cb2f1af042063f510c2be24fe74eacf42a6d176adb4260651263e48261b7fbab9a72fc3c471cc77f35bb2f7f5dbe876eb8cb7be39df6070d032b5eb6aa12ed02174d3e10fff77e7a92b9f06ad4d8e110bb3231f23d0b4adb7920793a92207bf0b13a24d5714f0e31bbab2c762a89330b4a1004ceefa10c5c6be4ef0c1ba6ce23b6fa6306c98104547ec79bfc8b6da2652fd664fd1ee312f7a8caa81d4fa1562c6ec78d0caa3f89e984e7bd38b4514ce25777c1b47a719102de7906a0592835814d8421bda037e0c5c84bc42a2837b6fccc9a93633ab3613379e12d11faf531f2d82e695ca5458c7e0078df056d8a303af7fc4ad19b44f0d94585d61a8ee9410c59a3a2dc7913d264cf43b305c454c678b9ea1c91aa1b8e28deb58fae05d62edc7d3848407112fccfb90e41334af3d80940e9cb472b464ba28af01865ce560e0b7d2a2337d786e16b6f6048200de500ef57d9cdf3b08162f739bb3f0397ba7ef33b782f9d3e44bbc9b5079fbaa901cae937c38e67419c49de273cd61a4a807296677a592b6a19bdfc2d5e7461190c93e8d56117e75e3e2ff4826bf3f7a61726dfb58b3ff57e53222a54b00c1b91267045dc52a9af97cabdf0da323627ef4a1232388a5401fe44f0df7a55b5e995e987d236ec671f3e288fed909c15515a3ca65b30fc10a152fc29d9a4c0550838d1aff2bfe4d4cdf42e875336583832d27ecdd16e3fd50399450bab5b9e791faf25d56a83674a916ff522487ea8319a0bd9409a72960be2b367bf9cc930c7f544f76f0d6042fca051eae22b8c709081516a6797e40095ea54896a6f85b0508a90c1603146602f63d2c696d09484a97cbead9c08558411277c4c80589f391491ce9ca27beaefd159db03d4a6cda19edd491b4e469103f96e31cc9e0890abeea865a2fa0d32df5cb0e411c1c3550b1c4b1d90330eab9ce802e9ba9c650207eba8cae5411c78e0f469b94b57b758a3c4f29a03de5adcc38b6f742d0f3683a81f33a480043af4c3de8cfb4c1d713c0a32a40c35520bf7e2d3f2df5312ec35752e9670160287bfebe67525f7b4bd2ec7f22a2d19fc68b9be3dd1fe25b298b0220c2ab509920d7e1923b5af94cb2b9c6fcd60991aefbb064b70d69a1c93849e5dfe474b2a6a57ed078ff8ab2bca558a2de404852e976ed811514ab70af7a2f15ca3d0d6fa3ae41f1982b4f785fe1e843666b75711e741492147f8d5e3988883c68846d96bec524dc30c1250684917391eb68dbd7a1f288f69d09c9af40148e94f1867ffb67e4a1880318127d5bc6e917af01d9bc6516e6df5a75452d4ca66be4e4d5c5fcd0be9f116587dd80d2ea467d9fd1a4c29930095044a50172e1777ef0192b71d0ccdc994efd2641bb9e0a9ac13490ee5f7c4e25bd1181ff456a79bc76d1d8324b4f74aabdf7c9f27c69a994edde0d3550305fba89a71ab32b9102a87adf06d4715552caf0e4ed3825036060c8cd9c041f3929082cc2f67804adb48287a71fb2f50e1a089cc736ab016ace1e57f672ca6c822d254358b34ba6e4ea4ae3736f9c66738c9aa6dc32349ccf2970cbaf14e2bb9a620966819f3d94a161b661c3e6e2fe04a49c15476e1a0c177bcde68a8792d33c84f462b75cb6e7587462738d60b781ead82aae6bb3935f4d0f0a3321b9b55485069d724838f6e882528ae6c8d01745d5f04282dfee4bafe6fb32aed6528c30ae0e633790ab478be913f0c0bbd4a8208e98353cc575f5712d853716e1490f2c9fcbe61b163213ec21b919e52d18e131ba4f0362f68f4e9d3289fc40d291762d63514148e5b6b4de4953414b7fb70a574b208c6088e18c5c4eaba5d7920053917293038123f4283d1dd6a3d31b1bef0a9d4322785aa5b702519226d3dd0c954709d01eeb742e78d76bc6dc77105e98b9005afa2ac0d5b349a4ba803397bfb28dea4b22a3aabb06951634b1a3cfe7f0f7171f202364bf1f276ca3eadcac2b61ee5d254f8bca8cc289fbf3d15af73a81d2af4302ba83a1129a20b94e6249aabca5473af5489a0b088df32b87f6be4fce789bc277f1af1931dd031ddbb558621f54b99807e5ce57d99e6480ef59b3ee3c9575f934173d1ceff1659bc9119a7fc99a19356e41ce2865d1d54ab1a4e134e1563216a2638afecea8f51d1e915b0862bbbf77dcf42b9a0436243d5f6b9957052513398952772f00de87715686228023c7d4512b95affb57ab988a92882a804c202c759f519b294fb9c1633d57037dc913fa3be073f0933fa6454194366bbb74a3dba040527977b805274527041d9ca4a9d9f321fec590cc4742c47c87aa99891d63eaad9825b952a6be338a5881f9b81d2ca893051266d26e092080fb873dd16222eaf65b4e610a30661045dd46b7fafae490b325f7bf14e5db9fb8792799b70e8db2525d61df4eaba4d7b9e7f3169603492a85e203af05bbd35e454aade858228a250bee2fec0a946d74e14dfc9bd8e9a46cf8afa89983f1025124483841d0bd421fc443e0e452950d37a543bb133e41cb961bb432b8cfdef67d805073fe79f7aa834b5a046d5fc39b21cfb8cd4f81d62aaf56b4611c0e0fbe2d5b47c8ccb76b2926041e135a3acc7a963ae8f05ca3c347c6d6873d43a5f40be8914a6a5e993ba7ac881e5348d823594a3b14b8e317684fd69d71dcf3ee8c97cbd17de81d391ce6950ff89a18918624febbe3b43f4edeeef056a206d6bf476dff0d271b18ca7f6f421113bfba636c85549f26bb5d26b99f99ccc82ff18194bec3d50aad3eb2e1f054129355cced2753599cc86bbf404dd34242a2ce1e3782a0f8bf326beb10d6acfc22c5c50fa47c48029558ec305372be3cce62613817a16e85f7c2018fa72e1f1c43ba534afd7916adba7a3d21372f0b2ea317a40091990ab6f0101bb39b8239e6fffd25b0cdd4fde2077cf4c500203de0ff880862c8ae32bd44ac54a5692c0115eb0ed314189ec83fcf40e20f12a7e3eda538996c4337475cf29caf3ed25b7ccd99024caab9094ca3ca9c91acd48a84ef3dbc39016aec0e49696a29de4076ca9e0103a476384efedba5d2ec9a1701eefe31fb7c4e73b28c8100104f6c722245275c573fdd22842c99fba99ab511b96e61f0aa46d6711ee9a116ab55db902558eabfcc15dd4b30d762c2eddbd8c728f866425c75d4f632dbe0978dc115c596ca9555ebb3b316bab7146926ab067827457d063aa2a9b0b930aa31b90e0ef6b8e78a5408fceb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcbd993a77ca0d4ea1595c470ff80ca4d89ec5cca44a3854751186a81c42665fd1745bf41c35f25e7f00cf7d6d2afc62816c117306ce92fa3481435ea04c864314b07c4b410fe34bbacf57dd4cde5f88cb28fc7f43684202848d73bcd4e7377f48b9afa0340de6a0e75b89f0eb9c72eb385748865abbedbb72e01b019f817b82741a5e0c13949e2983218e68ba82110b49684b88c71c086d6fe381a50fc3da2ab7270d0fac882aedc20eae2cb153f2bf6d7086c76c2b4666f020a11fe63945b6c5fec923d83149156701d7b44edd2c0401ecc3456f84365aa9e63f25fa4c761f32a160ea62b5e142c2395f5eba21d85269ccb99169733e3cca0aca08c281e057a4f917e54b10d9b9e924294b67456cb12aa3b6138252c9a8f8763a4a2a2d4fb09f3e634e3a65fbda6e199091991175f29f7689604b1c0d3b3d15aaa24d1e4736e35fbfbafa724041c8a76b8e86685ed7cc61f48f63ac1afb13efc24913cdc31dcdd4ff14f932244b7bc23943ffac858e3c2bc81612408549de8e1c8231833b64adadff6c8591918a44235b3d3b860657e738c8720de98129b75c5300e75341434ee4c38d0f53c9c4c491ddccd8941dd9008399727fef672ff09375928e7a4db38068756a31bca84abc592bc4d8e53c3c5fce4d25e5cd6d552953b3f8a0bde0b54070c3f5b0c574f291f60a303d6da6225e911dda28f2cbdaee32685ae4da9302838710884dca82111af4c78a16bb9e4c89b35b063ab476a96df01a74a4a7417d91abdc0d843746b15efceca604b6b34ae1ee12b4a694960c54cc320fc60edcb26e952c85595466b3709d616f4a16761b69b5eb8a4477bf558990e6fda42ed48802340136674f57aac7af45036a035556959c1d3c31d16a099db25a1c88e705e258c4510369e432b2155b570f5b54e451b35e53ba1f441b8f1652acbdd2106ab2a6461dcd7c3bdff85bd441094d4c16a42ddaf860467f89251068aa6d3669f2076e2ec0ec390b5189f9147371695746e9c45211489e2643867310456487959882bf49ac6152658ebae84c403dc0ab04fa703ddbb3e60a2e69d7ee68b80ca04c2ab04926e9addafd1742fdd6f148a52b734a749172720d52a40493dd7f5446856e2a0d8ad6939c6a01cad4ac898f1b1fb12ba462df28ebd5ed44e97eb67c344c5ada1d945d310348d0ed0e4e14b38a90227dfd5013482304e522dde16c05b88c63329cc9a623b9d91cdaa3daca579752e32344cbc9adc9aa3ab58db56a5b41140c2a5d30b0e59bd298e9905db8594765c1a6c867e7048b086da60e0d7e2a75121c1b0a8f807ef6af5d483c0386dff2f5cf735bffbb268fb58e8db3f38802094f384877dac89cb4b26c8f19ccb42b52640d35c01134f9038a637ac601c2b31690b31408bfc406e216471477b478788e69e87715f3d83b262934edde5755a66919a29243942fc1e64ee38833b9aa5b6413fa98b29e71146f832e7358a062ab759867c642dd05650e42b652dc48c9c2a03cb4a42d393e7a1cf0b7c707c53d45b3ca95a02db9645179ac2c7a75ea8e927fad71e4d8ec048af993c1499fcbf76f595fb409c8fbcb37d92c2d6e91cbab05b8feb30d5b1e97aac0de2f2b04f31f6f5b2fe9383c786a96cb045fe54abc41251c43c68537cf20ab08af356e37f77491a490adf11516f22c984a33034def4a21b1273d11266eb24771a66e8caa75f6d4ea370376217b215a5672942ab8fcd859391c646c30f348001a9f058135b3b14def94dc2561c77bd3f1a007361d46efd751f67f15ab89a8e693f86949cbf7004ec22fe945ac010c6c6e4b2a9e1399d72d674d5e896a32b99ff3c1c853bd08113fb4d959d781a656d1404f0fc8b0ef2af915260981751986e62f5c0d54d4d9eabf23d74097336d1ead44a116f0f54f17174b2dbc2afc4e7fc6ef718c4bccbda436171fe45d4aaa43f2306702613dc579990037a49ac4cec08b8ac36167da3e62b4cf851fcef55fb7b25bece48672d878a3effbd35c249f22370358b6c427ee7f87d3f75a80d61a2ce34b77a81ac6352cd198f33a519ac4c18bce361cb93d4d6a506cb97bb2fc37e44e79dcc175ce86e7e3ba51b684ec3767e398d703647cd8cabf95a8b4d71555b0449de8d86607c3e2922b994091ca7794cd158cf167635fd957207c99f0a3c0c10f2ad4bb4f141333d7ee969e07999be08341d69068c86f56e3447a5bc1d99bf98d7b4135db4f3303ac10e6c14f2fcae81dd4edfbeb823645d2529473ffa6447748ac1be5c5ae0d9d9cdf2353e167d6c97b7d370130a68e55157cddd4663cb7f7b55e3231d46f37fef79bc8f18faeec2bda8549eddb561ce058c6bd9c4c77e54265aac1730ce29448570f3a003fc807b5148c1adfe87bc61ee5ad1787ea094f1a378c64126d25498ee0125bd134aebf895b7d5b4a25f5914ff75b03c5315ebaa2768de43e46aafba69c05e7ce739a5255bd7684a12503f01221534e0e058baa78ff8ed17f3d4929f4f5348844a8193f64fa7929ec8696385b9538e906f3deaa56c109357ac41fc316c4d2637ccfb246266a6035ea039848c323cb50492eb64277759fa5f59cf8097da6ded81e5b9c5d99342a736d74f30dfa5c41374ff13651080d63af6f88521d0270367d031ba582cfb0196f2b882c3a7ea6e10453e7deedc94b32413e7b7e7586ffc7c0b62404e66a274e5890b616b55515e720658e81b6bbc4f5f213e0e0b5ed2a350334733ffe1cf476777ddedda14982d5f7f897a80dac8b7f4849f271f7dfc45afd0ffe91b89f346f04ea6cad7788257f47cbbcf85d1055f03cca8180698db37ac4fd576d7011bad39151501cd4c97adc58f59f79b21d2e7436be7851c9df015d3dadc6cd2283165e1a715b1d6b4f85e8e1610233e58236bf08c2510699df60131cb44ff1f0a3e7d18c6122418f2c5503f5d8f217b4083cb72873d72d911b9307cd5bec9703c245cd1042ebb05c1de058fb72fdddb1f35ec6e6f5c1f6b6b8d5a1f028d3fc88e442b1570a650ca8649e8d63d4daa6135eb045a89a62f754422234f084df5c810309b52c0c0e3ba52feedaacf571b1f95668640f3e8ff290506ba1ac8d3ca7a75d4c699b767f12706b297839fbfa811e1603076f371fbdab9e4c39a110802f25c529a280ebf25e2fa3839636951fa2df5388e4c1da85be3ad796ba30c6cbb5f6843a300d4322b06d383faa38606cc205af3fc4b06c7b4b580d1e882ae1ec5bcbbd419a471181fdc16b047e45d0d42cdb6c6491f266054bd42ae1457fbb56f5e1a64bae94b4d081d97e7a298b8e634c342de1f177b90c60cf20fea9f2e4295e24d4b9fde9af52ab3308b1f213f425e66a6e0c45a3e749bb5e419026b202f32c8bfb69378a06f062f3d706fb2d474dae125ba38f0d2ac215df651424873dea8d638bf2e35f2de018c36c9704b19d2936840f3efcd88cbae2758ae204daf3339f118b4e6239ecd20f951d484a1194f2e613ac59a67e1afb91c8fc9ace919832766e5a255cb3862400b234f074de37fa3fb66d80e8ccbe4e972bdb200e92e61e8f39b2a4e193b144d546206267e71d4658ad42a718aee77c55900ce07ac11bac6306a809b5e303dfdab39264aad0e75a7540bc20e3819bc139a5cf827a5e991e291d072bb7803dc4ab0c74fe1e5485d748ec3f95ac2dfdcead4de77c68d365b47d6adb2f5d6a184a447fb90418ea7520297a0944d76b2e6e8c1cacbf54c53dc9da3980cacaa9cafde3eca9cff09ef890a3816d0400579fdea43e9e65cdd7a75eda8699ad35e227ea8179cea4389e73cfdff219d23a8d8092e5715fc0520495a6cc7b165a062c9f2de3716e7be532c74d2b4bbe50e6d7276bcc50fb94e48b3242d9493546c0a257aa008369b1385c521ddee9dea6a11f533912465f9c9d9a593323e2c794b049197684f84520a02731f375e72cfc2c67513ef38be9e94577497d9384f6911e3d1aabf679e3b3712d6a32693ab9b5f4c005da2732523fff7d375956518ae8c2671bedd65278c8f3c9309d6cf360dc450964d72800454e0ade19cebbb872faa5320104bf9211913684ece165134a071130c6c87e5a97aa0d923bed012daa8179136e08a12623cd3a6b076dd3277bf2e86c4e41c64db69cf93a33bdbf6b4a50382e6d02b60db329b37ed946018d4aed79f7947fd6435989b83298eadfaff9aa23f2c5bae2fb40201fe905ca602ff5c3608f55d1b978bc448e77871f468cb8c3940ba5104fff83938dc1781472e514dd4d24d019af996ae9aed17294afd801df0fcb3e1d57dbe6e3632b8fd8c5e7be0159878b5247b81d787ab2f1ceac287f6f012ebee11a789db6adb55b67e66e0c9a5c62cd9de64ce6546934ce64b4865eeb9f9ea2f382d180248d0ee840ce4c05062e338af9a59646e49f779b561e789ffd87fec238552147dabc0598bca4f302de97b437f2ed097a9ff81f28b06bd83031a6c2e4772f4ea7491c38fc1ff31b677721d9a56005289dbe890bd828cece62da7cd245b257c372ce94260a5de2d45ec07cb5f20970377d4853aa834e7b804004a51c15f40cca9fd18cbf1a9883624f0abe5a7b37b3273f2fabe2f00f5b543743164e60e4578dd86f1039a42648654ee1e527b5c8549ab91aa49527e36d6eac15ccc687a8d9bf760381aff0c4a0cd88624d2e50e1e075c2fb93751e68918c7980f84b351293b78a026fe9a94102492f9c667deed499b63352e9fc5fec8df77c9f06bccf7e94a75a7f9d436e63e8c1ca10f2c6346e3a08e6615c78d6855ad10cfe3f9e6db401ed82c5f7061a3ef0cb75fb64dd8dacd62f6e3c45c064a6fa551d85aed62419f09d41d1a4ca8f57685e5eb3a9f7372032cec727c2b5bc7cab69432d3931796ab8396ee5f89758db80792fc2a4cf9e2045c77057945b9293efe5e13dc54be2fb1b0b0960961296657824f7082042cc544abc3c1432a606b397cd994d60a1e16c75ab6fed5e517295a456d21fb736d02239020cb32aa8cb33af212cd89742f1a10eec90a6d98437578776e4e65fbdb906182150861083efa5dac9cae6ade73e2cd2dd9475f77f747f855820b4d3b8c05793f3ac63260611ffff189e27d71b3a195304268b6b09d5d2fd08689e327bcee7c7fec310d4cfa8b494cdafb16732be4178341d58798abc7ef572590d63a4d5696a7589ce984d6d8122b0259804e44eef0627c9c7ce92915db96c2a458e1c826da61080d9a42e472260e46d8f3972ff06fc8cce3a79cad4110c32e6aff56e7ccbd0a97f03dcbd117119278743c927052d6ee5d3c012106131c5631fb0bf6d8d671bffc3012d86d0d6bfd1d995b39cfe9992388e8aa1749c394d09412671b442f185e5a99316b0e078ec2ba7ea0f2c2ab02f16317c19084ef44a8b31f58b13f9e91aea0606387de87803e5c3816f1213a24a80f3701a994ad7121d3897109317cef87cfaa16dfac632f9c5ce3cde269a22148fe19319aad305509a97bf5ad8d463fb49b70d08f48fd4b4c45d1498a8b38e6bbb33bc1992569f7d520ddc0ab75464efe37ead072e07f90639e879c3660fb3889b77592bcdedb5287538ccb1a8bfa6ebc656db0b6b0df3f8619e6b47be57a0674d167a173604dc7192fbca322c131742a357fe4d13f19a789435f3b36455df37550752b35b8650fcbe285e1a00430add7f6eeeb38ec84724ea852a907cf12d0b9c15c524d7cedb3eddfc728f9726efae3b2cb26fdb02c005791bedeb98fcefc248ece8d73f4d2648ca4a6dba527570230c43931b71cdbd1d132634b0d046634dee612234c153e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd57c060b11e594402b5ed2556f35a7c2a43629afa59b1720113dee2dfe913f142d4733971f7765c4f05888899a0236f208e1869c05f46ae41f6769f710596edce4d84e9eb596b8ddba08a096b418bf786848d88a0a9f182518e9e83204ccb65d3054325ef1aa222ebc6ee6f01c9f749a1247303c725502a0eb7842340624cc35d6aa2b8eb0791270f705abe6778729801e416e84c813c0e02546aea385c106a1ec2bbbaaa27e1a4c8a402348feaeb919a5c5fa158e5398892be5dd64543b81d9e708ac66da754a2a34b30755c84ee60370728c66fffaefc5c1fe245ac8dd0b50c08c107299123ed02db80d63dffbfebacdbee158885f8dccfa04534bd6d81ac22dbf3567c45b3d38b7fbf81585245657776553282521d7a7744cd7d06561bd25c851b7366d992eef63894f76497cf9c0cb44959c2b7d7c3d988440d7a86546a092c37b040ed95f7797b4335eec7604e6c27fc358dbc6e71944d8fb8a3594c8e730792a6f20927dcaa048d30763df9729ba58470878f07bf8641bdaeac505d805241a3c01353147fadfd13d6a32148ad053e2adb750bae43feabd336bb81447555f2c92ebd8f52f8dc1ae85421f626980151123f37f1abceeb554658dccf95ca8037774690845ae57b949526e4bfd6a898bb400758febc5a849455058d1effefaca457fcf842ac9668bda54b1174250ce9a56a2016eb0e85e684a43896cc721ce5098cd79106bf3d8f82bf5157a8728bbec66d135cb73c186ebcfc587e0330426f882dacba6fde3b76c7901f2576de9dd200403e6c5e13d7ff57a016db7b9dda2680f8e82868f189bb89dbfcb9b3c627377e4c30126ad40baf9462fd500b770f158c6205fd6a9ac42d5fc603e42e0348430f044e77c383f59edbd36eaa727d811b9981bf0088832eff2f4fbc745df0bb5ece0e9ff6f8757b14bfafe1cc3d71da374f18b47045f87282c0fc3b6503edfddb7c22ac54f3cf08a3b08397ef8d303b231bd816b1928f87702839c6ac4da991df16da460f80d5f596318a6978b76be1af69739a1ae5e7dd9820a89974f9df51577f915ed4a86af10979f66faf8ddb5297fa2f88c0066d0123e303652affe4440556898c4dfe4538b9076e6f606f572c3e389f1693d1412c6379f245528eb7812fd04cb926f433c5760de0c44636d5cc1db8e82a87bf1b10026bd5c2e73d4e23cf38dd99c86019856aee68a71cf4ccf52d24cbee08083c810fbcaf45c814c154aee56185c02c8910565ff39a84452ec9b8ae52af3d955a58eb55ce7841c6ced3270950aa792b6d6193308a91e188ef5833497d72eebd9534613b4153fafdee475ef1a4d095be70a7393f25ffc3f345eca25c0b696e1ab6e225f0f4e4aacc15509e64f31ee2d5f0d840dcfc1bcb8f03170568324a99fc85998dfc82a5313f848af8f7f9c302f8a5b66d256aea009791a8986b0c224c95251c0410fa99c93ccd5fd2ebf82d71ffab6f4e3755f31c44b7d0c00e846b7562340d93f12431c838527834db239de96300c5da5057fa62ac6e6303fd065e13dc42855b736bd8c66956fd7bcfb86f2988a14b305c7036a3e1acc173bf8ced067027be81f2f2cac930271fdd9ec66acae283098c7001546c824b2b2ed6e77aea052bef07e6c592a4b79d38b615db7a1e7255e004bf7b0a62ff0e5ab8123190f0ced2deaea57d7b9e9968b1a65cf737cd47a90e098dbe21d55a93c2c19be637e3d7a21f7dcb02c1337eeb02a7b129da6fe4119f07d48cae42a7406ea7b57e5b8e0b07e221d409a4f294b67ce4f8ff15a11c91ac1347983ee601ab8a114c476ccbb62f9f99e96bbb8a71f604acf2f9c83b2846183e05486b5ff4e819875e5913f02a316e7489870df87562b03ded195e8a7ff70acafa7ee01315fe833fa837fef99095b1864f034e64742c27360b7020b1d5c2b017ace36d5f5a3b54db311f43688d5a875a01f5653fd4cd33e6fee0ca9bf2de4ad767acfef7f9476932b5e5492ccd81544872b82e31289f486b3878f61572743ab7a209fc2c2b0ad352e1d76810f3ca6b35bc0e0e7b55ae653c768a90433234e4bb61ddb21afb86bd8cedd8f23c0f77f83908b3c693ebf27f6029bb24cbf68fc90688f8ee73243e3f3c48d71fd6dd5cd67e8bac91160f9c1f96000880349690f54cbb021ad5e5a55e8aa684391ee0d3ed5062ec9dc4772c9901cdd2e7063966cce75d8079af1e3170fac354b4272357216b86b50d09e4ae5ded7a8bfad16f3e445dca703cd1094a87654512aad5f36f8f8850b500e1bfd30c8717fe254c6e29a10ece0aa19c7f5b3a7441d62ab8675d3c257d92b3b8d5df692fd8bbbb0f20fdc1a8192b8b943f9cb58ed461acef7555010144f2776787939438ebbbb66c907813fbb0014e7ac10f3582204174146a2cfbc2764864dad6187981decc90c5df8db32452d8d9e9203a6b78eb72f7c3b132794cad392fc223344b3318bf6324d6772443e25f1cc29ebcacbbf5c83bad04639d36913de171682edf240050f865fde6b4707b5d9669f24ce778339da34ebd989ca1d0032ab2d6233d0681aed64d59735ebacc57c66ebd137649c0764f21c4baa67833860198b81a3d70fec2d1cfbaaea830f419386331284cf49936973170a7b7f552c762574d0b3aa952910abb28738fc4dd436689b62249a336cb3aa3a8c3d88e80771325fe8ff3c8c5a5578d6c69808463cd68e6794484d922838d2ed35290cd5be87f8b2f17176f3a36780b7fa3f7e9ee48e8ce1b5c3e2947452f91b0bf716bdef7c2740aa983d0171a0008e987621363ac6d83484b38d40e7a0ef58f0f4b0e683b35a503a952cd6c45cf3e15edb3d9d6d2e5510d22a51b675c58c50f2281d021dfbf1f86717890fbe7a962eb45dc44597ac2c2020ad1aedcb837b7f1ea72ed73e87dd0d444e976acac581053e01da30dd0dce06cedf8d552af37e29d14d18a9cbe47ea5c000d1d8506f155d9047212e28f4d83d29248b128f9ea908f6e43609e619a48be4fd1736107bba6d404f2626d10666906563a9771885fb2b809dbfdc52d2bc212fa07a4be55a0984d4bf63d1396c33b3f04c069687d66295d5f12511df2389f61604e36cf451358ad4a7543edd910bd53471f56885f83c780b812e440d85258f357993fef7190dccdddbcb5646d9632476b37433bd52155780a44203700d7dcd5ce56457990d0df5cb79278bf5f41aa5f2aae93120371cab80f4b66db0a682be6675627b15f693d33d968944aa0ac3d65a2286682956eb16a3ac379b6d66b26145e49cd23f2eef4e775b8471e6d5405b441f63d901adef77ad9adae85fae7f1c0c06a0b818a999647a8d5c876c7a2cdc4ac0e342711f44d56f6338bccc37929fe437ab407b6ef1fe404a29acd9fb62b20a2483f1c8093c71d247a5ce65ddb023634ad1012e81c6e90187a6a3c0c32ba04900e5dad818d81b20e44915fca878d01bd0711012e1254abc6987a3e963bc82a26b63d56f112f096902fbcef670307069dd1ca802429081cd7177a4aaa9dce61a11eeeb3b0c39fca259c5224f0ba74803f604ee46591810dbd1924cef306d3607a309143b9d303428af3396c28154d37dbc99955415396efa0972e3e9feee970544f092803db80cca32af443e81ecff2554611b71395894f6046b3db71172fa66c02c53e21f3c56a0afe470ef47aa1d4625245894b74c53ad3b04fe1757502b109d8388eb5e973eb18be5b16882c19f2e67df40f8f2ff589eb372124a5b0132aca2bd8748f091d45cec846ec76a9a8ba23ca3d84b9c029f589c36a85cb13bc7ee4744b0701ef90d1e9a164b8935f42fb9a4aa7a23cc3099a720e195a401e819c3e73ac8c902267a1ddc2bdf812e6453783947685df6caaf74949253c886781fc243592c3194bc9e8f61e7ec3350077719fe0ba89a2e655bc2af465e5b37a6be769ea64b4d4c4dff2ed28dca7add7777a6e9ec5de3208d82326b329d7b29c0a75c6f8f55418916e7480bf5c8264c80a7636639e6826daa27408126e9d3f15d96b8dbf500adfd8589654b9400e54b76f24917618607d7e0ad6a4b416669493b74970d22b3f07e139da21010ba602e727dfb726512082fad41014745e1c406a2d5b3d80156358ad4e27ef9f92a1c8e75475fc7f0437654008e6ba98d531ed85fec7a85a2638114205c24ddddf381efd3d5d3598f8fd0fe3567ad40f859152eef2eb1fa4b44b3d5d1925bff55234c8e1e06045bd708dc094af57bc81e267c8b206a3bd06b7a9ef4a2867681f5b48c709043efad8248623532d6ea892b9a7b0be4767dcbd13d7878f2418d282f0c07d552355fa8e6092c13fff4f6d327092032d4f9499fe2497bd77b61a83fa75c2bcf7b97573ef0438e487debd6444b766e1a4ed120a109e19c40b151132c48e848ad697b23491022acc21388450325f4ec45a492ff258a5243ce977065abbb66f75073c78011936a8ed99dbc03d2f203d35cdf2df010122cf66b4c55336cc78f45efbd45684685e7641bb3d846ed911c5d37900394a611560b44fdb2134353c5ed2a7c3347ba81a9d59e0b4080823cb76163cce545db5278f72384ab56314c66032dcdd281a24b523c65c02ffc8ece3e8ba654c6cc6b531568d75d2788dfb1dd1367e6abb643692c152df31662476697493606fc7a3e091bf151953a525cfa7375b8a6898d4c39e8ca3e1fe77ce09956acec9de04bb8faecac38f2853bb3e4d259de1cfb51dc5b662009fe782b4c9fbc7bef286d8b1d3314fbd95075b4084241d5595127676eb6eeb9472789240d8cb452be4eb97c8d5a6d26ebba2c1b463d5dde7419ad3d6c78c7c1907e5bfd4d3f6868ece7c4c7dc5a8ebc7e01f7b78d1ab29d209d6492473e8a00f4ba23283a31a63bc74f909b1d44ebf8d4ac3fa327d2fb9dcb3db0c483ceca05e3c5bfe72c31f7d30d98a609d19da1835b7ba47151ad0bd94456bf86537cb74c6ceafbc75e98b2ff383ff4a5032c229e81dea705a4feed69533fa551dc2878f01af3cc1244e66a0e6607479f16d3d4aa35233e8ae61ce0ccf3c9cd9062cadd3d86c0a5f6c9b8d6d761501a3763625906e88df7c913b7e9d8bc8e733c590f24185f9438b72bcb6a4b6b4f65f61393ab4fae62ff1ccf5a8cece0414f9ada7fed69e6ed2350b8980e7f2c5f839691839af2e693d6f099f499450f099ebd6fadc983481b81eb5914cc2fcb2f3373ac03d6a969191c67944ae5136f8cf48274bcd68ebaca278d0e3184c73c95391b003909a1c355addf1f77dc9dd02110b95f8a6fecddd3a7bba62f6704f2ed86bcdf961e5783fbfd1393c5ca103846166dc21da60ee070b1bf5abd24f4bd1d68cdf716df02c700f488f6dae15127b771f0588ff2a9d955f5d2f66c133ab9144db9a7df6f1601ba6b0b8f490865ae51a49ea84da8bb6f6fe4d3f8b36f48ea4bd84003fb1f639ea9847f9a93143a4f8610ae675e675956c1bcf9f35e286b499fd573b8cf6ca2cd857143b6f5255e054c7e7a5d9b29cf06fc953b5b002deba1d6d5fc9b7ca7f843da903ea1fdb772c667f7a55b8dbe629e11d567a13d5e4e75f073c6c4bbc14d750797d430de19c8b6857bae6b34857e60e9e4e25a203d3aad606ea2e3b6f75fede71bb02f89fec625b87f3a628ab775e154716f13f07f025754c8e90706c12c847524eecd899fe938d1fd54dd2f164203d17be65e6a774259b0f3483db8b0cd1fdd6a3ce462db691a4ff36512d23d9b17cb0c199d0ebe0404f4d6a2dd297ab499bbba76bb01166959fd0acbed6d409bb4bb15d628e689119f8a0edeeede;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbb6658ffad4513980a96ca9fe170de9669b357164f5c7ca9620e64f5435cf5a881d02cb726a4e418f87e4c555313e635961f86523dafe037b3f6f5add40fc6ec9eab22908d85aa65aa1d7be88a491bb34eecf011ae5597c8f5bc276da03efbdbcc9988029d1bfa8f54fd2453321df255713a43eb6ffcf92b69242a1511f6c36f7487f57929888f87809c4f46708eb852dd6b32d88811242daaa42237cc7e7108ea5f9f3912ab0c3382f42abfc9cf2bd55876f7c76e2f0a64ca45b1757b0e5873fc059390f7e81fea322903e5bed55bf556b371d4f6335ca517726cb04dd8e8b39a164ac38b009d79dcf13356077b57ca6417c2e63050b2b0e73c067b5a7f19d156fdc91e3f6affe01db22266ed1e8cb10a1c45c5c60ae2c2878f520fca8f021df937276b0078b5c90e52dcf930e58aa6d04aa19ab9dd2c8ea752713131eef749d43dff7a54919685f40627abf55472183a1496c27fcc7a13780dabab3f65322922f344b8ec40740f9bf1d1ed7d535e10470726831666b2bdc34d915bf1eb83ed251004eee7eb03b4499b28f88611e867098bc1558b0f37f8276446879978eda7904ff72bc9205eb3b78a890a29d1f6442a445ccc317ba0dbd52e4221cb95e97e893ac9ac2f906d8e0eb985b92e37a7698a581d344c7713eaa8698ed0023473ce5f7c2c808c91484c3f110a6eb1ff90d920a48aae874b92e384e6dd65a52bb3070c4aff15a646c6b451300ac956b70e892074e615d9d45a8e75b5558db2c16246f40b556b7f7c072737438de24af5bbc493c46120c720cf05481bec0cf6aa180d20b1ca73ed4a6bbba5fc1dc4c998a984394d25d83765ac6d418ec3f1706cfc32e33cea0943d7d3088de6975d41fb6e30c7de090d7f0030644f563a62a75af2daf388dd8fcd2d7cc4e5c7aff77c6db13f5fa2d0b8df57477b61b8007b56803ae679d8aeb5abdfd44fd26f6c9e9fe44292ec64421c486381ee4867c1d46133b0f5363384c2b2b747919332111de778dcbf7915cf0d55054b66ed3578fb5856877b68012cb8b92870b4e933cd9e080ce37accb4e97306c1543395e148ee6728bee4ec8443572c8955d4a807d3a47bf717d0c780f8b37790d5788b60ab96b85c0828d75168d4129221eba303177d4d12ac34e39d679755a930ab297dc4df1d1a6563cd00e324868aa0cc5b6635f568f443694566d62a594a53f5610d9b562e5e2300e1008296daeddcca87fa8ee7ef3d8671e8aa2a9a5446abe7876d6d2dd1aae3b138c1b54e9786c0882edf19dca988cf2fcd3c5be5d586bf30e37c5a867f15e712fff4111773048f32ad0fee99f8b4164688c56d5a068e6267c4be562de4bc12b7c8323a3486574b22760b8c26550b1b9081e57764f83604fbb1be9685054637243c47c1f3099f5c1a436b32517d658fac328de9ba36130423c3ace63df97bb880b880dfebb9c0bd13b2f69beebf87df3d2fe090f5788e76584ebaf55e612991b511c589ff80918dad3849d28c37c5c6d63fc79abcaa2b40147bbed2cd7528a7c8e2a8750ebac62a9b9c65f06c65cdb004a07ee5c5c586202f2b1e3527fd882b36d83adefbe1a57352153bdb888e16513dc3c3480bf81658a58adf7aadaafe002786b34721a67f12434c660d6cda5b314f308b87a852a8377972a0c3d654843e7aaa714a4c80b48216efe96025bccc0d501cec85696f8d5e9c2948964ffac25791cb1fa6b09aa413bc849d83ad04b57d8011993a15dbf56d602b1f099b9389eae414e6c8d49aeadc4520205ac5db8f02d120ed22da92218564f27b40f69a6f27dc41d7d07684c122c7e884c56438788e8e6d4cc4769b46643cca31336e41056569bb27cd1f0ea1cdb2b87f08d771507e2bb584d41d8c0372cec6ddc1b1d2d63ea93fd0b9497bf499f05709400e6c709a95c031ace46a83982450271d5b9360a778c8d077ed99eb0d032e2bd2160c2679d18374ae427dfa0e646437bca25cdacc7a9670bf8967f3423cec179965ccb9a6aa708c16edcb87b56cf787d6eafa796d6f379a4f26cef5fe2b978210e028f11a6c9410995478f85fcaf9f51b961178cabc2a067758326f77c2a87824572b9c4a779df29e58ee32dc730219f24aaea072a52fa39518385005b7814343af5d4854d7e5fbd48103f57b5dcefe2601bc3bbc73a0775f4a97c78972e6432fd7e89139d14950e9b451f7368d5f6692347e21ee61a7db9485a1cc17fdd0242ce60c35d994e1055fbc9463eca360a28333272efda90202bac09c0572addb21e7bde7f5cb61460b450a2f0a903d18573ca68dd81d0649e8d8f18d1843fce0436bf5099fb1eecf7a71dbf2a9e9703f4b433527559f7d782b528efbfa103eaae06e672b614bd3c29648312099e01afe6034d547811662c50fcd9f210fb0b37bdacf89e458acb98b3d02f1d61369519a55174443897ff0363506a839ee39fb2f6b89ec28aecf1e517b41def8b0dfecc3f3fc3f18ba305d2d322a3912fefc5d3547284c5dffe3431c0a713877c71c5f941d2c3b46cba27c868ffd840d1e8a94189a7408a3459170bc8fc7fb962a9de7a1978bc8615b43e5d41e07756d52051f1c296742355d09bb0919cf8833ebbd0f1dadd10dd62b7265151bda49f9a169f47192e0148097260f723c0e504bcdb1254893ec86e33d981f283278ec6f8b6f31488d8000c8b05cb36b515ee0ff540e4326269076512cdcd2c4910efa217a3d15e3e73b46dba74e7b36ac6370f5b3dc15220c8d671cbfe440d651e09a3dc7fffa71f1e1a2efbc5fe46073caa6690e2a8b06d0324d3b4d2658a1e895e0dbe4aae46a3681212ec66475847a15e139a014938c77a32aa1eec4d14028278473f239101e6b4c301ba29599b93fb19bc76c8e4e7b6d54d837a9b5a610fa0fa1e19402bcbd6e5eaa1ab5c5d8cc36731065f489c82cc059b1ef9b34c0b6c66801fbdbff0c9a67dc0332c19d80a42b5547b711c50e83218c3710ba86913eef2a9656a62318d6f4e59c19fac1d414484d5e833f656027805700024aed26ca17c6fc0865e9e4cd82e954447ba8bfd913a5d13704612111b886d8dd3febd9f696f0f3a943acd44a9bd5c78c72e148e006db3ac93347c3b67d48c16c9aec9d0fe4d8419e12ebe532bcdf2a2c4db39487638a43e02c0666405be51bf7cfad9ecb8f1f3ef36ac9f22bfd45aef6722814832f675c0050e5af3e124602bc8b30635a9be29023443e4bc8fb8575a6c74a37de8f64a8a3a3d43bc6f5ce65061866fc7cb9ea4aa18fb597255c8967ad027fec6328ba159e418c43a84785b4d76d0d53a35dd0742c9cc4aea07011c164437d4f461bfb7581c16e8d1f6632188d1bc18e2179b92908824c9030791840bb45750216db7435811af914a0d1a8a75ce8b564a87d38b1570c460583bbc761920fb9d355c65691e8a0010a59c455b725cec2e5cca0c0991d2c25ae02cd8c91ffa5439d2573c248517310e3fcd64eaa2457c2d8b5c828bc146e6cd1194606a84578a5703487a0b51d083a1b6bb928a55213d9d31ac726e55509190609df18d039a54cb2830033692ee1d5b2fd165f0f1c0785429e1adba0aefe8222b92a15bf022cba8346b8dc75d1f1303389b62d7af1bba02ceeae7d0b814d8df3712150deac68b8b73dcad10c38cc7d4c90051d3ec1ef554b2febc9c8748544a464024989ec0d72747166a1e6ccd0add816f0243ee2b7ea377a7fa85c798969457a0ff99236fa8fd6303b3840bacdf71c53a7207ab58cf9f0a08dc30abe75153795506d4fc207bd22616308dda14ded4ed5f03464fa31b45366f06f3b3e7df14f6e214fdbeded90b11b0fcd7b8bfbd6c2d360fd5fff5af8ab1936a9da251765c2b802389de53d20b998ec5c7a2b690919d65bcff321a6a50b400534f3b65b1a37fff705fed988775021209c7b3ef5ff13aadb7ee6dce1e3a187cc4f7859ad304f69bfce7849a9c2b91638c10011982f8695ea2e0a5969a36bfd90f5d337343c22f1f556cd2ebe66ac384eb49b8faf0d565d227032cb3d93b07dd74d1b8bcf959b028f31694074fd96fdc4723f6200c46df66b0dac952c66adf9427c147d581cb074910ca7c610a528fae9ba60fe7c1e04234c0023346acf0644685a0767d2b2ab5ff95e0007b078efa0fd475c8ef043617808b2bf8d2a1c1d8321574de155416035f0970325e0106f8504811d6e74546950911a1b8d81c0fc9b8afd9e5ed28e55df4c8cc1c195ab612f16790c83b4944768c4c3ea2db3b879067fa1c804d458369b780e93a5e32b8a9581a18457200eb6944343efef4872a03ab1effcdf7576d08357abf14cabb64c74aa6890192fdf6cda3de84010954abbe53ac04683cdc6fa196cfe07fb0f3a5dab0f77d9293d0b2d0e5dd63b8bdca062c56e6f5fdbc44a6b5f6a303af52969c50c7cc1f9b8d077ce66f948285df829dcd4e6d5f453070e2d49aa0c79f8ae6a597166bd71851275f391b062bf6113f5624975e156f9e0c417c4a9bdca5303ed0ef2a0ddc4c8b6bc7d2aaf52a170ee399f19ebaa80f5bc28a126ae071c6a149f67668398f8cdc11e7bde52da9125f9b21cd1c9159797ff0a7d2eb5ca1019946d89a8069b0f5474c130b1c6f9015c369c76da0818c787f01b4f26c90e610f20ac79f0ad7739a8f0f3c1b13982ce426ac9d7d49ace45c20c9e53affc742fdffd562827abd7313617ff04a6b619193f3f97fff5f97e23a116260f406e4ba7ad2eaad9098619c571f3fb815a28871fbbe459acf5e2adfdeacd54dd0dc08be67ead235786c5d681f57316163a3257759886781edbc61c127b99486b758d1331a772d66fd43485d9af7ac17bfde715479b20704525056f2862325b53373c1bc6f58cac6bb7d11f62ae50d0a874455a40394c0077750de601e6494c6581f6d30f7f59b9cd031a826bd714732513b11ec12413b07f9f10da56a745f579326f771da266f318955bd3364151ce6ef9bdd5ad2f24a3e94ea150593037e9cba82ef8fade6bc6ccac0ba0e810c7b0d459445f92d1a485709cc5094402b98a023ab246827c23a684ac64e6021bdd7e1b11f50fb3bc4b6840c16f6363819131787fe36eea09f7538ecd38be4f8bd41eed9bcc638ef1004b48a8efe86468eb688ff4587760e3a0e99512326573f474bb1ad3bc6bbc5e65a4e86162ae5b1f96b9767cd98e14de9ef56dad8d67b6cff28e7524e088a943e670abd139faa24311e7ee3c838a18b420455321f69ad997f1d825c8ba23bc9a16d8be67c759d1c7e15eb28996af7e35d28a6867b1a6a56005e843a65033711642a589838c98b65e07a1c86bec9461a8b456518b044134c2ba4e65ac48e6cc776fa9660e04698b2931d55950d676bac8659a3657729565a6d1b133648b7df9f0445b329bd78fe4a7815ab9d8116a616b3659effc5937a2c724111431792c56f912aa3db14e54f55ee6e7c5c14b2b4cdbe918a893e1180eb9ee99ebaf6b4a1fb0c4bb0e1d5de6a07a5dfc9b1c546e878acef36a2afdb8c2568ebe94eb00f438f28afbc3fffe3553e5897a173b1cdb85ff577acbc6398640f450f61039d9913d0d185578dd389805912aaab0ca7d0b2f6d0e3e7323b1ea6b0aa76c0c1d4f0aaa020b25852a91a682abb87c4ad8ae563e3d3a433bdb3b0ded0e454b048451de103dafcb38b0fe7fb96e1af3bd44cad235c775f71cf58cdfd3544ea0248c66c6a7da91e0704869ada69c9b99449417c8c207f2c8a6ceb3244279f765b2fb08aff1209ac31dba7e7339ffd9a50804dc6180ad43d4041eb7bff2997ab0f350b0eb3447469875;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5b8f7fda46ae45ff4e1310b1dfe581ceaf44ed2f0c03545965a650ffb7df3981915480eefec84fe9cb07655c3bb6149c3753761e26cf1705627a1d9e14d4636a8b2d9703618162bd550d92efc30d98505525741ce83d89bb6331906666a4cc2555a7677017fbc52088a1ef6bcc80294f233ca45eaad274517c936d2b806914a366df846adc6bde3a6ae0e4b1da475acd9dc02a738cbd86c43e0c5187c6a4cd87a529c2540cf7f17c3e1d975888aab6beb10485f1f7d0d01150c810a95570d1f2be9b09fb7b71538928fe50145c4fe21294374e8960ec6ede29aa8f1e480aa47894da60b1996c2d3d4214c0ab02f585439d94f371cfdc030c28031214ed71a06bb7379de1dcf3a49e5c310f5c80feeccfbf6df2bfbe7695a3341bc196d359162d92e21de782c9412377c490de9369946fc85b5e1d0a1ba0593a84e452cb293c232237a692b6d39d225eae99d36f8957c124c5ffe94d2112132af82653cfe49f48fe14d5fa6f6d56d987eedbf6eb63ecdb174fc696d208aa21649ac466b4d1a71942c1122288b69f51240a15f660cb880615bbc330a7550df392a072a51784ac8166114b7c21303c8d463c0d4acb6b21403c9a7757782c7c56b2d7936609478f94cce4ae31271898c179704062a9aac2103b786157ab4e6f8098c755485d3bda76b0cada876159f6c7fb3b4a28135f68bc4b9778a0c5af7a151a0e681384bfbdc2c9acb3ed5379a95f30bbd16e30960ab1e3a73c833c98657087538651e0058cdb963d32df6d672e520de6c737cd869bc6ab49e630e54751cd8598b99a2a541539a049f7956e63c9eafb07155f335ec4d09c990ab192b5ea5bb002489194e0eb002b6a418c43005c67d4a058e225fca5dd291a7471c8c085527b00440acc548e43ad1e8e6d1cb9733be94b369d7c31f011c38cd7efcfadf16760c922641af842454116b7cf7d6e24b4582154e0f0b12d626d863545ff1511adf243f8c8aa51ba18b783a23f06614b4c341a34336a5acd90d4c4753a0c957143c25d2cdd8f87966b2349255db1fa2915be090c912bedcc28c1ab0297ac7b5831b5e330d44d78b8aad44875b97f616d8b7c89f22d7dfa465832684b8282489f7004d1ea70c6d1b33e6d08546d9cc5545472be038cb08c9f4c34786c3e3d1e26e0b5babf4bad86a1e3bd704558f4b17d2403828319deeb468b855e33eb09b6a4f7135734b9965203854eef82e6e6c9765e74f38dc9a3323b55e9cedc66b27d2da3c921a856821c1e417077adfe2c0f6595a92be73aa1216f3d14366dad5e09925c13281dc800a03add4946695c279704d33eb8ef7d7779f73528de0bde5cc598dcd0fd7d45b35265a1116d6712d45849f90b504f7cdacb04ad85b2229ba6a1d5a51c5281382618a793199cee804cd3b3748da6c31448b7001105146c096393842d2a150accec0cc7f71168db65397e9ac779aee21d5d2aa32ee2dbef0c27072bc9dac459632eac07203ad6b236997d39ddb626fe1daaae6844ed11dd29b50ecd39dccc56a4a54aa9bf07038cdef9473f32daacf40c6d358b27ddbbcb49fbe08afef457a3d4b2c4f9f506d3a0229e17d831ae03b0f7352105f540ab4bcd26d674b598f8942c2074a5636093d91e318a3fb37f8f56062b598f2052f7cd99ac1d8648f9bf8b64339a72748a1996bc0284f032f312466a66acb9cf3852071836018535aa2b158c2c76d7ac7ec90d5a10424feb1a07c24c63cac119cf56cdf89c44d4f441965ec781badc50d11f7324ee7a88bd28a1e05063fde07cd463ac34cdfdf1fbee1f2a84fc9da69e2483fc558dcfcaa27f3d9f2ecd43e9a0920f9b9ea606c61829aa4f12f4ec9ab5a625c7ea274d2e5b9f35268070050a7123a6fe173b6da38e9fb683a8d79047c7d37363c68ee1d1742768188de3f45a30bbb42e76619be585ff95f4fce48e3864699f2255e21ffa328bc3913ef49f86517cc38485331dd9d41c1ab66b80bfc351dd90035ad0b3baf9b20f40c7ad9367f4d5c5d65c196c987b395ce97af7ca29479d180aea6b08b32bfccd0429398a7f56bbb5776ab169af790b06355bc145d4f154fd67ce61202b2b2f8e6d3f182260af6f4f5eb4136ecfcd587bf2a042949204f99c6510e5dbff59338c9e59e4f2abef6c34fc4859bec60c6bdda1429a8fbb962dacb02998febeb7237c5e7df5cfa8a9416b14e3990a1054811653967f1fdeaca34dfe7d6902c1ed50a9a1080b75cbc029807d14b08a91914a9e3db3c04676217331bc906f0c565ac13c9dc6b85409e9c1832286b2fe3e3ecdeabf7c0a06263a61b3b0617f9af374fa97d3483b9ea6cbe8739a5e57f24b02e78d0818c7fb206734d5888f3b1ecbd7fc334a4412792d25415075208748c9ee74f34e6e27aa21818654db05538167659a9db9d3613eca2f5cb669a051ed5bb5c75dd81d43b3d99a5243922fa0bde3acbbca1a1a0eebfdfd6e041580b2e09750096c53c2cc4b471ac6159bf06e45c6bfcda07b4ed6e3867d057cb822226428671ad5149159aed0dc960f436350a2f0ccc0d90276147275d534f3533f2eebd450de62e9f839748499838cd500b688a3031fa5e3893959dcb52451f75c2a0205dc3be59fbf2d98208b50cbb017d33efee0c6ac2cbd5b2fb5a6704ac761c51f0a4f19cee4e768596c42279cc7ad7322afb197891c3a3c4c022ae193e433718fca413a2ea566f5441235e0fefac10c92e55e2866277e5b125b4769c081cf623119fef4a33858c433f57d999e6f90e8d06b3a7503a1f29b6c6cc467243757f45dfc3e5451b27dab716c8c4a68b1fe59e4ba6a74c8916d534e02bc9a0a9f5d9c9112b0233ca27c663a7d3789a316e3960dd6a283a251829428715b16e0671cbc936685851c2193334d1d04c83e2534ea0d5d84247dcce514a94260fb25b6de6c7f5d362683fac03f3b9c2340bb5b3c257848645a1ac9b8df10c7ea90b9f08c593c421f91e582bbae60643239d01fe4facbd4338e10bec570356b05932e53c93e6c2c4b83695317c0aafe7f29928490eb87cb1be2e79be039cb692614c22d327ca1be25d5aedf9a4cb6c8b15c1d5126207b790f1467fbc36c44c568071b138a4cd5938015eee13ffacc5dd51a951a20ded257a06aaf518517804b7e6ba06ec161599c3b65b8c0e94849fc4fd863a3de13c8223001e4072390c2cedf854a053e8abc1d98f2982e39b92e99a9ecdcb1c7006edc0a1b6cc9b19d27b9c44089d8fdb38b87e007b10d1c9b6347b03bdd1af9d9a407f961ce612cc7b14ff58a4444fe6d2ff268824369fd9a70661fa7b01636eba4023c79eb16046b640d5e8fc8bbf224f63e549c4950813edd5417258541171fdbe5050a44e5f23e5e3f026ff88abbd9b69e31479cc954adf5fef896363206bf573429b6bed263e953f9bd6010f4552dbdab1e25ccadb37c9634d5c17d5fbf39f0d22b2fa2e25e58ee6062ddc1679fa6b2aca53486f94eb62ecab8a421d8dcb5bb48cf820c2c8ffe1bb8bb2b26270bef7e9b38661734b355740144d1a3de9303ef662d5a7ff9f50623721f0b1969fc6fc151a3addc80af6fa9b4d8530e45a73b72adae8eff6d3bbafc7040f859ddfb731de78bbe4d686eae0b772c7cefa4fd5d0fa212960443ff4598ac7437c068d710aabf7f4e076af1d080556ac7e9f85fafcd61f45f280186465733cd968c9f85ad6df5f4f9b687e07e5675e70aad868ce2ec62aa6148954ea2d4a324712d2588aca02aa5262eec7e9e48666377841d380121b390f5cc3766c030bbb649bfcb8a9456d6647187fae1d04c88efdee7275dc4222741945032949834f81f101e3af29e4a1293091db2cfc5bc911b8c0e838064af6977c372b7856eae83fe617fba5cbce239b2f8482a246ff6aa49d5bd41701fa3f6d6c63cb979df6ae125c1ca2c7abfc8d4f4b7f12f4513538da2f8daf60c6790885177e4520d3c65d4ec3007dfee714635d3a0aaff71748e02cbd127f1ad339b8dcf591971572aecfd77bc93f847dc5fc20a4352d4c7c2398ee4cb07b01ca3da50658efdad3ea11f062d2bc36c4f65e902ca7594c07c02f0b1ea5cf2f2fed012584c237c895485de32d7ced605add43ad704f478a7d6e030391cca546e79ab83d9413df658d071465af5a0afe2b691a625d68e5988336222c5116745a268183b18b4e07bfecbd4714112d0062f42852ae9c1503178f3829b9b3329f7a326b64a7ceaae7af081d3df9d0029bdd77df86c5c0355dddda442defb0975876bab54fef37e9179de2cbe14553ba0ed3edcff492819f722815b520ab8cb4b2b20c11e610351793efaa75d6a05de951f9b0f4c683c3735d48f14e5100896567ac92619ef4f6b57a2751b9e7d4b7267c733f361cde70f3fce34f72316d95d174bb016222239c9cc63eda46309dc47eacc02f3e8effcbf30612b714a65e0ebc17f1a95fd3e137c88f2b2b31327c814e0d63271b39ef7022fb8d24f3070c2b3a8a1cb0d27fd2cc84e6435ac5f17b47f30fa4345995f74d5afd9b36e57aa853e9a31c7fb651f9d3cd187e172dfe04e198b241e0c2ca332199de274b6377925197abbfd7dc4f9c0f7a0b9ee7e8ed0057c05f9fdd56c40717b3f9f0a9f2102ca60ac43c5cc9df3fd09b55249bcee8575d5852ed9af10c617a06175ba33e9f7cbe3ed49ab91df3aff14d032a0c7ebe53855fd241a6afa0c2fcf3f547a12b5a1c6eed60543019683a791e062d148fd5e42be916b3516d513adc0f24253fef464e0297adfe2147bd1f5e2d4e56c508b05a2962a7b7eb467db7d11efdca0fb6ef2d0fb25bf1ad77c69c33d0317a36ef2e598f044e648c2f070534905dfad5d02a6da66b2b3b050862896878bd4fcafa2bc7ca7fa30a11c4ce0a7003c3a44c83c85afe8081dd5beebfa773fb072e5196160d09f566fd1068c04982ada4c331a00cb118e27d101482af8bd00fa647f2848ecbe6b7efb73c3a15e34a39b1796e3464eef79e24de64f264bf39a682368205ea9182f538cb81d1e50a2adc2448a7199aa30c0cd792af4bd7a332431c9457e6cca81da7165e3f766e261a3c6e5f9cef94bf9311740afbb50dd495109be2e5c895d896be7ec52730027585bed003a8e3501a54fa04c6120de73403089b6db3e6f3bdcbd106e6b6d126f3fb16f324ac4e22144684fdac569cb5f865ce2c2471dd304e853bdf53a46ccdc09c7917dcf0783f1dbc7c1dec9941d66a0a58e63efc7c5621e146a84ea79b0f0e7a08adc51d6798c35a33e700fef092f55f04792043a292371ab9bef2e4bcbfc775c343c50401e1af46929a19d2acec0545adef46159760d4bf083f26ba53b1dbff038b540f8b0e272a185e2ac5165c04959c26efd72a75d6a2162fc8594c67f70d5d1442e83ccb70bd78c1aa5445a6a5fc989bdce00efab4a3e77191cf33d3f09c0daf746ddba2047716c431650d93b691cb55dfce0f7cdaa80e6df2703ce09760019ba50a6e83c2fe36c850667ac3bb18599dca8e951bdb85459ea6ed28fb15b169723b08ad82762d57fd17480d720bf9475786fa4f955d3881220de6f71e95b0b08d870211546da86539b7da654179d7143403e1f4902b50e61fe3c47d6c4157036c049367456f9ddbe8349ec00651d19274965fa7677de59368ece0b5d88c8741e5b77de5376dcf20fb82d930c9c2db175dae2d1add1839f07717d5b402c3dcf5c4b9e86250f0875caed41f4b443a1460922f0a382f56d28300141847d0c41a794063f5d8d2e93ec7bf319a3c08d393b993f459817042a1bf9fdbbfc56e044bd981d2eb37b1c9142;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb74dbf0add5c313c0f29ef4880f197aed8999787cfe005b559922874f98145b39de486572b574beaed2a95076730d18cd9c4155ac0aef86d697e761aa4eaa378cc347345d9ea2e25b71bc66bd92fd2d173362e8b3978741aa7078db4e5f448e446a869288e9cdb4e0e9fbf476f4baa51daf8c29898254582e3adec30027674fda92ffbfdd3f7d7291b6831b5c4de62fda5d0cb8713c7c8541d25f79e70838c9b98f1b8b8b5d0e2de6a0e914d84152846e2aa52b782d65f30029355a59aefd841f777c8fd1b1dfed87f7f7c5ae9b26da8560af38e8e28b726e62b435f6d82c6dbda18a516820e3d461d521f64985b220d243887b1dd62a155915c2fd7ee2a6ce5e001d598f42b687918daf8843ad8f55e81f25beb9167c88355aa630dc2b82446b867973d7f4d80d64a5816bf48d3a0a37e435285d3cfd54acffe11fa856439a4d6db1503e2486752f8b14a27481d66fee6d76c57d184ba7fc9f06644a2e4cc3a2b871f6cb029fb5b3740cbc46f0c11c36f0791a4875c66fc811ce0a94a3e75a048b4830a401536cbb545fb8ff5a6c95656e26f1be1be9119a01d3e8614112123190ba27ddc9f9ad4e3a6580bbebdf155ce93c27806e517638b85f11fa5f4ad0ef524a0217fc8d52a3d3a205febdedecf677ba18925084ea92c6f0fa25130994f30941e20d9f7026c464cd0e530490b4cbacc54ce10490a4c83c7aca17af105a08177391fa7c3f65bf9a280ccb67f21a298bb262cbb30d19ae302457f9cb5faaf793c002cc92faf6119f9d331e5d573d5c3eabcf03a7df010f25e22ed56f6a3239d4056ad31c95cd0b3f80f116443ec1a4225133a31943de561ea9428ad32f2eaf9a8a650f831144702708b75774534d709c8944719476e51312e4dd260f0b944674b2faedfd5e2b861648a59a4f50221dc6dca50ed372262bcb21ceefc6653ce52cd0cb39af86a079acf99df9907c3cb580c1dc40c13c4381dcfc65eecd37852075caaa4f498eb5e3b558fe10e479a8194785b5c06d81687afca56d264347209f7e31f1574a3c5738003101ee84b1ef6b9b129da6cb6cf7a84c02e706460b205bfc4550d8cb57c24470001f2a05b809d74832742626bde5e3b7034c0e3b5bbc74b3594b7635f3deedfcd3b2ab9b59544df2b6b4a9b12544b141d71d0d7d906d5ce5f67ea72263381bd20c25c37e15b8dd487792f0a934e5763996ae38a9c81f1a800216bba0c0d50dc0e1a23a9fdbf8fb759dab509606d107fc45c75c35e08ad07e943c48fa1a4307c9f455b6fb4766fff790dfbfc9f8b5d422a12c3d61e524c1b725fa27b9092f94bd98216289920792397b127e9eaa15cf2b5d07012c1183912eebf816dab95c0f6fe85997c407e166f7909b0bbb1d2539967240d2a701918ed2a9e9919a4b96833b9e3879debde4179d3008f38e06c30ee79d0520f11dbd9fb467005ce5c2d48d15062c7b2ce36cee4198dac9ee731b042df1ee179b0e08606deb1b6bb01b088388a3f7b10d39f5b0c36df79fed44335fc7cced730580a1c433ba110be76ea9460f777ba4594b5ecdc594de390bcb1a7216d905bb69e354132f4b3ff989f80dd6f84f9db46a0485cfa77cc971608a9d03e07585a5c1da7b39fb0fdcd78c69c49a0347dd4080d4b91e7c6e45ab883117a7545e472ef4b1aa405b48123af6e7836b2fa95217fa3f566200f5790e3dd16808011702895e521cd62e389b79374d08a0119fa1692e4f6f4adb078d352e00a7a7770cf1bee95a32ca3a5428776bd3af9388a488428443706b20e1dcdd0f44089118c58ba84f561030e9eaeb458c8222f4576eaf8785de95e0a7c3a514243aa61a54f079b51befe0a2f255e0278c4b3a29d2cc384afb404608acc16eb323cfea00b68beb14287467416f18a5c07f34ce2b9b2cb0e0551e627969406e95b4b974236c26352770f2e05ef2db64398677fcc134c7c7c53961846e603877a81cfba69fa8076ef29de9b4095d87348518328aac9c6f44b0ccfcaf4f9ebeeead4517f0e8ccbfaaa0989f2764de80207f83a32d4c3e05d3e6d0b4d38a820bb72d69b37bce3c82e61e68b066b739475794267a513b2edaa23f29642cfd98493c10a52879edb1090ba41b600325422ac0dee9dc96f031cb80ec7216a4107f8ab7facf9ec69c385535afb26f8fc39359af49b4fc280420d64395528a1b9c6506f8a9ef5e2627de0ce0eeea1756ca4dd085a476457dc6ec7212ed5517d1d2da47bca1d935bac869007c2eca83c0177a929577cc8726b651bea99a673f34c7369783dcb24be160e8802cac3bc9905bee23c580e0162e880c9c74ae32952e38c4c9af91e038ed286dcb3be1b4060c98266f759244cbce070eb44dee6cb03d2ad043ebce188bdc401044fb03da9016384a10b0dc89cdc505b22b529ca59fc04fad92dee2df16a62eb75c35cfb977302126a481aaf0d48d618d66d9b9ec44748f0dc980768e2303694abc181a06380ebc8b4457dc40734d703ae46f27fbf6967d3390708b218f64100a363dc4492f2634a2efb9732773bdab80c9d37c38d00e0e5bec1bc1aa92a085a0dde93011ba9b98ecf94962e266408dff8820f183e778af9fbd43e35c05e295b346e41659e9dace9e9fbbde002881f16cd26d0150e9e20c1fe8454ee6591dff9a22d374eb3a66aa3443be58be6ba1131bbb6226b9980841321df3d0740735a2448f04b493f87ec8657f4a11e3d653dd0b125ed5af20fe144433bf6c67e7fd75b62a9b7529996970fbd7efafb665d05e846d3071275a8fd42113d1f99def5a47993d1f64af7924a9f0071106331a41da309bdc07504e73689133941f9bbf7c92f6f35d07f5093433a7fc128e2e1dae39d90613c04579d999d52f0087f0b12a82ad958316753d99ead6202222e57512d16e89c17f1fa791a409f581bcea4c66a469c0df20752e120cb1fd1f44736cd7d45aa2d047a4661aa66f68f1217469eead75ba3bea55f356e385935821ca3f1f28e6d9c44464c839192d6184506b578e1074f61d15e10f50d8998e871c75ac8023cbc5aacdeb6eb7b90dc053d7e137da2bc59535be02adb41f967cf3ea31957f97b35df147a8e6af2a8cae087da70d3322f0c1a60c31bc8764334cf26e0e3a9c5a3c4fe356ff1eb3b6463ce57498dec5c85e5412e61af10d34996d62b741d04e0bda7c427318699aae65235773591876a44881978bea3e2386a67f49fa5c424eb04bcfd2c7d04c909b0e382bdd88bc501b1fa00c0c5e7b2aab382b06de6f9a4a47128d74521378f9b9250bd94d4a127306a76c6757510c929b984fc648ca15cd1d4745a1daedaae9e34b16278af07fe6ddf977e0fc52d62de2ebc5a8ab0b04ac1167cbd771e0b939456e1f4aa630c30dc673a238d83f9f4d2c8c703fe6a06e32293e1bd3aeafc716fad9532eb441a499ad54438978b9c292f512b8f0249e580e30dc0aaea75239568faefae22e7e2abf3a4aa53f0d14b8e13aec399559e72387ec443f3dac6b32688be64b6b8ee42904c1fb9dfc4cfee75df72703e813f8725029dea74df99f2a33a4c651ded9e4ea99a89034726836bc738259ae28ff07abd4984a27112ce7ceedb941bd8ed25a2c4a5b248285a4f961b7982b6854e224234b4c3fb3762ddfeb67a9d638b76eaf11fc67f28b1393d5b35a56a4ea7a43d503916551d09ca458f91060a6c8325dca3a32089fe141899ba996adac6e24d85db62a959ad5640e6bffb8e5ff12d26ed159e68fad6fce393de44a08425bf2790df802ac6caa8366ae53284c34177e744c73921a6adf251fcfdd6ff41209c8f2e3f6e957a0c2299104313c49031fac3841451c9b6f8533d9dc6b0aa74feeab28d83292530f86bbe08a0f53e21bcb8b69f8eaf00f389e81cf7941ce24687d890a1af433ab103014468f2cefe4cd25a9db2058e07852388a6d86158def5204d77539379ca90ccb956d73be49f3f9d3f192203f624a757c50ef5b4438ef87adde073a9e36bf8b148d17de80dbfef90e0964203ff4fd83dd345cb4f9af4c0b5679239aea838677f8eff903b6bb815e9e90a861fbb61692ccacde14ffd9c29d636758fb650b31df6a280d1fbd773888fe2d8073606fa55801fa3272dacafb2793449991e294fe60aed215491d2b7b96726ace01e8655d48b0513baf322993a3e2eb4c9476e537980b2c78a8e4713d67e21cbfe58edcfd82616c33b529198fe37415b9a0af85a52e17808810bbcd69cc59463734084f7f4cec6ed0316c3dcfb3df8aa838d731ee95ad38e1b17f4e9801b5750c4d0327f236c4b4043e219caebbd11dd44b60d94de4b5f66f8d67921c9e2ecccafe4ef0af8045c0dd66a3935ccfddb3bd1067b986ff6cd94dc9d9bece11a4bdece23372e33154608dd9183833d3aa7c919bf46004debdc13fb9c9ee7f4ba9e4f94e9a4ae9b1a2c5144491f0cf17e9a6b6f4f8cff0a159c51da775a0224e63b3cc21a980896fda23cfba457fa578277d460997f6ed084386b0340f1084f3296ddcb3b1aa7236d50287cacdf6d97fa38d364786949ba9366d573911bb47ab0460ef4ce4da3c854317fcdd462fddc89a653aa3d1096c0d734efedebb0b6d485421cf8bb7848980cdbe2ff52266d04626471bf5594fd6672cefac1feb3a9e331800e32534fc37d37764942846971c5a8bca8ef8ea3ecef6b75183c5dadca650aee5c2d8185f7ad65f050faf5b4a6a15e6534089f96923d0cd3ec65d6ca9c9ebc7368f89a82807bdf1fe8bd98b721070dd3fa6b2cf516446e9e00fc6554c32289548b0b37cbd9dbbb6af3d4c30b59ac333d093be15ad60355d970013c8e69a73ef4711870158c0674fc7b0d814a04e7c94fda55efab09596f83eed31da4471561b208f738464a73c5eab74d9be946e3ad2ffa08c125e3f13801fc030a84001101d05650f8fa55da0cce009ad268d6da3e0fe67f92243179447c146b32376feab00f46c387589c7bba3645dd07f240c12182a8358267d6de7f6fbbd4ba4318246fa430bdaf1dedd55381bfde92eee7e1646fec256025dec848e269b3e3f5ed4bc81652f5b55d4c3fef216aed45e691f58389789c5a28c40102d457fe25b14d8bef4e175c015b24870626bd2d288657f70f1f9c089cef943460e8fe0cdf4425d62a74486d26e28ffee197180aa69e307554aa4ffc5f65a207a4e967bad28f8b15563794ee4063b6689a389783012f2a9237ec09ad08ce0aa696326941495e940a9e4ae0f013836942bf8d7984c2aeab8430f051abe257d3fba991f5fe840c5f06929a9c0501a77520199812a10ffdb24fda47cfc6e19bab2c24d3bdd299112d7b0625f58b48879f56e416647d73ef591c9a31654d96a4f2646e5ddc342694672633baab7b4ab22a7a4046d2a5260842c0321db456e5b34a30f8498a09b29b2daf07c5911b24a6c263bb78591c6098cf608ee2589fd9f23d6cbc0f6eb157296cabd904c988309cfc4814af1d7bf50aef6f9ac6557ed380ac2264d1223587bd20e0eb45866b3761672be08609b42405ca6ddd9a622e6ee24d9fb8a6b0187e7664abc2e2ddca319fcf82486da9beb1d687fbdf1079e3b122381d6ca87bdc85d9ff0e677df4bd9eb51a2e6ba45923b21aeb7da34d4bafd216e9cf801233ebd651ed10384f16704399382d6301e3495da67c23d4ffeb485a60aff8e73a35de82dfa0263e2ab14e963375cc36c75308034121b8cd6e356edc8447ad8d1e31eecd280d5716c1b181d64ecf789f0cba9264810bcc55ad5dddc9d67566f4b9687d7271d3c885fd19714d67cbb1396c4144be6a4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h39f793a4953b4d3fc62944e568d4ee275a75f4ad1e96e153c4717c9af489e3000996b58f72741b4344f305a816c84f23e25d8e72139157f2835291b29838cc706b067edc1c2011f1139d79324b2bc3df4704e8ec0a9d805f018e376e3336a11f1b9272bcc2c19eb7fa463097ea3078975dd137863672502f62408a3ba8579bdcf6b8ef6535e9a3cd5c93456188105f08da6a2be7d290638b14615bbaad04dacc1ac6bb3de1f6bbe642a5a674266beef2455945ededf2007bff214661f87282a3a9052088b0bbd9f0a48cfa01f54cd26e0ff2ff655f17225f7f60dc445ff71603af46a0cdf83b62feb1a1430a686733c17e59fa346c4ee68ec347ee53144bfba7342a9bed6b49027621f3a4a911bcd2116c925b20eba47ceb784fef218c8338644b1d2955c46cfc83b5004e9aa40a31913138a528346ccea78a4b143c5b601ea67dbc1d0d82829c668509f7d267336ba52ea59260f0685a65823ff4a4d37a9e4f18c4c6bc2d6da934bc7577b7ac85916c54eb3f64cdc2c643a0bc520d84076b857196c40a35cfde03c9a28c982f957b87af926baa380553421455024b0558a7f739f7631b90a610a3a557243d7fbba13cfe1f8ae2e1a33985f7116a2688c5a7804f3ce5efa4fa7fc8f897da3201ffdba1cd8511f58825e9c410caf8e4ae30ef75cbe903c609ed79e2e6fa38a652883339e03ca1f9cb5d78c9c2b71a7c47207a05952adb3a71812ef21b61e4a194f7aa5a619cb3f829e6114a8dcfeffcff7eae6760578f870a4d99037d9629cecb92d684669bc829d5d3fc411c59cb5e6df679c99ce7de5e8301ef9eb20f368b42b79ec15d379bffeebfb5832ba78b3be0ee3b1115b1877ff42332e54423a8d8262b27937fc30974958ab1f78046f016c9facda19f50807aaa7e89ed6ec7f20dba930dc6b69c893981b0bd0db85a31aec7422a65486aa171513ec3e6486ddf6083e2a7e6d845c90a7c31e441ee5d1160fa3448a17e7b895fa176a40944ca0c5529a502f1505305139297172df6a3444f99ac9565293934fa9f242de7339e5a274fc278df7189dd40f3015e041f78702e6deea9e13a19ffd4cfebbaae5fdbabed02ff6c04acbed3bde6c0e78f006bb8cb027c82382ebaf0ed3db20752464d7b37d29273419adc1f5ff4c260ba5ae64bd617ff87216442dc85015ab31bfec5ce9500d6d9fef6738a9f7e58e175331eba72cdb4ca4178ad64fc040b79deca9c4d0e7c984431666d49940b53d62c6c324d1789d3901239912d8b738be8789c709da30e1c57453ee6f7d33e835848b199aa54a5a66e77799e66668cc1767af46f5bcc025fb4da20563ba0a37cfbc0cb26599eedb27a4ab31ae95798232e7f0966be7982bcf217ff5e010510f73b9df427d027fcd2b47f77f41307a78fe1792579d4981f0688cb82360dc687a5fa322368bb90d87730b56d1e5cfdd7fb2a4bd3917167ddfc09403a922a1ba2b4cc198ad173bb2116f80d026082028947a29743deb8fc5ba6df6f2af92e1d31cda169df6970f3694a2d7ceecd73575976065118f659c9b1d11c165b4b02243cbafd935c48f219380ac85f5b2a2263ad46b559c8b98a69491084c4b132e5b835fb030ebbd2039e69b0a73b5a0a40aa119f566c8142e86f7ecc0bbc0992b72e45fd8b3aed7225c82fa7ad329e857ef4ea6dce0a9a7d59ba8481886211e01c011fda955bd68c1565d1a592860e37facd02b5dc2ecf80e23fda5167deb1cc1408a930ae224f627d58a4e5463ae7df4ccfd885d6fa280d057e753430f5f1d4c82236684d2ca5f1c6a2df97cca33e27b0f10fae46743ad5ab504333920bf0bfda2e2c1e32bf8cfe7e129d94d0c4c4e7c52f6cdec34e379fedb41b1f18652c163320f9475f98cd3c5978cef839257db184f32a58741a1812cf66ebcbb407820c874fa00db7cb1099807d2f0a2b40c3b2b80f17494e71c1baa8d7a9083a90aaa36b212a66c905b82967ce801a9b69589038d4cf896bd38f00e3aa0da4ca69766b36a962dc6fd03bd59913d3f9d58a1c93f63d2bf4d2290d534968b32e542372dcacb4d48206d55f6c497cf99f248a624faecb1159de0847603c319365bf76497bcde2ecffb976c6397a95dec4f730ebc1e3948bd93e3db4f1a9592ea668f39ffbd438ae785dffd40cac438a0d4e1714d315a92753b08e1e27006915e3332ebb82f7a899f68d9714f3ee6086e2ce8c9e8cb9122abdea6b1ceb14b5384c9122348c88d9c80a59a8b6503d84a8367617816521d49251ccac511502ed1d64f24ef91bd5c4bac186e882bc63d7d5b918745c2a64eeeaebdab24f1ed12ff314ec631183d167cfc4f95b23e7b9f7f051c2f31e70bb9fd257d9095a658c72c3b6f60bcc1ff9d9fa348bf506a1071fbde9b2891fc111d0db157af68d8205869854cd19d6707cb6d171e46df13671c0852f79e6fb6800e9482c4e369c3f3992845f2ce30338d6727fd9671e0305b1e0f6fb892b016ecc48e168071ba3ed836d1588eb7c60aec2a3a59225bcce64c3c19ac182f6dcc463d7e77c052ea9be46472bdbf77e3d5d6c9c1b5532cd8cb9eed400bc3c2f552c40c1a501f18c9dab28bc2f7f22865c436bea49375b50b26c547c79babdefce1a9ecfed1330775a903152002e4eb293dce1bf2c3c13998dfca72d7a3fb44c86038657f2766bdc3c4eec74444d437fdd1940964e93e3b94fa99acc0f840ee9c170f5b787a385f8953969f519ff2f1e8ec0aa17bb46870ea25dddcc5fe5992d8058355f9c2c47aa23d2314a9b2ba1aeb8eace01d1a3ac24499771a799972841b10f18cbf584e80748aff70c19b926eb408102284bbe80a95bc0f6ea6505527e23291ff82dc6f0f1bb4ccdde6aabfaf111b5a5ba8d709b1901159ec993ebce2ba3657c18b29bd128cab44ea546aa9cc2bb02efec0b1a2b295b723cd0de42f10d4e8fd7cc3222aa7d982a832849eeaba2027c2c3187d1713a48bd2e47eac4c8b1ea29adcba36005a31ea5e173aa150cc686a29d0cc82fc89e2bc5051162903c7b50ce1281915fe11dde5840294245cba43197aecd30da175fb81108f68ba7cd179c3ac218d601f20b52231abc7844928c4bb820a5b9d7c331e019079a4b6ef00d3e9a6eefa47e113a3edaec04abcb127dd6b09038b5f3ff9d8642c0dbc982b1e88f07906b63ef0c5a133005210377d07f1e73422af5f6d86327ac09a3c46b2c2ee727ed288393ffa996183d0fea97f5fe2a991186c192091aaadbb48f17aec58a8222810fe80fafa4a20f123c2370c75d6a73b417649d465b64a26a3ad84042f43abaa40cd1abaa0311f4367850f09c9b0e822ce28c4f638c2fa26924b3003511f4e1af0f73e9a280e1bf976b8303f2c4070bc3d07b29d9cd4c29dc12c1a3e1ae670e9245bd5e03c9eb9c4f7ea3bddeee11a976e12a7fec2e1ac7533044076459a5f6804f590cbd3e6e87a3c416ce590e702effedb1c167bdb202e2b1ba68360bf23a99368fcc639a39522feb59f2cccf54983eb3a9b80a32616c316780d6ea0ce586b8785492d8334ac8afd493b4ff9670f311d52b9d42483559fd886f038db93220844649d81563d46f07a01b1ee15a2ba11ec88ea2c18cdfb70b4937d500b1e69189e7ddbd4b968a0c53c9bdbe92831a9e5ea20780e6d22295f0959b5e3956fdd808c55a7ddc0480cd6bba6b757f50979391ec7f0624d0fbbfef46831f70042dbe977362a2054dc78929e59fdc0d93ce49e0e56f66471e0c78380ae28658ba2645ced8615c2fd297436d4747ec06d1059d8eb7237682bba5482fd2364750ccb584cf268fa678d78a2acefbd00db0b3c920f11aa6bbb3b2994cd40f506f77237b244de016fed79da1f1e02eb4362ced98583046317e1d4fc6e6ad802f5d97374c6d99eec1d545498f76da05f2d690278d33fcdeff93ad842ddc63b88f80a7761afe0d7395ab0ea8e538e0c7fb8058c6f6244951f59281335869cd4038fd08789744259092df3945314fd5981835dabdd11d63fa789f4fd7320c2f585db04c3c165b11ed624c498a035402d046c192a9c8b75f8f10c10b5577f9120cd5a1a027c38c2a08193a88c36bee3953bcde91cc9bb65576a53fbf149b639b346f65cd621a8b3fead2b97cdb92eb6562fa2a7164bd33928320ce83d1dc2c76b5536c3d6664814b4d4ff7bc4468709c376365f5d03a7919e999198187576ddc6fff572d2ee3e8ededa68fdd9eb730d8412bc51fdafd4ae7a934ecb9c2089bcc404874c4e8930806b34833603552bb5496362538410e80bffbb94d6fd50593f66d6dd03d804695efa0ab66b86b7870ab9de713fe330f1695127f7d9add2a6bcc2a10f6f89b551254870198c1d4753727a3e880524f1fffe164bbba84c6b44c9ab12c1cb0a57bacbf8359567939ea018429a4dc8d1cf8838f0fb46f27aaa4dd614c5d898c934f981787726bc835a7a5c9836922dc35a2f07705d6980a790e32e3e2ee48fb223b198341cc462eb21f66a9d712e482bce610f5291ddbc2f15ab22e86fab2e115f914a9fd0a09a1cd5eaad94424d2611f722ccd78493b09902c83c8ec9a1be2be6c678d47f4eedcdeaf24379ff0780392a05a24a2a44604fe3f005e122786e7b51e5bf9b15cb4edf47785f0c7adf9b8919437dc04721fdd58a1cbd9d468da3abe9dcc3d48d7bbd8d8bb1323234391ab4e8cce6d708fdcb9471dfaceca6010a8c1341c07dd5bc1744ba749100164aaff3ddef19362823cb255965df8e233ff1445ab360f55c9461d939a858901b91d86c8312414790d0787b7eda6f6df97baf925a2e1d615d0d0f847bb6cecb0f5e72c90e80c2ff283d22507f8e1de81a3ce5a533fe524850a7e9d1d04ce70614bf2429757ccb144a13a79b549f9b6f581475e02bdd8851ec15a4930455025ba65c8a9418cfbdafb6a8e8e61e9633b2d18b0ef042e514c375e579429123ae8c44c26db9682ca24c588acedbafdae0a7b244684b1a24ee580e9edf2d5a86d5cdce1b67d93b20586448d19e81a161c1f418c3850f6d283f47d9b8c3757726c881f86113488273693c511d960facdff264784f720cac3e8bce03870a57c3c4897e537624b7daea428b0279734e5c4f212bf1aec5f5c4855c49f0fd04be5100354022da15c15e7def48c484522eac53712d9bf0fd942931ca285034f2241170708f67b5ad84ab4c9b1705a8a466553b26b1e4a51db857737e4824784df117c5c5d42aa69ce78a9018998923f8fe0c76b89ac053d0664637c41b1e322176563c7cda80e6723f129765ff083874e4af3ac8cb9d978aa59917f6992aae11a869f003959f9385838560076d31194bde7ff37941c986169c530e4bb8d95efdc29a264b30c245b218e5dea1e827a336dad24e148321dabbf73e670aa4abd337a26b2274a6ae6b157c8f59388944360fdf583b3460b8c997c68507152712c9a1ae18d1d770a3c5b73dc920a23f74261cf94ca597bb2a9a21d1aae6202872aa4b81c0c7a0fe7e2cae2595b8502cab0263cd95493f7bfebe9881f621c05eb244ad60a363b589c1393ab4d3105ffd60f4421ee5605325fa265abf19e1729914197652c034525a4d14c4ed8e83048bb58f2b6a9c9d68095ae9533031deb7fed4a3e2f56643388727d94b38f442e4a9f7a7d28b7f5bb8f59bda4209923a99c761191d9dae44dcca36500fd4a576e8a47295da716b0fe35d36f61dab6ad6c1711c69770c575deb499e46fdb8cd0aa81a8dc1ed971cdea6e7ebdf8a778b24c2a3ebc1c699db871bb3cb00c82b9ac8dbf7d43cbe2ea0ad5f845e637cd5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h50cb85b85d5b28fe6db5e9243a09c600bfb66dab12ca347b8eb450398f7ac46e3391a891eeb7c0e5817ad29cbce83d1873d8f3753a33fc31c6a3d85513ce55c518c5ab669d07ae0d300bbda915e7fba7b66c22a5d3645b84269f60cc3f7515d5614ed5c25e41befe1cc64fd11f4f95a8accbda58dd33b353b891e84619ec5f108c5692b126af31873121567f59618b2e465f9fd3569b187c45e29383eeaf7b86b7bad2dc46e5b2b96cea5b3c5b7079d06e4ae3acab277618969a7691949d41332a7a150c10d06fb6ca2f5cdc0ce922875433cfeea09f42feef58f0a6342745e78e727bd9caa8fc77e3b5b5c4717d7814a288b1c0681b94f697e2510ec2583ec745ee56f471c34b4df5a5d5bbc0b92dbe5fb53260d0b864199c10c05cb5f0fb23c9a027de842018f08ea4e337e7370acc23f3ad887f3139a10e305606b9a17a1f966d26e96c7e45a162dc430c3b1c7e669485b33ffa3e27f88c3c331c6d4f86707e70d24734cc61ac1d5a45fe6ab6503c2a254003dc9862619366120646716c7a6748bec63df2688d004f93d2a883edab5781d02b9f5d21fa26e5e4120d55e90bff255bfe659ec06067724397bd11becb96db0917ff7fd25a9437492ce616a161fe36c77bdd4f3c523ae51d075d6a35d7cb157b3f51d489bb1ea95240098ec71246876a2a003674649b7d3289a3bffd595753dda258c25996efe7928e49ba89b7e4a0090f7d37d46377a88ed448d835b49f2b79f946b07d71391b016ec649143f966ec6a921688585291ec833b902751e97c2f1f703de7542c45ae23abbda7dcfce5cc9bbc4bf8c5a710c67799eeac2af1303075e65a391bb9ac699a00bc7f458b310c0baa2d9f0f986715ca627f180919a80b3ecd4059a6ee5a2a4b203cfcf3b1f93ffbab4499f6b96e674f06dc44038abb9a546ffce361242fa5b0892bcad0f904a5ca582c77f5169a2f87aa62bf652513b25a17f8fc9afd3f6d336f875429cf04d5a67e40f57e375dbb6c89ad932fa9460a31471f6308d61b007885445ec3a23f624f7fd471f63b67d7ce8cc906c6a11cf9dd7749fc9914155702be492b3336455ed565ab4b8fc9cf0604be5cbc22980c45acd786a95e46fc29340fa0ff6b4bfe90262407f3388f9b66743fc7afeb93d67f2d655989d4c978421e48fee9d8e23ea980921f11c0d07e9f68fe98a793aa43a675043dbc0ed860e38688a90ca87ff247d9cfc64c01cb1079058981275b871c25d89579c29affc0a8b36bdbfdfd9406e021bc07f3429b4c4c3e7c9602456cec3ad161af96b9bec0b8836866f5a5ceb7047a54fb6d0c64f8da305a836f295d9a5d532f490f3d53597c8f39145836332aefaa521a276c85ad9313e48baece9a8e0168cd6f288e598037728b50c38589f0f81e4441d0a8dbe20bd74695a2e4db0d6c626d4cd4846db151dc24ef902f3645788d69c1cb3c0570fd53a9c888e104fb16f07ea066f7b06d9d7abe6dd2d22d13a0c72fd7c7c61cb3c2534f6c6f3dbd9d79a93781398b03ddf8018cf05b4fb2443babf514743f8deda17a63ec6c7cabcbc7b0e7789eb63a34293790f1289c52327730fbf653d6a125324b36a56bbc08e8913c3b5e8753dcf578400646e7297f9d322f38b6e92c0ff65ad9abcd1c5eced76503462946659bccc1760f8c70f14c0a2ab24122ae2cf195dbad23097b5ad7a451398ea1baa21daca4d8b47b624a38caed2c925418e5d2df3509db97b908ad9222d1d4e6a8f81659e225ac32fabe0c605756a2b343e75dc1a9bbdf35e1406c85c75e7369c422fe2b3dc504dea9392c4cb303f6b45a2ba72ba3ed51db198af7b2d320394debee061c7b5ac2469bd7e3be275a54a3b1e9a910781f8f81b806ba0a89e5d01268816862451e3eeaf6109dbb73510fa7b1429e18231f105833ef2ee9edc17dbda8631f3a70ed8a565dfd9dbef897d7e437282543b3685eb3594d2e363dd8ae7d48c79ab454821980d672cfd6e3811b26d30bc290c06343d8cbb64c922c16f716aeee8b0d0edc2e01cc41f7e645064225bb66db1dc8015c7cc067686dd16f5557b9438e404af4d46e026c23d9c51f23fe2791c637c998d5dd015f6f9965b82d33a0f08b6b8cd32b8089ac34d642544aefb3a4115dc033109632ce3b71e1f573ce142306ff1377a8e79084ecc97ba7b749865ea321aa517718f8e7547fc43191583aecb9b7eccefa6f1a08143ee1b488b32a64b063be7755ed62e7ff1a576cf0a5eda4fecc915a0bec21384d4311d4be3f7c7fb6b147cdda9e0b28ca99fd985c2f24efbcbeea584f3d3622245a8dcaceabf412ad7e89ca484b7963c40337f1388715da2c6cf68e1e13d77faedf0192eb4890fc4163b57e45cc3972e46d6d48efa7fc9766fbe3c0dee098f3f748dfb0eba430215a1ea3340b5b1a138e75e9c0aafde263ae4e41cac6af3ad4766304c287c6b78d96e442d1f91f265f71c51426c5176aaa274e337774ab0349b942c6a3f9908207b2a40c0c181f4493a264521ef34b21bd119888ee228dcc9464f507d161affce7f073d950c23362a30d8dc9d1dce606ccbd8b1f89c84afdbfbd1dc0ff71a71443c8faf4bf2d46d8e181e44c75620c2becc8c1a9f6584c761087cae72d5e18ec1e8648037f6d21ebf2cd70cb40b7458888759094a79a13bba8f4a43b376f7f4eeb8cf65384bba47db913ac449f99250c047ad37e6c64925f17708d010b0bebb7687dfbcb02a254eef96348894d17adb16683a8da2e50d0619a0e6a1be85277aeb96173af330bf96f5cd125be4fc819826543c36f3691b5d3edaecb97ea02bbdebc9d6a4109449f9e9eb9828e11b17aa84c15ad63f1e03938ad74fdb5bd01f8bde7c6ef684fb896953dce14aebaa61316e9847ab7da10f3c3562431e7fd7a187e555749c487469b52e35b1af882384506cefb6eed4c94eca5573f98c4d2d868e51c6501ddc26f7de256d27530495077489b3f6a1107757d83a1d557d589e72ab2fa7e0be6fa9769c537fdbe9389cb4a774b2ac90421cfbe8dac748681497263622c902c89897347a0f47ad6efca03c14b603118d8c045453fc9c1e939ab0efc7de70646950d7a61bcf714d42b81967fdb2e8d6b6aa7ff646c7b6286b463640ae5299a6e3820c252c915c3e3da28272f3427a920d7572d18056be9df92046f788ed79c44ee65e59cd0a5785bc7b9956b490a9ee1a5df73de62714c259858fd5db02fce5b586241fb656ab15466ce98249537c4e8addfbddf974c2ba3211f5949e2efba7e2870dae60c1d15d368d10bed53a6a51c1bd7947ab23071b8e3c9d8bd218a43bcaeb650dbce01e5ce4567c7325440c6c3ed7a947aa938e2a01e1fc02ef8948081053a4eea745b95353b8b6e8868d9100e975f9b9a8f32c63459d2d16e0ceb02f81717e1dbe5142c77d1aa0093f1eb8f56477ca1627e9832988605a0b234ec04d0e68d130607d2f9c10a873e94fd5f93e5cd1bdaa656785cb245bbf0cf088f3dc757d7000a18d9fc616aa8322c5dc903302f091fa43b1198ee808345e762256d9367321ce1241869fc76f8233fb5601bf1fb0f9a441dad911b6a7ca9c62ecffeffb24966caabbc99f4b7e269f6cb3f3eca30f47d51961f4be50df7721a4e30c50bfb94252a7e2f03689e5d7fff4bbbe49fbf317e15741c03a0512e929e270d3163e6ce50f20031406679132742dfad3c39591c1d8ae9586d51d9cda37c65beafaae437d75621ae9d534bc00775abcce3197125b3c2356abd995a83b49f52d19a3fd0bb8d3eacaf21de3a38461b08bd13b7de5c497468010416e4c1d0a4fe13fe2071c2886c0e3765e49cd3e9a5eb5024c048b12fa8ebf905d9c318d3af1cee10d5b3e6af0b333f07043cb7f35768e15426d3abf383ee43308a949911e8e626dd6bb5e3b1e0be5c167fb3409d65fcd3f3b83624770a21dc6493e0aad36f214ce7af6b64c5e726e7ad3a59076cc2195064df29e508dec99246772f98bb769029a7bff72556977d2a5878961486faa79bc3561957bbf908ce31429dbc7ddc80db3fbe38ba3c5ddc73222fceaaa37e4c303540eb3b8c35012fb4cd55fd5a587485e31fa8a53d47efdc050bdfd5dd443cd6ebd32d382378480c70018ae677aa9aa03f37cfd062fe907ef6f5edcb593de3b5a51e9c711d298b9fc6247f0f30f24dfa92861f073eb7c5db9371a01561d1fed2555f6411bab6111f038c2f4553b8af4c4222447165696bd0403b31a27a12112691e90e1eb964d0dd339d6f7676de850e35092cbdf98d1c9e3df2f3298add478c0cf0208ccb074d5e1d6703ab574888906995bae72c00e6ceadab440edb759ae46ec3417c8d6d00d7a060122250a97184e589b772726fdbc80a1f59f60a0f6fcf2862ec846dfd0906d0996efc8cea502de11fb24a8d42cb32073c0e1920343d87dace55d98feb3c02fc1d5eacafef928fb3f8994919ae3590071424a7555f2598c63e41d4f7bb46596fd2534d61686bab4841cea01d1df1753848756b6df8e4ff81b5e2ae5e8d8242504c05aa6d57c84bee4ad8c4d9b8e2e446d9feb8ad9ba1f2dd8da675d3a4da3a5102033d3f6474a1019b6125591c67a40cfab3e22ad4355f2383824e7add41acfbfba93bb9bd6beda8533a13eb40f700013288ced60f7e157c0571f0ff43ad5854e4955879d16ed0234fc9448afcfac89100b359fb3fc29f24e2c1a6efe9a8645097b4a5f6760004d7c205ea793b81dbd773588936fad955cc8d204d0d22513be6e6e2dffcafce464b5cec018d6d6dbb66e71571a342967f1bf1775bd540c0d783c2f49b2e11e39dfff4a573c1119dd380b79ed0636221d32c229ae2570c68957c3b8dfb7d0942211cdf2818a934063867dc3d2ef7d3d9de720cbfb7b7fd4c53efdd2cab70ceffe0960acc64174b4d3d4850f40afb084a269491a26d59bb540b00b031ad6831a671951ab77cbb4ddf5ff9b39eb3f7e72d1415793b0751044e81dd36c1e32102b3744e1b9211421a3ad6fa5dddfd912a2bd838f866f247339c8e6736f0af2098468f38c692e15becf6d6520ecd7ddc27c258c59b1d162546abfef45c388817b5fe720004113b066eed40dcff40e211b3071a23c0ee60c747b2a8d7a915732dfa58a9ddb06d5eee6c59f3a380ab32de3f7cfad9ef962928395494827a3915d8594458748c7fcf72700fa90db669fbd5996b488472280522b0cfcfccd93e56c0e5f62d37b0c86ff35ffc929479bc9ab5d35d436848b4f20e1b81f8812389eca9501382678783a5473fd8aaefba0fa56f52b872aa7c025ec8ae81dde45e077edd62344e18585d28cbb770a2d0d433ee97c24e4729e8714eb8e7c757850bb737903837ab9f98eafc02a5dcc49cf568430a4691c4559a79ada92a3a83c2446b130bc0722ffb6b20987782efd4a7b8e803e4d4e4023db49468d98cb23122ad9482746e919904947a1058069e6a07b4ccfeee12208bf0d3cd9ddcf304dde3a00ad5576d33feccdfbd2e19ee8e3f4bb4d4ab87acae4ea9de5224ccdeb6afd7e5a0a71d049cc51c29000b87d1d565215223fc30b375781a6721103a989fbfba5156cb8bde286a4881777c2146e2e44d37d99797bab7906fe7d4bb92d2128d02d965ffbc492be6149215ed9903a17def2857a548c3787b7c37e1472a133bbbe8b8bb47084a146d8fd91bca63e29283fa1413523a0da63abb0fccebb08a478e8c8bbe6d972202bfe32beac568778e4ab1224bba102a2b85673fea9cd096c6dc1a2cc16b11e92b8917c94ec8170b05ee0145fb1bb96b2ca9fd533fc6ee9c64f7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcff4735e0f6c6eb2ad43c8fe5e663e48a019e0422dfb9c1a9726f76e1b199264c8577af0e65b33db215f2b4ccc1ad75705f308bb65b54ed3c05a2fac3b5e78cf5a71d6f19f4f475a35187bf57fd53c4341147e1911a9e22763b07efc06046713580d8a8bf6df2d1a211bd40b7ec36f8b136457f80f4e29f823ce78f42c611773f1029c047a8fda9f63f8495b55edb3bef66956074ada8c2bce2a20d4139a9ff5d715ddcb99211cb4952471979fffdd3aef042f75dd2b7d658f82f32149dee4b0661a421976209f08cef6047c2556e81d96573b8a191eb3136c38421eac23e5750564863595a6a136d0c9331f7c9ac143da662879763e6d7bf9d27fb0c27359c9d558659caf872af7f971d332e94c6578d92afe924f50dca1b3b9beaeec262630a1572fbf730cf4490f143b1fe239ec66d84bb86225f98a1b766b475bd940b778dd068685082335614dd93b33564257639eb6129e9e04e42beeaa25250598aa0da2bdeface2c1282b4901766b9be15c947a8afb3233935e0c2a844b8a869c18f79c0be28b7779987ae9dcc61270908bec29f3831419c22c555b8f93bae544d5068b033bcf689ed3ca0a9829eebcbd8c03e20639c03183eebc392ec2e46a4ef477f9ba5de6541ffe8a86bf0a3dee113821f1c04ec4e6ded7a8f8017c649955771da42217e305186b3a8cfc716a4d2088f8d6aa351efcd48753c484e733f5f38dcf7ed91f87fedf88a8fc0b6362b5ee5a428a78b7d32a838c9a70b119445d816b938e531a0a964deddb69af8896d99d721ab77039425e1923294484183525b5ec9856ffc0edf35f6a03473583cc2e34a8c03de4984adc5968b9d0f3dbd2b387a8c4523e14a38a967113751c0e6d7bc8ef4729c923810fac045dd2723fd333ccf906a282bb8cc4d2182cf50e6708dfa00fd2603def59c279f3f1e70ad8ace39d3a4a7aaeb740e76e142745a74b0572d55f3d5ff1dc15a938dc67314fab70180e879d7bc1407177ec55c41904540a9b78d08d77f1a01f0fd36b86c44e8319e611aab2fe08ab6ab56f57587b907a1dd27c513ce088273dbea95df18b15d08cab41c6e9d5224a01a74b0f6527af161520a2dae5ca55fc3311a156e315cb0fd632c9bb0b3f106646ebeead29a58554238018525f977ebbb0825ee090a587241fe8c276414409337fc217202218879316ab771833bc359d17a54fc70fbca7dc7346bf0244b7f60714b2bab99855ecb3e060bfd6c5651f6d202e7fc6aef013da1b6e4178d6e451f8fd1d25ae2094f49d50bb2a3c229b627393526546ecc71fcb07d3d270d391afa46b1fcaabe933cbe9e19c7c945bc8649fb89f7680f64743cd3b5e9ee378b327f0a1184ea6c8e29ad9911708926adeecc1634e578532ea5c8bfc34242e77a1702eae78d1f4bca796063d4b0fb7dd1747b6d61ca1ecadc64d1188bd38b99da033ecd6a6df6d2f9faafa406c92407312436188429242d0c9be74917bffa73fecca4463303eea8020c94a4ff8080fd07237d8e9eb082f3879f7e36a99714fadb2c9bdb2682218f021c5dd08315bfc112e60013eb8473a3b39d12e9a251cf5178ae678f55f6827b105167f2ac41c7c7e2a82b28f75769effa4b6735ec53ea01e703e7f77d1f7f5b7d891252e4a066416fcee4172924ece18ad86d4a51e64d0e3aa0af13ba2832a179a151915915460396a2a8470f33b480ae88ef1a4ea115b98c6769d0dd51fd41a728ddd0400bdb34c2e99cb1c89d232fa416c9311df907d3f78874a593902f42d50b60246e4126b33a3f9a7707a28d8238c2a8599efa229d0091f677e27dd01904967b05b523f0fe7652cb3b38300f2d8a162baa76082ab161091f0ec896f332fe1eb0e3746c0bf693dec5342b52edbcc5426d6bcbf3929eab336a4b4d4f3f0aa4e22e8c8870e45926d9c51542fce4df3a78df1abfa3b3be0700aa3b01ca7034de6551d8aabf540eeb28bc881779fab90ac45c5e3ea039b88d04dca29e5a409490b4333612d5d888a9c44f655e4e774914884734c7a92460253d01a96bd12648035804016d561ee5add8691810b59d92d865c25c1de6b3657597df6139c9474ac7b498cffd5c7cdedaf0c643fa6bebe6c2399a26ab9ffc07bd5e7b1e278b2bee4f615a6cc9cedb0c6f9647b0c9ea440f110390521dc1bd8e14ca3b45c567b66c8962da9f2a0ebaa3c3b81b6245eb0c3ddbf03e9003bca4da4f95e6fbdbcad9fbeb4393ab44fe6ce34e386cac2af3dfe2a9d785f5b808a890614e2bcd8cc72d6a764266a926173bf68e1d5ad25374db301a657eedb7eabc865cd41b4f01bca16451dfaf2b4a11ade8f458aac442743235935e7b774aa1389808d29f61c884fc2f934483c5fadecb1682b44e0f008e14007cb7af8d7672f23609025cd27ad61fcfebd0eaebb608af827fb2164bd945abbade92502661b2370fde9e3e4a32cb985f7d5b71b47b89c3bd794be6d4904825e6c5172ab5562fc51533ac96bdeb26fed5e830dae45352ebc77cc5e746406703ab46963e6239774f0b9d53a0e5e0ca511b4d22212fb725027eea3944aef8d7e4bdea13b7de8a03cdf639ef519ce10b62be23cc9d536bf5d8fddedf5e5ab5c9387d8015a33859b4b85fd30f9b52bb52c08c5444bd3b861fa30c8873e0e4536b21d9ec80398b0600259cdfa23aab5c6067ea13e99f63b0e8e01fe9e3423c25a4e460eb5defc5edefe8edd95d15fd2067be5fd1583efdd0da96e2560a8619afe15bedba7d76ecc9acfbe54e895d940af90a676071b02f78952d973552c9604aa62feef5bd3907feef7f0d3ee2a7dfc2551a90a9762d13512f201f51c75e4066bca5b8ab0b4ba1c6ab339cf9527dceae3aa0557c40e93e90ba6f6c6536149c67c7ba796c3d6c7321534d11b756776a70918de76c03c3546b77e92ef99a6fef1028e9a25b716bc67591778ee8cccd9ffe51aa25f30ddf7a95c23f1e4f8489623ee214fc9f1bb17e6f216f58aa9e6ae6a2dff06fb84c1076ecf44d02a344ad7c5e37a3debb0d45302884fc371a5ecf8af288d7fb47758c2da0521246a894a40dd77cf185c37eb336187a9c8c91d1101b65e117a335892253097fe042193dd1986e27808242f15c6a0308e103af67ed1bb7221b4f3d4ed89f3bfe9ee37f883e4ec45b2cb1a582a8c9e9f331377b6ef32131b2b091e506a2b219f75880317f8b0197e8500c5d6a26f4a7407a0920322001d928feff71677eaeb347558db22964a121dcbba96f96ccec716d9e086023f94cdbebadf6fcc7e8bf49253cfa7d482d5963e0fa3d5480f43cd0fc78b46224f6005f52403d3400beb5da106c167bcc7a3603dbbbbbb5664b6768d71b1be8f8aaeb609a21ad11a2a579dd4d73820de259198c014ea19136cedc7f1813f60dfc20e78f4bc390d6df04fa28bd9609532134f2887256b803f8a4b7d7a23d1f0841ebf03cf396627d11929b1f26c70083b309751367a32cb6ff1b2e397c9dd840f942343a6ecb39fcc7a3525fe694bd254ea16c963682e4fc3506a035ca5606d7401ac601a34e4f33376f8abbbd2f7567d45a3787fc463b416987401d14d90a39ae1a9f1eb7d60862e76fb694e8e28e813b59208c9ca5f7f75b7f3949bc89b9c857f0c930164129dee66cc47854469f7c6ba22f33a73d7608fd530d3fa1e0d63e2c22cd81ef47a8d05bc60f56f674287344210a4adcfd1e0d3433617a1861f3cf62f6d2013f7100318c207cf5d1b726b9846241f8f181a0959b5f723b2b7df8fd8398a4aab86bb78c9792ec4000afa8ce2b29d91d91c526581c7347a04ea56da4b58107dec262e72fdb1bd23a39dbf87bdb530c12de90b4a065e61b90f99c5c0e1c6d3045be29e33e4a5f1a843bd1cfdce5fd57ad3b026e7ec271d8b080f8f9a9fa94a7e00e08ff8899ee36987504d4c8ecf0aa16600f86b1d21100fa294eec624cc6575d4576ddbbb8950e19a07b86d79530077e8448c1ef4de2fd76a1c4cbb9f0c08456722ba81fa18fd709b714ae0d85f0a722c77d13b126ebee48ef19a6aef9c9788103ec06b9412cf3198680857642ca46375b9dd4f2572ff88d6c7089f19738b9548f09dbc94ccbd5c0b49649cabb8859d06097bc9f0de5b690df6ad1f2a20e004f77106bf668b0ac0785290aa7fbfca60032f9326fce71465d80e6a55e7093b96dac16c72defa9300c5c05eb90e26731c5c66091989c01bdb3f43e7ef31d0d17045c5cb4252d67ef68d82e07f2fa4c648936ffb9f49fa511251d992a5305892004614a03b0b127df1ba44e743da17e79fb52df07a87acd0fa13d85234ddd96a3c9ee427977c194d19360ce74f3e40e7225d8cb169987e1bceba19f5dec36b103257851ea593aaf74b036ba0584a0bb62e3dcc827ca658042c0fbbac4462f6a74054bcef63934504ed4e8ccc3165e00a09f34b9e18149364b2d01517d25ada35e78aa9ed799b891a8710f43e0c74e0b96b13a3660ba831d3030e1f2b5554c679608c77ae7975282a817b6489b5a19b7623b8afea9fee2f9fc4d9ea44838446db9e606cc0379e2705c05845c2b84fdd4cffbd2faba726d097504bb244d6c0ec2c2d448a5f89116cfa7cc9b44a5681296e70648c3c76a62d9304f64565a5008ad96be255c2529f3516f899c15c7f8dc4151d1a0aef7beed584570771d3721ed90f3e66fa4c6a6f8e1c275406043c4a6a3c1d57c341728b83f438c8774f74162027472225dc2bdfd67f3094344115124241138ced144290598c9c9bcd9075dbf7d3dbfc0b578eb6e05b3d8369b0f3944908815ea6ac570fe6da3ac5c2d6d897d73321a4095a0dc625ffb0e7b5efebf10a242ae8fa8207b09ed1e05dced71c51b3e3afe9a8031a4a979340e8ab2611e2015627cfe21319176129472659b37137e1c0119f4116b62245f3c608517e2c7e361bb576e1a07fccb3d432ccb529d4a33cf459d681981d5e6f2cd93aacc9cc4565a051b04664638e0f0920c73463edb7b684db6869f1f6aa2293bdfdd00523b4580e21a535ec77f3dd08f3abe9e2ddb999366c079cacf3128bb97c9783bb7e0b76b6dcd6a31d4a777f35e7449278626c35d9d4a4410163156588e4b2136cf192ac3e45cb35db91ec7c47eb28ee176890387ede27b6961c8215473fe04eb2d2dfd6f54329e3c63b0a8f6bc4c644894038673ce32cad5849289504ee2fa1aa1e495d330e428bcb3005ab598fe70e908b78d398b9169752ef0f601d38a20a065c62c26a0bf81372b34ba05dc2c8642c7b58dc201c238781c56c9dc2997eef8f5c5b3e07f25204eb4356e16c9b6fa93845dfa2d40c6f792e60cf0feb69a912b5a77de54dbc3e1919e6ae2d685bda87eca30b153b91a361de626b03a598d932da28e0c8c431b8411b7ad661ab0c7913664a6d2d8da7d3b03e7cface44a569440a4f38c00e8fe25f61f662f36b035de30aa655b7e6482124c194d901ca3c2244745f0f6e4fcc8853856221264f85059287bf0efacfd29c9c87cfaf945e817f324f42c9b17695acccc4e8237ca89814b5ae1d365ded47315d65921b6a3114fb398da59e723fcd4681fc69938523dc9075f864a1c9a7e09c4654f6993ac54462ba63a45f02ba44b41b07a59cf3c7cc2089c1b8c68648523afc9fd9aa615b9252809e388cb27eef77b392faf26848d3bea7623163d71e13c531c103b0bacbd938aeda52ed6649949a8c8e28587ef292b3f8fb70c04b65a2f2b85a2fe3abbcedcb27610d1189bf51983e4c0a7b2c945f9ad82c00b128d9e68da272367cbd83242df7132ef284f42db3ceca024816ba6ab96f7c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hddb5179bc00419f2cb808ff5551f90384e3fb56d8cadfb5bf354a270da44edc22b6b1c597fa81bf319173b5f2515e56beab9ecbc741c4dbdc7f52f3f8f7fe32112e398f11a65ab4e5e1edb722977d6b6b89880dbee48fee2e71ea5eed10ff915d1d7b8a162278df6dfee33537fad64f98c61b887056a809e7f87ccf5e5dd3ec580b7aa631375e8f4287d91e572337123449c13f84e1dcf5c2635b9be98ce7e19492870b75c4815057f84c065d4a2ecccdbdf42e4a9d1d4e1f0db3acb5569275a050407352cd938b36116dec66c5ec10a56426138ef210598703427ce39420e16448a151a3a9b4f1ebe8e8a4f3ce58bbaff5f18926d90ed8b3d0ef6c9a377cc29da7088672b07414430efdc8ec640380d4cd8779b6152eb8376442424603ae296ee6c1536b1c6d8ebd0fa40a8232043264f186d924869749ef4d524f7c6538c45f7f1b3cc3981026327a3ba8a8224b646a75b2421e76f37aaf56535dd8aef8cdc2828b32f77f2bc8e0bca2a03bed1c7542d73f940e027408394902c9084f4d2e53ed3ccf7f10824bb675228804efc49f58b1abaf51b2c0e7456c7238074785235b61cf359ced74a39c14725ba3ae6e352b42abdd05dc9b0dcafa0cf99b440a8282e57423a793c96e27a976bc5a7eddb0c9d53ba8362bb0d52b64716ef9258719e683a26632d09014b118098037f4b68f27134c7e9df38a875abd7e77e5131db0ed798c12799a4fcc81d03999320f65603e3b495768c12421f690c96dde7c726f850e0bd6fd64f9726e4524b29b9262dc2282b354ca0a4796406f076945ce2fec5ff481ffae6e49e06e534c894856a20396f70bac0b29357afff6329a3ce2e85f83a9d4084f423574b8c283ca7e334597e30b186a40b206283985780c2f1eb83148669c90983eb3afffc56a1c0aa409e77b0ed81f8292f95337ecb0d77054afdd23a8e65cac3342b0d8e1fd578a4b32f43a296082764d7dd32b5b66ff6862102fd4884e5925e6cab299353527d54af49067d6d367fda27fde53bffc22d966a3c12582073cb632d36247211b756e2eab2eb7460a4fbfc68a293fc2600a0942e5c9fc9250d45114229cca6e134819b2df56486930716c25c394067af02913ac35ab8b9b1a47667f170ea8dbd4af493fb9bc9724e0d0075b40dd0aadd6a0c7275555cfa15bd727055a7763bc01d73ad8fb0dc2e87a4095c5bea3ea900bf36eb342f48408eddd06b89c98db051f456d178d6f18665b60f20dcdc993be2fd8a5c6129e5164c9fe36bd5243085000820cec97406cc0146b99945c9ad522a86b56529640da9c7750a6b6e3e252d004fb9499ee010b7bfcad25b3586608d35f0ab1eafa60d2451b9f34c50c8b0bbbfc679ba97e6fbe9b25c1bac1fb67fd9c04a8ca82c5c8b2a3556a53d5a0d5cf2dd9fc6bce309c21b9b04f3a32f9788e21fac194a32a139c03ae50afd3abb677d17e2a035de495352e486f9a5f87de41b1c977a64c354b3e284e811cf58e1895a2deef7367d3a9522d5a710bfcf22804dece9c67be64058d443e28bb3aca8e538d072c8cdc0d7b9295334334666901b63f17efb01ef753e19454fed6b975a036e2b906efc8b24d5b4e047e27a688e7a47b29337424cb9c5c0263ebfb4236754ae490d95b91f3bb264e3f2eb90a331998e82eee2ddf042081aaac0a76a4a7f2ed9badb2665cad69b59bffb495bae95f96de3fee1b33fa9e123b66c4d000ee4f9cd26720201bd2a6429720ce99e923561589e0de1326e32ceca3afb5a8a9c27892f4ff99ecba11cc7904253950cd573bcb5607aeb5c3f1be634a78ba831342fcfb4a80b77079fa8cfe42042157ade149886eb0fc7a42a71641e909fbb526fafa209259cc31221ba7d1a6a87ef531e09a35558a17e781606d0226bfe4f9562b8103e5f34fdb4fea04c69c57f17183ea8f81f5027b2c0c78557c4038a87622b38e60ab12edca820cbd85fdd380592aa326d4d1a732c6c1de98440e00c15802388a1655ab5d6087d6a986b1d3488ea6ddebee3d37b8633ccf53621baa7b63eec0b4ec023091c7d07fb40547fd0a0c87d828a699334b91e68b9a6a588128bcff5b850e6eacf4a91f2e6b6cf6d131a1e0af68efd4c1f99dc5be0971f5fe6cc2d1b1ecac5b08335eb994e313d48655a4bda61e7aa649029cc25d87c80093d58b8a7a0692302b688d19debdad1031503e07bdace658810db78028488b5afb6c5c8abfd4ffd687b142eb1e106efeafbabf8203261b7c94ad8916d5c28346e5a793058fee05a74e5d06f07dcf8438be67bd33dd581559108eed9091199d2dfeff7d4a7a818417bcf37cb90acf95b0314961acafa5a7ee33595fc60643d429d18e17b7793565aed7db42505871ea6858e15a2b975430ff4b47d0e798947209271f81eebffc1870167952b9df2e85549ed61aa4e508a9d627e1148112b2727532bd50e760e8df3fb648492cc95b598a4365cba3300c869f641fd7562bac54c2b469d72bd61650bab1d90fe5d7ada53088f48e8a4f739c93b484f9fbb6884e260989990be86be28ee110ee97dcfe90b5a2193547308a0c90d0e6651f5f397dccec10ae639708864b8f7fb1181357735f084b98c323a2e5ccd93d4cfff2891906ab8a86211489e42dff3be9ed39e0e9a15fe127fd797f91981c38db0cf083a74bbf87ba2502c415f2b7a6b5c2f7863c9873db9fbca8394f023a1094948c448d2c276f05083210ac7e800b6245c72f1310045a907710d3b025a3406db324cd04bb898f83279ebbde7bfd4c84d0dab5235360b811bd4d3f2a908a906801fc08182979fb635dc69716159e5cc928cafcbc0127225add2cccc225a4057df8a6c7134c14a8d32fbf97e5f26ba252108c5eab7bc9719275f44caeee03aec04dba23f869d0679411ff5c6bca145d581dc81f3bc141db19cf8fd609d3c198d37c7b25b3529da3633e10b3d1eeec352512e1fc14908f06e8d012f8a000dfb34448793ed19f26c020fec1d57c71239a9d618141d6d6443935705376ec1266f4048c773ad933f83714a1304292c8494970e7975fba895954941b15cbb409d0b0f85489480e0b16e3bb9206920d1691a8c5a8556371e8099a9a3efa8fd24df8745973260e5373f90224ab1821f531672f9f1bbf170f3e9839dae5c6f4bb4e7754ec4208544045de6e4882828fc01588805cdd6fbaf74445e724371be2a92e5ef2619f81167dd05d2e9ae42818116392fc85a90cdcbb5ac83e8d90943d59cd1f76c7eba2fa89ca365fe056f6310babdcd2e2f3bca41104fe786560663930baad47b8a006ef7b2e0333e7a4697fd80e4a43eaef1063f0d5fde993381d2b9095a16a254844af5dd4c7cdc8b011468c71b0252e9388d9df8ee13257b4d1c8ac33d5745d73852e9dec38a7de00cb6211e1455d420683cfcf5af83572ababf93db2c593008ac866f6041bfe65d151deeecbf0666a1c7c03c65ca90c487ec9120e814b4c228608b89f733bc36966a37a457c96ea04f2f5f19f2455b94eb2bb3ad4fd45b442b8e86e682e7b1bfb816e2d799992bf56ebd8d6403a8e6efe53cf56b1d24f18f2a9f334f9fa8a23009f36a128478968e9c5878ff672700f2b90dc60e65ac213a2f7e30f12e085fd15579dc57859df249f90214a999b74cddc54fae15a252575b53e009b7e6737dc9ed2d271c7daa2be0206f11ddfab457acf2a22b5364773eb34ec9e566dc7d41de1a1ff847eaceb305c9f6f4449de8d42dd701fa8aa5f53b50628ba35fb7eaa78d12e2b1c4dc30a8bea6b7addadced0cb5006d767c9c7a42671dd2981d4c02eac4ae64249b87822046223101459057405f60012cd8e036ee5ac6d84528bac41af49f13264ed9e662c99e56cba02b26406846dec708bf58ba2344562e1a30eb1e176ecd91bb905ff628ba8c5411ac6df9bc68234809a1a3b4db9b7da4578549c9b8e0dd57bef92191a6622194fd50095359f4389cecc6815215a384b805edb49c0178817eef7bad8df9de08f2c6756fb311bba89fbe561a87d2d70911d674a7c3469f858c024932dc78da9ad95f5cbb6038c03a56e3d4cafc2bbb36119a42d754ef42b69d5b64d842d914ad5c91558ef7302d1919d7c72bb3090cc4686730978456a8cb53be64fee9b953e78f662c9a52d009cf2a9386190fa374ec2f11afeed87ed926f174ee0cecb2992f253a80cb87c4118a20c7a4aea35ab60acc6a604228e6c8b2e4775ce873ae561787d8dca3a285707997c8004366062d9d71eb9dee4735955941281552774d9bead4467420a01c48b88a6a2b97bccc7388d4cfa50aed563de4413a01bb6bd1c69949d34a8f047981ffd875083fd6873e4728d4f15948aafafc6e94fc473650d7bec1d5c12e7778a5d53e091836245950789177f018f711439c711ecf2306ce5f84ad1bc9413a6144b530918527629732352b4392e210b5e3fe41f50a5c41384f74b64b7a16c5299a625ecba79cf1e926ed49bc632dbe683c1d68aa4ce3732052c1b7415844b2c857219c930df79b0d17cf8df4d95009029fac08360d19c01bc9e53715294b6119c762f19f27a7e52bd00f19bf78031de0e91bcda0b998750cd9d452eae1c63b7d3e8149e407583f610354d260ee74645f60572aae41bf10225e7fa4493262670f9e39608c29af94c2f01f2abf3516ed1c95a4806db5eef815b79ecc06d0f2e9c54d2bc00f96655e7dc04224f257915149bda774f468da425b7ebdddd6a5e82017f457546d6b0717ad91f98f027ec2effbaf1b3071ce7ecbd041063a2b3292cefa4b6ad29d0666828892b35a33b24a97927169cef19f28c169c4dca582bec65d3bb7eb2209f186ead7d8e482607c309de877499e7751d269d5ad37006afc93df88b805d178336ea2043b2fa66242bfc65b4b492af5cf5d782314b4fb5063e441a3897b189e9739d11e7e443911a1bce1cb685fd62a0e986cc2ff8a7fefb36d55dda319db2fb1295039891cfe115e314c0cc908b155912875223391845c883e74040cb07491622e9ad0d805a5d1eb4b80754758b02008d1202900e55eede2c13c70cf0c5627596688bd1718cf208ab705729cf232a77bba2deda42171728185179e13c7607f82e8dbfbf7cf255a0f37e7edbe71db6e98a353fccc5290a16f914f19017094e873f2d33806740eea630201109a7c64bf2ca4ee47f8670c79412ebfc27e05898fb2d1560fb4cfb53dae66d7aa63055944bfe49cc4575a2083ac32f2c73dbf4805822a9a9e8621736c4ce15b585fc153aa91e7af6e0c2507c947f1800a67678b9d1cc04464bf73613fd8710098ae97cc916b799042cbc7655f3d15bb6aa90e5074dde5ab143f7473e04c3400894065872e47fa054a5250587de932b45aedcf8c6ed5a978dd2dc2207266564b297246992e205c2481663cca7cb092a998e5db9eca0d38c3d02f279fc4399719b2acb2fb072d6e6e839c335be146b85c10a540ad2c9d5e5a0474ad57690fd5752b925597481a798e1c313da035cf71696c5d2ab20816a5463f8b5658032073c5f6b7bb0aca356e00e5cf46cfa129a9dead9bc2cbdf1b363f4956bea90a935e4eb2854a455ad75ba5bdf59e81231cea889c935386acfdaf8c3b343b2ffbccd14dd38ca7e37b2aab00ab5c0b195c8c06fb835ef9a2ef493caafc4bf7c0075109f3227ca7127350c1697beb46cd5ac7b1fb2294fabd9afb9ac90cb4dc378bde3ba9f0e0fd550a6b1cc233b8e5bd9dafeec7afd0b163b09f0e5de5edee8e11d54a6600eb1f0995acc297942a9cc28ea7e29bb4fc9390d4ed9c30a7967b8fcc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h166f55f8c95e0bc457e0aa0f28c3e60e9238e9bbd23bfd76a1ae4043a7a44d1e17c377627c855d9a7ed4cb6f5a7026bd057ddf576cc86482df7e407bc34bfec531468ff77ec3b23ef9615a62e59ee4f6f782d690ee58ce24f39b4ac7804f8b8058c4039a2fb5c019ba383e61975fda6269de11c51a7fd8ad5484781e7f7c70066381a5317109be66599588eee3b4d194a3099eba7c2c6015dd98a903539b281c0c3e6aab0581830d70a35b2ac92f148b09ddb9c12db76224387ed060df348075e2e06d487ecac3c848e020a396cf8f5c38c9179075840d9cb6db637cd19c759d8cfed007d62a77e3bd491f02feca40e1951e05fb0ec85ff235810ec3841bc4e2aafa953dcf5dd3c6363265e21cf3642a8a568d2a279422237be46e0c97e1bd77bdc4cab98435a881b588be7439039e339328807c6499d855d423943b6b29dbc6fbd5e86d3f19b54eb179ebe0c5ca28ada1647c7f744ebe256c4efb6c6ee2d44e85e3088d3dd8c4f5a5ea926467c57c7ef8a01fd76d50004f0c90dee5dcc02a9b3158887ee73f2981d633dea0a9b92b437d30472a5b8a07a64c54bcea019edc12730d2bb298b667d74ceb6acb0634738c79ec3af9d9097f358431626b6e2c19379aeecd714f72117a36f08a11e36745d6d81fbd685c5e2912581e0a8f1ae58e4b3d94617f77944556c2980d54c218a77c543eb332a165d0adaa21b6b4ed83324bf4a8a5bf002b22558348b094386dadbd5b9e8154a85519bb5b03edb8036efa3ff9ea00523402171edb80f96b26ce85ea17fc8e15827f2cd696b2dcdf33b8cd9622825cc95bf93d57c92195cb13e88c2afa7481ac048f19de2601d08ea0f1043fb56cebc9df2a8a8292ab24016441cffbba732060827774bb7b8de7ba036cbbaa634c854d3bc534bbd3ebc38398d8516a16a07bafed6becdeaf1ee87932b6806853a4ca3a69eb07d7d2aee67df6dc38ed8405f6ca0f6c85d5fa96cddfb0036f2b4eb3bd64ea887c73d84883a3785eb75be5cc28c8204c913cd09d4a519911685c88b2766cb877666aa34df759953f3d9df106f05aba480c487991d2798f78fcab0b5e636e9a34455f45cb868b075888bb817a4a2eef4c3800f75d10470ec7904ca911eebbb015d80c754adee6d185cecd147001722ff95a38f24f3451d1aa7ca563fc0aceeed92dd7f333e658dff06a6900f4e7c8af123232071783a7ddd62e8e94d786c0f3c04436677d13c47c9b7d331542bb974c829972b4444d9ef209ce22f21e0deed53973e4c2d9c84a40fe9c7e9e142e30c8c66c23e5bb89c30a99582155ae1dbaf9b8a7eceb91a15007bca932d1d696393be5de55f73a12ab43cb2993c373b41dee3d7234339c021be06e45a0caf829e115b4c605bdab0ae1470271597c7081350258ba8b58d03b1ec9d1bbcac8fd53cf59366e4dd09e13896040a159528d355414c1ad4600ad19d85f784ee147ceff222066358858b3cf28767d0addaf015835806bdd82d8aaa438812b56faba7bec3c3858d10a21dd7c0330fdd04c395e3facfba6b3bb40e79aa8e0240e15c49a9c8914cfd1ebfcd8da5831a892c7497c400b391d1621655c6d48d531d9fc9c540883fe5b04c2f62dee636b94ddca225b87e499749034d31223cf58df6fa32f0b38ce375af62fbfc3e474cbd2d3e22cab7fde25a6c3cf6537766ad1d8a452dfe768e49566f5a27c10e03d3f341c8b8d62c6312846d6d21c52ef61fcd2c9f639d9d75dcb4d9939d4e8133c15815998ac9156bc6056ae7b537a4f9776f827e78ca636081572b3e5217c6ae88bd0f4ee87faeca91d86f1704e02ffad626a203192cda46175a377ca4d0f462006182de16116f426ecc214927423a3d7d88c125e449a6d6d71804659d43196f6908ab46205183f24bc300e67e60291489c2ac25c4c9729da3d7df17049dd01fa94bcfae152a47f074d8114661f1c4b25452b6e70dcaa413aa75811abc52b642d422c38fba689cffb1e7d34c1ada065e303ffc1eba144baa95c423083bbbdebb7938c6573ff3707c95faa6d2263b9d17b794053809ca8dedfd29c05d433760d5ecbaf059daa514e186728604c3dda68a3147bad51c4f2ba8e0550481afc9df0391614d7cc62b886bb15d81eb6c46717d27935d8b699603e2e4fa3f7199d24ce15a031b2b93e467d3f6dff9e02e3e1720d8f15d57cfa22a1d5d17264a8c7f4df03dcad68aae6785c1a21cfecb18f56fa6578b8b0e9019f430bfed05f0d6a405e12e3b21b6756d3a9beb4f6b1276ccac67956b6e373e5163a17c386894a538fc8a2f01c19267b548e4ba7b6aa5b6ae2e694bc9db7549e382c07071b09eff86ace38818308c26b86d4db5397b84c06017b82493f016bbf3a018f78c43635e03f3fcbbcdb22d9f5b5b0eeed36e9e24834269fd790cc29afc5bfb47262a1212abdca3aa63cb49e637c84f1b865897bca941ea4fb664066b6f49d294be80b050d39f3c6324eb33557ca498dd64fd8991f924979e1eab7f91630f28bbd947ec2800829910a698b9176a84e22ac45b8b128875ffc575d8827aee5e573cd9d1dd1295c8eea8791bce4643a6edac362123c622565b5ebe73df60f4b6e66a5392594d9380e777d912276a84961f32b67fbbfd699bec470879f968c025551e5bd1f0a75a423f1c1d89cb31f4d161ae43da30640b29c63b44563c96e8fc218da6e1c6fe21663fd6758280a2cbe3e2c0e4405c4ff81c19086909f5834cdf3a52572e48c842d93798226d4be933a2393056b50ab5a108838c932a55b903b4dcfe1cb89181e84ad1c8f0c19387355c1fa04bc7efd4b1043f95b49a6b17a7930824a90c001c4394b7fd4027123ee9834058c7b5d31509c5114badf2faf4cab25195e2ed56e5ea7ee5330021069a351e0b6079d097ea942e2ded27f5ef643d7111004d3e7abe28916b09251e427f187ddddc80f25437854a362134ff3b62859e641f1b230530a176bbbd0a30e03582617e4e699af05941b56111ffe1ead67505116619133b7ca4b4354599dab48048c983f6ca928f8d19abe5cab899e12e457ba80afe5c202902e883bb2a156fbd6c04b1f7423206899c977c180553d510f8521ffbb291d39defca01adacc3bde6ac4565cf0641f66ba6840a41b738f3a2e6e88a0a2d210e5a9536bd782f2a2ddb087c0425eb1564924c8fc67c5bf0f9077d3cf463c5d169b6faf14d6460f98ddc931795d1c9f0d1498202c950e0557d9535be7131875e07d1da6b057e0c61cb6822a483f99140bb17b36a05b07f12c788f490881d763cdd37c2bed44bd05e74b54b5629c508cca0cafa541ffe3f91bf55360fbe2ba6409c6d9d6b558925c296b7d44005e6ccbed1f9c24d015a55caf428af7762cc358c919e62288d92c74217f0c1d9bab1b48a23a5efc42c89007fbed34df8382992ab95de6c496c07a12a7cbc3cb37ee9a541dc917ec16ff4db7c01d486773f9ff2f3ab02f2697be34707dc4392475db0db49df2aaabffd1404b4387c543f64673d0bc3a9c3de8ea1bc2ffa79d11061bbafd8c7587668b7ee3f2c60ac04078d045e43bbf689d27a1f8314192f8e2ef440a831b5fec272613ebd51da622706cec3c9b8b8aed86b2a4fca95a91db930a46d72a4afc02e2891ecd8d4d3001eeccccc428f2e03ea73bdbd1ef9d5160a14c206fb2a132db4d1d648e345ee987b6fcf5eff41b7c6d2fbe8d9bc905afe6bdb256f9c962468115daac27d77181a467385d38add343535ba10683d96d4cde3afd91a75e60f8a1b43d84f203d1985f27773f5d6c1880e01eebd443b43fb4ce5081bf540e7996754de042d009b11cfbcbf132413376077b2414824896a5b41d46a7af022416819b35443af45482206182ef960dd1a2e014ad8bf58acd3d9d1c7138a7bba479552b03c9e42390bc3704688dffc37797fa1932220f0cf763f60fd6dcc4efb7b6a5a45cbd02a41db6e7599c44d201ae0b8babbde28f028779878685a675fcabd4109e5b62b60933aa62eb024e8fca536c2468ab0854177a8a8611fb1b3aeef603722c3a3dff76a2f0f0654dfdcb42fbf48c5610179b39c37476b94ef4f926c8e3bdf6c1bc3f2c5301058c6819c60716bb6ca5f3253b46f95c34225b21e731aa837b3885d6d70f0ccbd5cbc64d5a71c9b379b07d08766f909e5dde369ebe672868ce18e53a2e82d2a8770c99e063d1d7ea7a0ae79a18c63e334eddda4930401a10188d5cdcffe25a8e9ebfb75825619f2422e9e5762a5d3ea5ccdc8a16fe24065439ccda04ca49547e816b7dc419cab4e2de34f9f94e799f6284500cdb474a511764cccc91946d8ffada50fc84b54be562131e9a006edbd5ec3874f9c608175b914c1a47209fde4ff670a9d0acb70dad4c760b20df58d92edf99adbf5b13937bb6eb6acb35cfeceab93a1bada0e818c0def93c9c0f3cb61058caedce81cf243c2c066dbce938509fb6b925176d459eca114aabb312154808e2abe29ba7b687a4cda557932dc6d2acffb920a91fb09203f9d20e303cde0a18a02b38fa8638bc962d11aead2ba2782d8ead38074f701b845e727e874b488ad909d028907759fdccd0261bcb2712e604aa61eb1e6095383c7f675015ad6a35c992da69ca9254e1505dbdefb06c2c51a8c05430a74089e83d7ff0454db48dc3c31b06159c8dffd21f220f887b8cfebf17e63bfaf42e7e7261e359d9e156765ea927a515185abf9b394b99e89c9a8f30510c20d39fd5678c7ff65d993989914abb5b51cd820ef142ce1fcb17b333f3edc9fff9a9ac20cc485a3cda51f5a306ed3f7b7d554e068083c3c6e5b5afa7012678726692cab53e143fe89d563502693ac8cb8f55c1cf9d8e5b67cb6b49db9be2723f335585ea7aeaca6626f107dbc6e0ae44c714f3f3fba1ee6049e0161d43672becfe8433a54ee2fca6a8681711a925fbd99c358c682fe066eda5a17a2cc1405698ccac715188b60a15f5fe0a08f0d216e201beab01f8bffe072b77a061e0f4c2eafc9c949abd156165b23a95e7d826012244f069cd29d9196ba5cc2061809ba46c48703fc8fb0480b46c7f662cd72b6391e88f812ffd0f09e0b92be27b2245fa29f486316cfb1c609389b3c062df5e0af99b238885c9a778dd3922d10b33c5022d3f2337dc203556292585df7ca72f0439654e8897a9d4b34604a1fa05f3e1fc87125e6ae291959d5c6e1f3f3d9fdb1920653c1a33e4aed19697ade1c34c91fedc13ab24f977597c5fea39fe1f5cde3417e860e9b13831224a176cd076ae4c5bb80def57cfaba931b2f7fa21518d888abbe118f816c8271dde2291d282345c8fd8d40a2780a5308f839ea5ab0f387b3a4e7afe2a7f87be5d4aaad0176019968905dcf0d3d8b943aee4d3302c51b9db7efc540f1620656fa99cf627d4380931abda3e16c25017fc4803be82c71809a4d2310e8e9cfe8721cf2afb27b536ba27362c9cdfa36794556dff3464af600c6d93f51a04b4c8b8e0068c169a0bb60b670aafec18b86fbe0a9ce0812333c700ec3df5347253c61cac44a5026a862694ccd074d087aca3af2a47ac6c9c97913ac2f5eeb04034aafafbc1296441e5f402c91153d759d8328ee9117f99a7bea0281150bb7519efac4660b85d09784b55bc377d9efe6ec95a760f6f4524329b385bc805ab619f8bfc084300d86bf17b0659a6eeb15b988aeb6a1eb1a3acec9c7a56af2ad1e44989c2d97a316883aebf57201841d81ad9ce02bf4ed771642f03e43437d2f057a5dfdd4d4a95f94acd38d38b6c55d4632f67090626f4ee3e4142499aaba93401;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha93403d0bc707f37554d4020700e930c3b6fe74b6554a34b9a6a334398364e23c824cd088bd99e7573bbf74f3de5fc6d85c001818346f7980b7ad580f0fccd8085ed220eb74db3e094c21f2c1aa5568f307a5d933ddfa0e3b692248731d49d7ac8dda9812e870b7b7e094d964f47ece67a6dcfcfecbe856abb03e4e35f0cb48156e2758be1d3b1eef49d276f43efcc6b1c27b7ac9b37a20ecf123e94bf3cd04a807917af5f35bc811fa5680991521e0b287ad6e115bbc14780e4202e033c51d899f74de6b3fbc796a0b4df223a92deb79f9872fcf293001261204c13affe28b35ea123e821781f7ccd0d6e89a58bd494c447ac32a3c492c27e5511170df7fccfbab691883da1858f8ae6baa188996932aa4131ed82dd7dee54573299459779a300c7c403072b091ecc09cd0a67921ab8ad3523c971195c95d3e8702fc7ed0d007f42d0827da40f7bed9e6b98a88d99bd7296dedc93e356ef384541a6a314fbe7a940a177ad4f3bf88705570782de4869b02059a123b1f0b18f9edeb56aef68abf9324ba8393970fae6c3f868cfccf16eef8861aedbb66bc34db78663d55c8c7e0643f7e363a4f478786738228f7349106c4f81d660c31a1163c4cb80e893fffe43e92c303cb811ba8b171d057f4905fc7ad70b44e2548a51fd8f39d51c0bbfac898f6d193b448ada53ad7b8b13c8b274c166aa2431bbdf4874896f38c0683b973107df7f7c41027d12b92509197f08e84ae3ac1327e40b277239e7777211f65ae941586fe4e5c70680730d5d4c079fa7d4a920f87e2d615bf7b29ce031252ba3d0060661a34d0bd015614433423c3e605dfe9cfb9911a90805c5ce26be6fa011c301030ab6defd63f62a829772a318c019889d813055404f0a610f74257b781f92722062f73fd814b045e0c697b6c6b528bee05d1a3bcd489f15c265f4ccc41220b4b49d08fe477a6182b2a00c8b43c04381973dbc89a25cb125f0bf644e7e8c2421983758cba9036e7f662a398fd83bdac6eb06874b5a492c47d74b7f28e98f3093db8df84bd516916db07fce70bbf897ed8e121dfe1abc8e77edc205ae1b2790a1a0a998db028564dd457b5a66951aff0319d995b58cc6ce591e5eaa68d3bb617578f33b78db7029959a801e588c54946847a8994ac97fe4bc4bca56358901d532d0a3bae48c2c7e5120c1e42b77bebc949fcfc671b1e059c530d164b1bdbe5f3724dc570b6d922fcbeb0263cd1b7e24816981612ae62a7a7c368a7168a175776a69bd186e9a3a48110291574748364f6dab5c483b33a70ab144c9fd226a36fb1ce2fbd997a9e9fcfd9aaf3ad26da4dfe04f639757f3f0eebd6dccd92a7cfe72296f19383859fb3d730a760958e4a8e7ffebdeca1822b66ca02b458c74298366e1fff500e816af34a2b7647aa946a71bc3e918d8f09e120d3cdd58ed54a04706274e10fc3f713e21e7ff14d1b2220cc55f173187a8b144a4d6ee1b3aa42b466440bbf3b929ca881e36948d955dd850e466f4a2b95b31b5d14f5fd77b64e15025fc8273797b8ee7d19290e151cf0f73bc9978acfe5a948a01e30c239b35d09f1da25a6fc7ef43fa0ed80eb5dfbc2f303f117f4c65ddfba185cba9bef891d7cc2744626df9a265e97c210c790939de3c5eeecc1f1367295aaa88d27e2c2adcf29c5ffb887998cec960c12fb3839cc76ef0a1049a868e1df80b5e8ad27966882c7a803d275cecea80a9e64381e5a78e812523de0a494653a1ba3114fe28cbddfbb12ff588b6caf57ca29e41ab4119548fef9ef4b930e4905af7c9c39ae9e44f00209974516c5c76b8df2a84e8f8e8fa19a2da39f04774e22bf9502644189c51a5ddf2af7a18eabdf776ba0a13eea83a0cd56c391331f4dad636ac1ee6401e1dd5ef3b46bb5a2e19296a99abf916824a9d1c696dcfc59ff399a32bd4b156282879c21c3ff8a44757d49526995ced43ad3e31c145be8dc73bfad52cea3bc2e9bc527437d84da2bc02f9edd7a89a5aaa4a1c3b675b3aac64e91cab7939e62abd6fc0e9a12b10eb9de7b004690394555a6d83b1d76a3ec4a595fac7edfde16b1a57b079f41e7fcb2ff9055e492b2f61c2c2e8fee9bb6547a368ce3ec73a5102ba99489e30e5104f2d2cc0bfb6f52b6c7d9e9b7079aa661cc019a2b135f2d883a5a76d4c59f6636d90a13c0997ac3f1eeb1084abde47d169965ed752eb512276f8ca578e7a5ce4ad4c2e0f7baac405a15a13655a324bea17a62449ad0b6314a1d62935137813e9fc96385d6cd5256740053fcb4502a50732dcaa47a3ea9fbcdf27cdbdf449a629adc11e4859f75b32412129393f1ce14c305dd039d514aa99a12e1719c1b8c74827d99f8f8c0f53ea90cd91a5f90c8401a4a71a0662a1ed445bc4e8eef000fffc4fdfc6b2669bc3e4946064b6bac63dfe19889998c1613a5a1cf9cb197c4a5c88d53616232536308e03dc448fa6bfda355e740de0f40192ac96b14118d136f234a312fecd9e36ad326dd3f61130ae79cccdd4ab2da26e3412db72e9a1a7f0f67db33806503ec07c8d25d625807af300fbffb3fed3238a655d6875b6a7f3a9371b5799a39766833ae5a8e1498d59cf4f688809e834fb957878138333348daa693fa250f6c4881762f51e6f2941e1cc0e107a179d073c2e4043ad926078a63f4064b0304df5f6841cebe6121025d1f1e6569ed99dcc412ffadaa82aaa56614492ad7b98393396708287aa83aadba0d83f36beb9f46a8f304d28f4ca068cf9a7efd3a0c938f6ddcd6f175af244812481e347bd88ff343e8870c0d60d878e7e0a4962e2c4428f7f31e585c7925f3856e4f94b83be333e7e84030c178089472d7f296ab999146a7c9f05cd42952946da777a7b12224a4c435adfcc0659e2161bdbb6afbbba4e23bdeaa1a12c433e59b212ee30cc9b99161bc7aeace9b185d27510565cd2a31c2b6f2d51379a8d023e6d0743aa47456327005f71470472657041d29bb219ef5cb5855db2ec28f3d4f4c9c9a98425f51897de9e0ea6d5c6aa20e02825d70b11c2ac91802b99cd8d9f689318959542c24e16e18fb48939adbb09cbae3517127c033792926f9b8df622f19ec57526bd4a7a506e235720b8a322c008f5882f604946749a1842a8b6651b55b29fed0e1e8dad9317654f8163bac50d1d3be7c691aa276c68d3cbea64ee444819111d250a50c64058291acf9fed759d961aabc0e6539c5e74c902bd605be37ca1f33cc876578b3f6580f40595ebb603430cb3bdf85ac6c09cf3e3e93bf089ca915193f2b793ebe8d3f7ecd662e659bcb5b9c86186c1bab85e6358cf66b5067495f23047c9f7089573d988c5ed0f58f5612ad4eb728319742234083a6fbf1f81687f9f81204ca4391cb17647f3a2d6571bf69d8d08e90f78f2fb57505a7ac60beb39b6535c8f847861b57bf6b7166ebf56184aa60bf8c9df0757fe02293045dff3761ff1cf42beac8d85576fb5ca9cfc40dbe4d626da660f1c34d3afcef348bb91df6718ce984e9d80092fabe46bc8fd0d577a8c45d62240d721cd9d7446ed5f3de6e13d6c7bdeb40f3a41a13f79a67d2b8cf9c033fcf7764fa0c9155fd361ec24e59a8ded4b1185044c9a2ab591ed72a4d5c083937f3b1522136080a1296e7f94a0ef1b39e2839543f9e66b6167a4aee3ffd49b7b6ab33c078663200ad7b72a04b8590429c873450fbb632255b14958ab718da50c69f4d612dbea587f5d7f43736d1388aa056b2446f0c9b643bc5411d6008b6e9a0e45041e039c252b4e3e3f294a35998dc6cb3efa6b47beab69b37e49a3892dccfd7b0a43fbe06e2c37059dfd25ae384be4044da9719ed12890481afca85aff6d3e1e6451bac49b44e1d03cb2cf84adf168155c400b8a842bfc1f5132eb0e2f810e3366b51f82d709539adf7c47de1c2d7946993228738126ff165bf6663f55796a2aef1ba2aa49972369ab3c52993d8f8058ae0ec02a3765f4520934bcb09c3a6ea7854582892ac349c8a12ff98cd742d7c7c6b67b7343bef95a621090a9ddca94a5fc94ced94c7d6fad69adbc6aa9f71965bd453ec2b998f065a15b175832d7407b8c57f5a9e7a7d59bfba89188f520ab753e255ea7edca84ef99c79aca476ab0089f600eea80a0d2f60989948c4c4413fb2316478e8830d3fbc992b16ebc088ca1cdd02129a2db9c6462752b5d3ce4c559c43c275eed793edff59e9ffd2da5c9ceb7e6fa18d3986d79a33eb922f015819e6a43ca21a494b4d12eede54376933e2298f7316ec1ba5a3a0de298bd6b5c22f054e0d1b8942e38d45a1cf264466818f8b0ffc8068a009172fe59335a7ab95839d227ed8f46abb5039cf7c6c95ad9288fd0ad6896c58bca64364b165965851afa6c9a5da79de1d31e69c281366ad6dc1eba95168aaccc2b8b56b150b619b4c7f2d822a44e0d4ac596a3361f657dfcc0ad68ef9fb66705910241f91c8cad2f8f329ad905d84fac4b2714541a86c16efe0eed27a7cb13439067cd222ff598edde65788e1dba0ef2ad304115c0619cecd74c3e1053bfbaa19347f18435404d22d8dbe0f57622db0fea65d80883612dcf7ea94aea80add07f1d0db1106db050c21ea2cb3e0598d8759d8f5a782b526965a547bc2d740c83718daeee21c80f5d93f1dce6db549313c5bd107ca5a9c5298817c4a9d5c495e236d7411ee750302850cabc2406ed80a42a88391e62df523b4f85122388de9b956a51e82869ed74e3e8f4917c36119b4cdf8dfb8a6f6b50a73de535bbb652139c2acfad0b075423171df16af89a47a834d43a16ab61ce1dac1eec6dfcfe1164a6bca8bed1f90832738021d020efa86c1d3cb41aad29d0f749aade57fbad910a6dd6fb03b22608227153aed49e296a5e53a0e338b9763d2f314281b5f08138a231c747ba2acaa09a9fe3300be4bbc0a958ce4827d800b9b2d17ca42dc42361f5e02a4106eb34fdf9889c7b161b8417b304181f7bc3c20e33601ea314e9c1244141b262cfa953b9e55474c23bf7f09faf22841b1aba15d4393fe0c98f8d92dca2ef30e04154488760341ffffd984719b9552ab9110e077351591a2d382355b9502783585c1e6570c19c2902b56f8b9a2004530a3d0aae3156d092c1832d8509cf49e2cd16224365ddd4b3b41e7d40406d760d2dacb2c9a1b102bfd59c7778065dde6094ca90e0a38d0daa2e3226175b3f5f9830b79a02c83329a98c5108bef8381f15fc66c3b811583e1dade97c187cc78352fa46b2c75557dd8ca3a29e714c0b13090801e5aa043b5a5dd89ad04d97938401cb407045efb8529d82e2b582bf13e91bfda91569ec55d730ec5c294f8a2d6e486492efdabd13cce652b646a9fe53fb6aa88bf6cac5426a3a83935fd9d39a3f35459a4447ca853acb2023409b2328a65a639ece8ddf8f229325ac4c6a93aa3d39984c6a920f2d165b9f95635cbd0bcc36ba4fc8e60218f09c87c650ec1964edb16b55f16bc83f91cafb3fd3ef68464ddd87b10f82d0454dbfdac23b78f837c5996bb3241e9fccc6210ec0851d331776ebb392331537224af5867e9343c07c011c5b58c657348e87824e325f038658bf39ff5f96697cb83a2383517c3098d6250f690011c0139fb7e2990a88545531723da2b3a81c7ef221958995357b4891d1f8eff03a1dac91d549fe98c47a8c2a8eb0f9c4bb54b224480879fa65f6561eb28ce194f4276a28a0ab984eaa00bcf64fe431285c4ee9211e8d92d6261aa1a82d4acae3c9b15770a1a0a6d4131a3b9628d1476cd2ea89104383ff562ab6b82d16aa727efc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5178434b1220ab3a9c50a2464a07a4e0c81c8089d3d237032d01ff0a3e7b9129956146e51719e09f404c5a64d67060c5379bf429a9019d9cdc4512cddbe310f4436b68158afb0002a82ace7df530e4fcd4a067ae8f348818ccf1d6a270acd21f3e6b710379a64def2337c4fd6cfb2786e537e57045e4a4e84d78760f07119ac817bcf28c677188f5fee627c184555a70087db25a5709775d2057c4e587d3f0ca4dda0a90943bfeb1a5202b6cc54b00abaebb2559972f6527dd7dd8276d963dc484cae7f6c650d56bd90a634b1ea4eae35e4fb928432e1dc6034db524eab716a7fa47149b36e3969873e81087dd2c49074564542088ab14d6f18481f3e274962afd9a43a34ade7bd79f7d6a391693019fc83525e4d2e5a9eeebf9b2f2674e1b9ca0de9344a6dbeb25bdea4ef5403e2cf2359cda103fa481e550b718595dd8515388d97b9fb0b8f55886ef0b4495444c7f15a0e30f04581c6ef071b70b0913e48b737d2ba293278e87f6b5519b44b55b80d3aac1d162e2d9e5fca3e41f1befacca2488ce94547108e8053254fdace3525b0ec1590407bf91b1f69d1fbbf11bca28fb57bb50f17bc2962812185da46627bbbba8a3ae249bec1d170900ec309468abd8e0e89f2adf56db3611ed9e127062b3cf6bf97b7e8c277ccd446e25b6db890a820e55908b8dca297687690991ff4cff110971c7335493831c39d910a704ebb1ccfac40939d54ca504900282c4295f48ae3b5e65543bff0a82a11a7a5ebdd09a2fc2f8a39c708789d658bd0e78053927671540f4cdc46f15bd3b3cf0f0337c5d03cc7953c6a910139579f8ed94a749d6b2dd2c86a9c9bd7efa56ef4b7ebf8df4f23d63f1a296dbaa02025f766ede9cc3dacbd2ded4f8283082ff254ff2c106ef8bf7384df08f0dff0d164c7d6e6a1ea617ed04edde2aa578a6888ab57dada8e61bb1a09033a7166c9cb1f4213161321db7917ed20f8c97262db74a12002d1c50a1f135118a1de130ca0c3a4769eed1808f5054752ad7de8febb631e2c6498dd937532e52d4bd9e1671d04f8dc3bd3c4bbb2acc424e460a7ff955c4e0f042ce6ce1602cd19ef2b6ab3d2e802b6fad821d9f4ea3605f69ea0df5a4dacc2367d01cd8865d2318aec724302d543e604095b1886a0e71c1088280203a0293a5fd4708e6691a1f9c5460fffd53a8f80ebdd31eb3991ac22a8fb0a8b1397b620516c8a4f2a63334062ba02528b4b297c0c63f85ee03ea07a32b3e7e690359e66a78ab6ab429e60674357857d6b2b77d1fcb2c5687b1e6e3868e517c08c3f0d3c1123d3a3f47b5f0790b34d6180c924d45e652ae3a8b64274db87a92c824dacb50d0f24816336fee69bfe518e4c337a161ccf55ea1f5ffac47ee8a76cb97b76960387e74aacb85eee7d304aeb65688841bf49a94b4e986942ed2e2bfb92e7851badb73ad04bcf597af4e1b37dbdd87f442cf6afc43df2365b26f0593d3b11d603437df9302476891759cd01cd0a2a08facec8745c16ad9dc3951781b64eda5500851567c57ce00d9b50fb66e46039426a5231b2ea419222dd0a67e1e32d16e5ed810543d7396197c439b15aa75a742ee74a0886af5040084b9108fef442eafbed836c8ec412986c9105df95032120ccbe6d05303f22c080498555ec492cbcf6e6c38c6fe3be98a51f694d37b612c20255acc0895382c14119748913c574506e35d0bdcdfce6ad6b05bf32aa0dcef7556c8345d5b19b70b2f3f951e3111f2092a5295f903fcc7b6762ed20b7423ad1e7ea46d2cc0e8a32925b3f4a54126f47bba54efb87726ba755849aa76497c577cf8d38ef25093acd1c983fa3dfcb414fa3426fe2c44c6241fd14679ea4e4cf0b6a08dfff8fb272596310aaef80b42427c603b9c62c574373ff555ab7dbd37546359178dea1cfe7b3d0eeedd22373f426fcadf9a4a0f72a3647ab7871cef206fa2be919297f799c741c82e7328fd0a98230cc89b6f09e7380986663be44554858614b1eb948b277e6ea2b1d45118fa39079ed572c9f2fa743aeea97deb7c73ce4c60ec27d7c8497e834ae6e07f08c5f70658c6eb4cd9cfcc25f3594a54bab377e87fb0af75761f3153f78525c6e37cf828a77bd5d68781cd122dd507483875f421df2bfd2829e74a5a235239cc2c759965bf501def5ddeeba05478e69ecdfb0de9620ef4bedd3becb03d755eefef8ea8a00291e769b39c2d4ffc2526f3474dec87138fca1c276fa36cf54b86b154178e142a3346555c8c0fb5ceb63f2fdc4eda93ded2f53b89a67db6a0cc99d2584df81ae9a2ce100a4c5e94156a70f3bf264b8885b052baaf11c9a5ee011a094cf40e82954da2ebe743876afe583d95d9f919d0a678435f4b96a1084659e06fbbe42374b1cf67231e2c00479cea505b13ecf1b7d607e9dc53aabeb47cfd20062ca2513184e9e8984b95417637e3a43777005a774b4f8af4d4f369e494bc0f8e6397caf7b79abf1eb82eca22ecdc29d65ebe9f14dce5a7ad09ba0daa37ebf9ab626e470fc0b40d8ddf5769488725d3734d03f1c815919b67c83243f58f5d19a20ce60fdea318802e1af39a1872e1420641a9327047f4316db708c1e12379d32ec21db0ad9bd8a34d650aaf1e830401effb65fb531b4520cdf082e3900da718c78518960b431c047fa849e633ea0a3910b39b4336c29b4cd7a83976517c7da0b0bdcbe34a6db3a428b0021bd7f5a33d398def252fdcf33ae961c738c3bc94d09e26b1d1e555177f2153d40d9cf69de9563d8a84d60163f50699fce0e319e3deeffddf9d848798d982ef2372c2a3b3353a01dd22da6b36c8a99e578edf1eebe8795c1cc5462d27f52d0743613b13293344c50c96053d87c990b745e6f707d0724359f0eceabff00928b942052368da671fb44cf5cae424d3a64c9854c47482e449c867979f950afbd2092550ea8131cade0bbbc5753cd900370fff7f582bffb444e65056642605a53ecd9ef42a28d4993ddc05272335bcf2e35deee14f0e7cc31539c625315fb71ed93d01b00d2e39073ae78db22c0c6e3a056c0ab96aeebe8ea9f55454b0143f6333eea9bb686e054227495b610e34f391e957a258a3b3964525939fc088d33bb4f8ca12e84f7553a2f0b61db752db541169927a3ed8f2ccfbceacadfc1007feb51028bb7726c9478aac08f7b34a32f68ede57dba1bc0269477ccd8d74c6dd067042e75d657637e02e96109b08fac2ac9ff32297d7bd2790ba5807f93fa2074c3ad2b3614e2e0a0c0b3e3442bceff23987295b9a2306e9aa43e17725e2ec040856affd8be80ccb21ff42248aab90793c381a3549107dbbbf44721138974dd708c23f8f85447e1fc3ee50838eb7cfe9f2b87420d1efae99a6a3f94b1fd715419af87701197110562faa28b8088671e31fa51cead88a5df7db8e4902a637f25ec9770c2a2202e4462df5700383111f03af95d513e12f4993aa0471ed183dc3ff2258562bcadfd3c3f63483ccd0711731e0d54dfcc9564d699d71cb989b63896c22c2c0532ccee349a915c8de40ce1bb6628ef450a1feea415ff81351cd853c8025974023176dc2e2965669830d036376505018f3832f2136fc7ba1c9f8fc7605bb19e783084262d90c5565f2e6a1dac39358b5af66817a2000f21226c904458a844f14f301e3d8287730ecbac38847a6109b24eb40cb58f2d25fcd6ff0c1803d87af13324ef36dca0ac573421b04ca92db2aa87c2b42046f23ef637f272a9bf83eb29f8ff1e9821bc05833410aece80d585ab8a9d1333ed3a81013ae1189c1ed93f56fb909106e7ea2a54f4711efbbbac44e4985ad97c95eb4f414d9acdcc52da6e71fa8aa2b0640da97bf883a3e956ee4d9d606f2ab8754c062e033e852fcf787251cbfced9807bf5f6e492ada0f4b58b604c7882a38843541b69b17a24cbcb9636dd34acd4f0b58d360b9c88fb55328b74f18868198dd8204323d2056641483dd77a19e5ecc2000d4ade85875491250d4d364385a5b2963b7229e0c8a4eb0ffd02f88d845cf3036aa95bbe924b9cd5fc587cf83d1b5f10d7c0384a092d49f3829ca32ccdc930de2ab5cb59992e4bfc28d43f2a3741735dbb85557923733eaa1b6358c9228cfa42cd859b12c16aa6fe875b811a86388e9a895be3b7029216a0210151e3f9f71817ca40383612f0b95798cb00237f7575d4d3ec968e6db09e5e6b6d175aeb03d7260fc786703cc0b7e576fd85f821142feb7e436a2994d246be1c245a043e090e4ad1c5e1756f818457bbe49ee1168e49df6f599db50056eecbdfdc9a52f69bbd346f9ecca4aa91eab1662d603c0240f4d970578faaa9b8331ac58d6a8a4a567b107ae39099425ba7c87fc34c76553f0d6af2e22564196f22a9c7a862badca7ecd5293354e4a5809ca884fa2dd351d0822675d074eed0f315c06b94e6563a2a692c24e5f23929c19758eaeb1811f5bf4865f77775fc69c55fa89ddc5e3650205738f1426520a4a6fe3183700e2b0efd6c3d154cab0b47699a3d3284f113a48818b367f2131ac686be6a7393f9467c4e81630d468c1ad6cb7419d5abe691a8381ec57e56d9f2750549a49035f09130d5d945b7723c9b6faeba52e81043a0875f2125d66bfbdc6ad7792b33075429362da49c12ef2aff4aa611f7aa920f6010cf0098555d65e615f71d9ee6f81c192b23e803e25dd282f15024005141aeb7856fbe92f667fb93d7eec013936de82fd5fca1474a590666077d7e6a918f6a181fb6d6dbacb85b62e2d26e7e69054065e4afa4ea2ce900962659013e8c3790497429e401871b3662bb7a5444f37030a5154505d43db2071a82947f4f55d35a404ca0e0b4a670fbfeb82abfd836ab85a8531a2fef5f25c1a88f0881e3544da226351933504f72636bb11b2751decb11c3236f666635c91310e779de1db16f508753134821fd5b89cd654728a90c3d2f604cea17ca35d9b854a855d19ba2aef904bf085b7cf53ddbff71b473231a0a323f4c096bf8013efad9f7bb2800db10ba8d07b679596ad3d77cd0a81097ffec7ec42b6342b88013564a7c19a611fd883c7d34427eb05264fb0be4b2a559a58b44d3e005606bf032874bc7e858391dd7b64c2899fe42a96fda4d656d3fc40a9349cac279561ac72ce5698aae54db7c0a17f40e441f5cc265bb77208ef1be7c308ceeebbc6ff479b24c26ea94eccc2c308356376e569c5d47138873673261bb9fbc094830f868550389c330e9bef8088e9bb50f9d1ba16248e85af94661d0886f696bae4c803e827dc06cda6d31969a6f28d187a67068a0c54a36200d9336e09dbec3fdc31089d891e70bc169fb1a6d50ebcd7874a183fd8a93bcf80b1e31b017c89db84ba91a9825c845278943ea72347311439121ad3448b70e0b9c588d4b2ae8239a3410f6b878f539eba596838cc8cab874e960c1b3262ce9533cfbb0702f97ce92b95c6154ea6b2b012e490b93db36d9ac2ac3a1b6b308b4f9f03a4b2e782485ab223839f299fe0cb26d1afea338742a2f9c79a08ece40179d2df6c35236f3b44234eeb46822371f506a71e0b233258e03e385405e82de064cc7fed6e8b4aa6a3416c478f54d29faed8cd9bf8305744f0945b8c4fd9bb5f7709b816668d6913dce2e13d8957e47c9b197eb84f23cb7b4ec12bedd15c12364e7354ac7267c3093d3b55f36170a210d8a36d125c0c0fa8120ffc267877c12565a1514b6dc306fe92eb9872569c008a2229ab6684c0d70ed735047a350f12ef65264b648ccf9b6c24bb9ad634745a5f4574cb9c3436cdea7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h86383824c997144e9336fb7cccfb3411653d66e5039cc8f322f7258701680621ac21a80b36876922394988e90b9428ae70633ddd688ed1558fdd8db2e2161cf99bc5c933257cf1861bbf4df905ea2bc3d5a37800d4f51564f57aac09d3d90d18f6d4cf26b6c572607a65e5d2f73717a63c14789f44833c85e176fec682769019df678ff1557786eddb1ae0a61cffb84a04c247e0e79c86824686e78200964f1d98fccd67377da4ebae41fabc1540687946492089e1f4493825b28ce83b5a8212743d1839acf8a0f7dcfd75a02d4fbe58b3ec9f9d31d118dfc7f595440e6844170afb56587c6e8ef7232d2dfd581d1d0b7a4dc6e830626532455c964b80b0bccb14355dd53face8dd12cc2ef6d8f2e513fa448ea46fc0c87231c8b79665b7eb13304fb87aaf436cd3e34fc2f38cb3c263fd97f8bf510f6d33b87d8aaa3e4b27da3d5061910d6914e1c5cf501769178006e4598c51231f3e1c5e5881270f73760b82293a352b14aaa0ea30e23d73891e39fd8fce02697e6f2527529a8d33add0343c06b6deb67be169c05453b35820751ad5974ef8ba07ea0b24c3c898254a0df18478a80341cc0b11f4116d4dd6e8ece77640ef63b64569516964b4a1123beaa745e99285dd3f66cc744b6da0429c6b77b791138a642dc9dc4ec74a6402ef24c275cdfe0b6bad28830d61b9ce1d55cdf2781865d7e9533d2426019a402eb539c61a646dfd06a25b3cf7f9e45f138267801b7e26f2bce5f2a438f6246d6b65714896ca41170e146a1b8476ff3fc1e5a8dcf08c5c161480b565d286754279fd3a842066b037768a24137bf9702bf06885f850ef8d1898387aab7d505fe26c6209b2ecd864b99db32fd080c250f295a0adb74379f307fc43c0a18925192553f43fd2812e990a080aa2a4d4ef95d9acde7d79d9ab3701a6d2acf5e22d2e3f22b969099170af9c242a210b4c6f0f8ff88c85aa290b3ab7834d1e0c9482b9919e147df09edd3ca548bac8e0e9468117042d8ef00d9c3104d0ad835ab9cabdea20c5d20520cb1afbbe1637c3e98a85673fd1dbd950dc8c50751d0679cdd2496417068fccc73a4a604ccdb12e30e2604b2bdff81093f5495333b2e30020b8e3057d84a5d286eadcff2862f0a03e5aaefedb8b08d5340edc226cea9052e1d5453929ce1902656e49440018390e8eceb4e7572f849a3027d1a43f5a5ff305a39a8e28f1229131bc4e3bbf1d46934e050620ecc6fc1f42a690d82e5edf04bc37d7dd3eb29448f20603a52a8458664bafe8f2eb372b205f539b7ee87ffff233513f560fa51413c270f3de6440b3d880ff24c662259ee9143eb6ce3358bd3d36051e13075e7d7132f54145bee9318d6d550e62d656593bfda931dbc0c05606f8ddc572bc3f8a0a9e5fcd3a90e57d5bf6952fab06dad23d9bb20dbe6f657dd6019e77f7e9a9283e5e34460f2fb9e511fd9ace617142e215e08dbeb02f8e2e8b04878c729ef9607c279ba7c985769477cba9824a9fb4f65ad8a19de0a561e7e90c6d8af330ce7b883b34875ddc1cc59559074e83927ad61a0cf82a98b5c38e7700cfee87450e387e658c3c81628a1104a1f2dcbd7d684761f400f62473ff245bc6940759a81e34c70aaad92b344bee7257ad80600af193e4ef1d26f117634c0de8114e621727b6982ed9459e364f1f32a7d52f218488c7a5fbf8777bdfa910a39076cc5aadbb19a536eaebbfb9e5fb3a2c559477c6ef457c61faf398f0ad8153cb6a2d3154c23e24341af36328f3e721ee08e928a1597714d3bba06895d12e862214e11beac7dfc4ca3c7f795ae6d62bc1be95058e0308456cde0b41c559ad5a18ccb2bd1503b7233596c87329aa9b39ee9aeef3867b57266154db2f667cff54f44603f4ee8866429df803b710bcb5d9b8502f31f056844c57ce9c2b41e7117f1220549da8847b3ada5930a351944b64cb9969a70a6edac345c44436eca4f59aa05f6701c4611be521c657b96f6e2f4bdf684fe925b057d6f5b2500b30101b7ed0393e577990f86096824f31c711628ff3610733232e7fb48045344355a1a442f2a65f842b1a12a447dad8c55c2df5fd92124e67fd160c8dc35a3b167249acbc49b78fa37d85cbece76eb440882db03d9a66bbc2fd1672573e83700be083abad441995f87e82a7fd79fb6a4a68a367175ef19aa3c8c91478333d4b81527ea4ec8776d265680b7e484bc8e31a02d275547cfd60d1267c744b307e16fa4f09933183e2af8d8a68da085b43844045be262aab27fa751bd5d93a51e25dcd2b09d0fe07c6925e190da5027354afb6625f5d1050fe4c9ee01fc2342472c9e488409bbefc533d3afe8e7cef5992c8d1591d5772b7e9a13720280315be07ef823769849646abb6295ed202a1946db34973919bea557d9e9bd5004b5fac7071167299916758693b5416fb88b2963b10d0ab8b782baffa91c78928863cb37c41af8102cc037f38b304dd560bd956df5454d9eae6077b442155eea8e4f0a6787c695c8eca1b626c0c59d3d097a6152422d172cacf23b046dc5ec954c5a9a574f66ac490dccb7cbc0e858a22ceaed441d195c0d65e3defb71e1167fde63624fdf40893a648958a882bff0bbf95599f427bd04754da9be31651a55a4239f51a7d20eb9162c04139c8ed8611fb13de1b32b8e85971e9d0065ce44ba6295d1e1400f4d80957968bed063b58a1c5186ee5ea98afc00772bdca2489459ceb74b268e0607da0e63cfb4bd08b5a5ef1528a45145ceed3a02f578b0528280b61d1ddab7019a8f731fc109630d0dfa94d0804a789c0c4d9b08145e88a3b47ddcc233f79d6a6a7b04195187082c5a5c21f9ad90f345ae5b1ba87cb04b000e8e9a0954eb40e106aeb7babf0f140ad52dcf66a22d34bd0ae0f0b8a880c26db21ba685fdc2c5aa95a5ef60ba68e59874de8c8bf24e5e4a3099486d38eb5ffb8df2022005d81bed64f15eb3b078bf41fc9a117591c49e9086fc3192b676be865976c6737969287079d0eb421ce56cc42045ac2486afef0b5fbf78d850ecd058a11e88b5d42c04e70da4eb43fcea77f2ff1fad80acfe4ce5aeb955e9f19daf892a6dced85c444a28f8aaced28e302e8c2eebf13aadbc9ef7b8e2a95348a16547dc4acf5f9c127e3ee95eb12d6668ae92ce7ca00c4ea412785f3199bd800ffbbbe4496828b07b9ef6c866cf704a3b188847cad15791e4944e30f958f4fe9e4b450fbd45430cc8980ccc71a0ba05fc9820d9c8c55109feb0751a0221bcb5c717a6accabec924bb91d53430cf6317c0bb6e171b5c3312319cc1cf0b65496aec9c976e9e7f24d212f6818df9917572b8f27d6ba5ce37d4f465d2b7af47ca686ea4eff877ccca396aa8edffdc08672bf08cae9b02dfb7f26a3e903b3c4ed82f458f98beee6939429ca64b211cde2ed1844edecba64dfc5a92f89de7529d1d7d83961e4b6c85f8d23b0a4ddf0a0269657950e3f6351a4a674268b0e72f562daa4e6865af74e9276649bbd1f0309f6568fbff85b909adcf5b88d297748c98e5e5a6fbc5b3479509e7588da661be19ea6116f9bff705b399c1b7525f14c05063f60669e3394b6ac746d7cad98375dec660d6428b09c308c01698e74c4dfbdda55362584318a11853d3ad3f2328602af21c1aae89dfbc6606b296eff922b14057f08d1d8f480cd503249e76f018694fe15f770adff3e93c241abb2c5c665fd55d14523924e291483769634b7062b6ddb77774fa0174a938959ae99b4db95aa3f6f27bfafa7e8a0ed66e9836180f3cccdac8d7afdb4b332e9515f2118c48b94417e20ee79d4f398acaa0f5fa1df6928a2a805c5be7c6542ee500140270e8adc55fd22c826b9e98e3d9578c6d81c72cf5683ac0d2679107d890c6216b492be443e46ae20c8ecb35bd670bcfe29ae5fe6ffaab45fbf543a17372983e560a6d5a1f2183c3a61771a7ced6419b40fe268585207f81b074295cf9b667006784337743ade2581a38338bfa1c04eeee27356b87a7146835f972dec78c9e4451f7892adf62d69e0db2fbc34c4359812f8fda646a6fdbe7986dc8af2e2611eaccf93b0f896086277912a5dea3753f0746e8623221cd2f066542b6a19f3d836fd6d976bda5aba000b2575387c77d23b1ac64fa3e60d6e8c7b08abc9930cf18f412d7bfdbd287ca30bc814f97d8e3008a1bf67ab7505a3faa094ee55e8266cc89c8f21efbc7e66d47a76476de959d39cc07639ecb5ab33cae2a6f41988c2930d7d21603cab49ec6440da7b44ab150f1649a774f0a570406a2fa1b20f9c21b92e416d40d0a2219d0a91fb5bef6ede38199161c726fe008bb9d621d2abd5e3c0b419f7f00d26fbcf48d421364335395f80c954c93a9fab026b449d7f44bf40136b9dd65a5b889a4c2a6441c3c00c01579aa5a13fe32c8a5405bdc830804905a757194721001ca2370a94379c60abe441bbca3b914e4669e42166e78fb9706de033d6d8b0ff75aca5372043fafb88e23264d350c4d86849bdfae5bb65fc8a6e91b3eb3fe739a017f3e212926c0c3b866db6ed534263e3066cecc9b726c6c22078eec7d73a89cab977ebdcc318b789cc5cb77f959f727a99aa7ea69ae4a7d62386786cfac50267ad68956cacd162a0e0e2cf357727b3e34122898340b13e262c362ccb07c1243e3e7fddf518e235b6223c534bc55c1c36ff302726b2702f0675004f5ac0c640ee9d3d9aea945a9391a424b987ffa3e19eebc89f7815fa442f9458ea226c52dd02cb88804d195c9e4d0ef605a7ec27fe56ede12ab446d1c690b96d1f73b5f78c6a28c7e76563b94461de516fdca77eea3d043e55f1165a49f9072f44bd5798b823b5bb759a8381da5f03cf3d77dfada09f182dec9396cd697cc2c38bba7dfe8b4c41dbcdf47779a9ae24882a2a10cbb3c7d071e7d5bd8e4fa235adffe1f5d388bd91f2c4001c56308532de57f3456965b01a6e5e0e77c8ad03f00e697ea98c5f3c1d850c56deb1e0f88efb7af861cf0c5357d10dc09562e1e4298a4d73e0295741bbe985f53c9487c8573a2b0e765fb3b21e108465454dfe3bf9ed46cdd4e7749f144dc32900dd427a83e1d1a7e615b48dc95b43a1900096f0ee8aa03af22c22b7e88da57e7a57ff8e27b4ff13c606d34349ddbe8079454fe4672f971b6eac83ff10df761a410d8516bb15eed228d152d4141a05cd040f22d46e4060cce098a8fec067e20f2b87ace615f3af3ae82c02d84a504cc0e009f5fd4520c4a77f3ea0bac0b620036636b864094bfbc0b786c1f5f9717286df453fcc14e39d10a8ec1059d1a2e63410d75df22906746af783fa1cd470952f15030cd00b4310066beee990d1db503490ac15f0f49c7d2542b8b161232c0a2cbdadcac26b965d8c0f96ed14f205d2adc4bb3aeadc4016955632b7d5ae94ff16da943113ab7a362aee043f13840216dcd9b72a4b35a64a022bb8bb1ff069c2ac3b7087d9a1baa3670bd80fdf1d54ffc1ed5f33326deb93cf96c9d346c1c0a91c5b37db9ccaf2d141a613c02c6eed7eed6b63973b82dc8879c71f90f24e5fc5c24d6e2c7e4f0899780bb70c5e9be0bf5b5f1a4e69e84730aecc1caff1957d0d1b08ad3d01ed1ac5361e8ad7c523fba1f2b7c639829d24055cd3c2fa5c50ca1680346bb7072f3075fc7bc371e2d60542e90548e6f219cb6d3d0e99f64c75902b15049327e9becf7c7809e5ce024ea790a35359139f227dfcfd4d7315d09b3f3c9a0230b890ad247b3131ff4745dd3cddd2469de59a0b5f56be2294f812b58ab43b15b757d5114235;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf3316292c3ced419b83e8bfb1ed39fe2b38186a527be99b20ed968bd53fdca3b6663b432edf3fe1a2d594e65f641c7fec6916d40668ca4bcf718e37f0d7d398c9cd67929d2930df0a05e504cb46898f66323880494af7e40d733bed9769b5a4730ac7f2c8274df2d01de9bfbd8d01ec575d3abddbdc2a2d5ba2f3e7517945d3b14a1ef297d1d5cd39e9e68a798de110d71ffe5f8619b3685220ce878088cb547e53e7decb3b2f38250c091f23e0b69e37ab2e167ddad003712f1aa8eb891427ef36d272c8d1cc0465c0e016a96813b815275818a1e7d5911fd0e5f151402ecea16d135b4079f9897a1e1cda7189ee17316e62bd1ee0a37b66d10dc8e0495c6b0141b86eb8d62bd62700a0859842922522ddc25631f7ecf748ba4b39a8906116cd679480cc22987a3eebcb0152f1199449147fe992d8de12b4a8ccd698c06d6b6bf1d2a18452bce3ac733777fbde8b4057af329e2f472af3e36e79450860ffa3ae56c0aab83b16aac4c30a8207b35a946eedcc4271e7d88fb91a8a18bf1881bfed9f0f1dedc256f8656dc0298a1a9ac97179c475039dea2f82e85295597a580b37521f5d127465b47aca5b12d9b0ca965d17b62739e5bfa9346c9a1c4ee6bf2ff8a0bd39603fd313f300df04a8f381f2b579c1393fd59c6e72c7ab85dd541234491a8b15a8eea773629edb25ed9160df6c620c274178770262e2b36229a28ee6a76675cabbc5c0cd701cdcc558a2904d3c9bdd1cae015c599d81c44ac094a8cb5531da8bcd290da7f98294b0097ad45bca840a8f074bb01a1d26e700e891c774e3fb3f8507162ecdbf97c9054d4b4e90c59ffd38f2e8a8f2f277286278233db04b781f7650a36b0b5df8a6a0646049609fbef00735f53216bf711c71bdba8ecac97f8608d42eae019018afd1db6541b65681d85ab5d74be792a5bf32554b442de6b6aadf5df00b744be5e06ce59b6f2bbd51c6a970286ffe9dd05174716a842af217ef009f8e415efc2bce44946abfdd8472d51f53410db61bd108ba30a730703e9a829d546a7e5cfb6504025fd6493264aaa0a369caefce27c5680e4e3a362db0c0bff0a5f53b6a1c4fb4bb9bcfb458731224fd5bf761bd6c1f0d148d96f30b26aa5df5f44209ae2cad545d495cb6b36d6f1212dd23cb0f818a0cc01d11bd0407ef6cc405b7d9c053bd97ef0fae1ede3dd17081d643b81346e2c59df9ec2a3714b031ea4b9d829d2a0e3b755541145b6e7d0718668d9664790d9044aa170406ca0b2b76ee4c2cf6de7ce4bcb599fb5e80613f7ef4c50e67fb633fc8e79379c6390b18dd79ab0dd2051ca425af15c1d13ef2b54db3f4395a505f3ad0ee0c2ff2e00881927e38622d5d38a1fbf5ed21c4c9d783898b6c1b4682f4fd44e0805abc0fe4a9af341c81445e4b1e12af91a6e28ea9b25bc3c61027cdfd03022df2a548bc0b49921ea0560606286b5c0486f7b6bacd16b46be549ba2e42ffa7cc2e52f8ff97fcf322ace87c3fab1e3016d4ddff4ef4a7cdeaa70cf750d5c00d3ef7cefac71860fd98cf553c8fdc3122d0ea924bb8904d95c2e270b83d5fe8a15b1494a1b1a71b451eb7e12e977394e347e5baf6048599f2bfa1da3de127f9e2eb22152ccdf104baacd7b5123860b4951b2bec88aa7c2f2c559ac11c41fef804eff5ef87de84e090c37c4bc40e0b454d2f36989601fd4cef6f9e9dd585e93a327d041618e1250263102860f37cf20ed55b64bdd4c5a811ea7cfaefdfdac777248de78056ded4f0dbae56e4dffd54010fdc0e00534478114ae7ba0f6c9e4c0a667a6782aecbfcc14790da5e91d50e8a62cbc370d10b133506c99e1625a2cb50a037f1166f80b98ac9bae69f9cb35d348b287c00fd2c2c7267e881f197081bf822d1ec03916d5e2125e95b0b916a4c74f53799689f84e1b270b63672e3c0e49e5ff36a983dcf7793b0c66834598627f7086b64dc28f519b1d26d6844f220837a792bc09b633ae5eab99367150b7efe1b0b6b43fe915e498c5c9abc10868bf1b135bad8b0e2ba903554e51be78e23d3a46568cc3eae63d2dd733ad580e37959472aed42ae84a5268eeda8aa5580f6c0eb110dba0bcd2cd7a2be24e78559dfab9a3decbb3e6f0fdcbf6d5be0e9fdece8eb35f1e2b7b26968e0e221f21fe19ef1a0c1e046b20bbc6fa928fd9a573b5fceb2630f87d0e7c4d99f6c3e176a870ab37bc46e3e8b045871ae5b8f3e8c9c32a6392ec13d0adc66538325206a3225e3b973566d4f0fb34759609ad68a1e20cedc81ebb7f08eb14d140524e79ef5343e26870501ae565d1f4ab49d0b2db417f895ad6c57f4304cc53734541b568d71acd92e708eb7e91dd4f15b866dc2fce2144c67f5df03308ee960fbf9217a277a0aeb3c581b33716fc8ca35d124d1443a85fc4d31c16744dd9938a8bad509b5c9ebe7183e5a53e028f7c2151ae468e3e6f66907e342a1e505f829a531fa0b40ddb2ebc1482deffbb8721dc619fd26823064470ad2de400c2874e9f9fa70ef6c38a84fc1235914587b745d85bc02d0eb26fddbb08b5e579485b5cd3959f23a430a4b4828bd7ed21f6df69ab99675790189f1fe5ec6450b539d6941e9e1ecda7402a619bca3aedae27a422c8d19b9785e0f2b06954e12a363a2101202a200208d681edc90799e3ed9dafa273950a9eae58dd0a8e186fb0b4f02b9f4cb940abbc232f78336c62e7efa25e693232459766a3ea27783c66681b8769b2168614b7fc27117906f9aa73ed1a6fb198a5f3908a9d9c900abffeb3a731c643bc554119999286d4a92c9a1d43ec038bf963858bd0fb77ee7227b08294e135b0fda10932294b22719be35455e9daac54294749a9e4c1756516bd5b604b90ac751d94f9ce3f5fa11d3a8ae6bded800b610ab4f232bfad2e427f7c9e7b5ce05e5e275f89228a3253bb3a39eea2f7a2dc2ac50c135b1f79bbd3fced9ed60a996b3776611c7ef2e6719c219f8624d6f64c11456eb25a0d968943d40118899dded327fa6fb534852ad7770a5f421ed038114c3d0d6762c16f274c8c510db16a99a0b68133bcf33e922273b10cefc19bbcfcf4278ee0043a893c001e885d7c897f08196641216abb82f7c0e1b8cbbb528f3caffad2e596c0a579e077c88e1b5a020314fff7fe08e0aed2e006a3d2ff3954329c628b401fd02e5ed1098bb6f73a0d5ac4ac1ff3f8741e4264e60a5b3af930e76796f2d4bb3c80dced2649a44d232a906a409e01ea3cc240ac3e249acec92bff9d1dc7a95a733bcb0ef172e9d9f180028be37f0f2733145d25bca3358f4c51d66fbecb1fa34d429c2dadb2a33b2f759feae61cbc1201d11eccbec98ae53cd6225a961767eab5189aeae4374fb8fb3d6b347a18d99f597a66a4c5668e6c8368acb4149ff2455f32b768f86adebf253e713dbc02cbe57f9ac33611e0eea2cdbcf8a818c3e11e292044321d01cb35c5055ce04b1c24793bc0260dd0f68d376d10eaffa6afa1d6ef86a24d2c45c1b4e5be9e1bbcb8638abea58fde24fbd3c7b99bcd1e2a23887ff5c651f7d0ff5cde828cf7bc9b9df818a647b5ef84a1abc4d2a1fbea439dff3b94917af58bea49181ea8e06933487805a581f2e9f093e1720c57ca75f0c2d92b9dca605f5951a62457919deda1cd7c83f11cb8b19370aad5909a379ff14ca80467c4c9cb51ac898ceb606bfc145fd6476d7df67128afa6f74dcab06cdafe7bb6800bdd824b0189e4d1c556c82464871489b6a6e731c6cc31a70ce0a4e37b7d367905db4b0ab80861e0f7081922af012d3896d3c19152798219d85914cb4e981c84c86642b6faa95907aa7cc1af2b6c80e0d0f8d90752e01847f57c49f39074648a6aaf8a36b8c6fcc2b768590aacf640716872041b1d0b2ac56eb3bc3d4d832f4cdc3b1b45660bcadc385930014be9b355cc428e952d12e4cae2710b90d4b0cfd67a442245a484a31b64ebfe80a4690019f8be07d51eb2e45952956693444a92ab14e085618f0cc09e127d9ec125a768eb09a0355c826c0ff795970d8df46c3f5b435ef486b418602f03cf1959858a3beec0d11b8ba7f64f25e336fd313e01e35174ddb7bf75c8e1e444eea3cedf963f29cf8082761ab66fbece8a206d3aba8870f0e972b5c4f7b1c8f6e541362499298a5afb7eefc234ea82fe3375f3bdf54ad92feeffef02eb6a39080be300461571593921b4333b84fce6e3e0e1ea4b639e2663571fbc7025f119c34ec8fcf33f31b1adf821dc25aa060e40c0e2032dde3d840b0e9664d01106c207fa7798e9502cf576624b6be624ab14e81e4bdc5cb1a62c525d75bd894486c03ef0ed4dbd4ce5c79504dd0fd3f6b440549d17cf6e0c6e65c389b37d1c6ef294f77d003fd3c949cecfbe80fdc5c4b1adc9398f4a4ab3e0f3c1d74eea40090537f58d6109b95ea668b70e453cbcc4c27ecabf26e021b4ca39d9b8fa8ee6c7c36c8d7cb7e6ad4d752c8e5f557989502f0bcdeb985de9a65b742883912028f17d22876a82117784721b8ec294ac28b3745fe78511e7347ba81ea0a8080890e03a45792e0b7e3ff2b3d994aab56fc7c289a373bc24f45ad89eb5794fb8b92e9a94c7d80d351887134affe71a1070b7a23798152188c834fa803c7a10c462cb23f5e105b2248d4f522792504506a0e6b39752efa3a7f041b6acc36e9117d9788c9c2a88a8df4c90e3b0b986658f05b66ceda6eb30c16d211c612920b9281a83f9bfe129b9f75a6fe00667011ae354b9356616f650878f962a4ec79497ee4127f384ac051048b43c22c8ef509b61ebbf3e4d966f79a0b350524c54767efdd52e9680bfcc45d937db131ccf4640c0b1b3d886ea4a28919cb44dfc609eceb6e3d3885993484ab8ad9380c65c02d494b33be6dd772e1c7b97454e166fa5a6367793a82519eee3884e200ec19a79a354ebfa20ec5e2a584daee5b1e2fe3a200332444dbd231db74b5eb18c1ded6530e8cb8d52851fc9138b47b2b0a1a80fe64cbe768bf92e51874c59a941f0a6803acbc5f165309796a1151c2de8023b380782e86a87885ec23b0365dbfd543c4112e12410655c799b4e45b7a9eb99d3e18d01b713aa8570034b82804db3e932f080c6da050b23c68f17555cbdd5889fee9c7a5f5db92d84867a29920037f71718b63c7cea14e5fc3ca2c4149cff73b7f93b671e1ddeb7ddbc4c27f9e176851db954cede45a02f9fc60bb5968417a3cb301750c43ed86fc96e155b6e27cb35330e4d410b0836665f34344804983a0d127981120a59acd0d4f971159ebc88d4bdc9393304b4fa74898804e4f2544ccefd65be2c18ca99c2d2908e6eb507af3920c1036466445a578a02a28618108d9818b9989224f846c37c20ddb39fef1478ce1d6f9f531f8ae7f9c4ae331cdd66574bef0b59390c2d205a4170fc96d968df83c8b1b5761eeab641d3e7f71bfa03d8ae03d0317b7e218f73856756b77e05c8a4d8542da5e9de49390549265b91c448d5e118174bcd414668ba8040bfcdf5e485e0b16bd1aa3c503a08ee3b38d776287f7ca10e95fc3616f3f2e99f93abb547ba6ecbbac916b02bf53bdbb84b509082719b115c5882f06bd6e5dfc2dd39638fdd539da09f3b4b30974f0f3e0a30c1fafe91eaf3f8d5666e82fdc08abd3b470de9eedba558fb3cf453162a3b6a6fba7475584f2977ebd1144ad314dc2025e5d893679ac444014a6f5355ec14a22cfc08108dd385b653cba52e2bf175c79f29b071962b0dfa6d86d076c2af789fdbdff2be528617c0a720a56af33778a182d343cc1cbe88e3f8ea7593595a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h13e5ea4f4f8a50041f24faac761e44ec17b4cad85ee39a2e48a47af5bae66ac159d6582a095052f2c82d8bf17804039526af5a1e841048865f0503894adb3db7da7901bce8c76e626c546b097e81a2be473e343b6b963c06c02247739c41c37ab0cfe3a8a087a2f5fd6a627053b6083b272c74c18fad53e9435cd6c8b6f41a06291e174c7d91d6c3f698f2153017d498a31eda08f7d4ce59dcf6b4b949372963fbe8b8b221251c8ce22993cc3b5d19c0d90997ea87c3605c98efced363c89c6c741085039976f5909d5e81fb67322b5c3b04cbb9b29b839ee6f75245c3a52f285cc91121597fab4c1de40135c77f015c2d99efb4107979010548b9df33f8f74b59831ff51e4e68977adcc83a53811630d3ffda3b70969ea72fc3717ae6b86e50b3c44b837b4325d8be2048fef5879ce40401b6e30af2d437e85067aa6d1c179818ed52eabbe4d8c606d591738f78e6ac58562335421b02832c6ed434c18b935f0ff5e0e1c5451421789173b13f07d07c067bf8bf72e6cf885a4f8a697b5043873dc4633967ff70d634578071a042601b93617bd46ca450fe9d259322b5d01ae0f65d86c247ae3f7cbee712a8d40eb00ac93cbad076de989061f832341a1b4303c98a1ed425a653098f547b4b769a02647e13945fb1761aa1d2722b39a93d072995574313f6d7d974f905dce2404409eb960b033432fd6736469e31f7f754dc6e832f51e97b692798d17f65bfd9cea89312a6650ed42adf3a445904e8c184984e1a431178f8288d3ed3f5c7db2a127915631e4e0947c44c2f68ca09e5efee0ec333768f5ac5f5430471317364a04ab42be0c8853a28e44cc7a7721f5d1ce465e691e3a59d0289c9618d85a53fe54e1f6f5c6c9d6ee1a0ff03ec72a0b7241cfa47c04f1d05cc24de75874b3c1e3b71ea343f244e733206d5bfd4a71e52ecb466ce23c61543803153b21468bb8a58509064f110657cee13a3a8921cde718706e5bd9f09447e006b9dd0f049e971b2cb1f35c8e0bb2e96f27aa37a04de43a1d0a9be3bc91a19ddb18819f9b91851a55497547eccf05294a7005d239d606f4dd8dd0a04eba7ae3f28094acd6c98e4c49e1e1e1011b5bd293876c60be0c133b00bd131a9ed06e08e088015708a35f381ac11b1e1e3657dbe86b55026aee42679d86dad44b5a775c4a88883ff4912d76970b3226f2d79593fd20da0f5f1309ee9d78e3c723830b64a88539e6410a960a302d3f737dbf9b012cf63af354799c66400573b82268b33240cc4a25c4fe3a5649451cc4b00f18734213506c843e7bfc4462c7adec1d76a77d0191a6365bf4b5ea54efb78182e2b6ad254167496818bce220f1f45eac24f68b6e73dc92b00cdcb3bf3dd9f78a4961c43f617bb287d2c481496c9fb3cd84cce4fd9619f7dc9ff3d17941a99ee60a5534aeee90335dcdb16c620641062868306d124320f2f57d82b928ecd835652fedca1908edb573a733aabbdc5e036c189058cd205b9dd9dad96f8b715a0f9d4848e2e8cf02c051e6832e88ce644e93aeacb300e35d24f99d1bcd62411576dfe9ab5d63b2ce7701aa9a5ca9f8855f7b571d0a3bf6e21dd6107b5845343e9b9c9884a89b5d7ad78c081fb84ea2981fca21baead795b3fdc2b45058818ac0ebd69f25e46234ef535b94b207ed4fb0a3324aa9853421e64363be9040d8abd2a82be61c98018f8af06b48b2c4fa92b71cb527a866206a557061e4623a0695bd8c37f55c61c1f248eeb6c403a74c67e503403986442f9dccf9b64d05aeeaa666a898421d1d84d77d10ba1cc3533d4b22daa33f0ac49e0c7ca6159b043255bdf15f9ecbd19e0173ac7135f885b444df6b0da1d9a96203f96f8edca371afbaf431729069126625819e85ef07a2d3d194de806806a1e37ded18db7033348f70344fe4780fb73b2dacd4b03d974717b0c16fa753d1f7167fb98b4b1762c2be3a422fa421495e17f35351e933d6ec2895d829e35f0111c3c4840ca98bcf2e09b6a13fca3f230f7129acf64fd3c62b3fdafab5f7e64cb2ea969a0ab02251e1a8e9dd0d335cc6eb2a94ca361161a2a2e9001875007fcb2bd6ee3fee7c99cd013f58a4690d65f8677a1d983c8300449b6facfb429f7257f01c3eb4465db3638b6165884062a8c425c6a64aee4dc9d3deb91dcd50a53959258985fd050172f25047bd94689ec85a76e6dc02d292b553c24c0e8f60d949a1d5ed0ea1cb236f9879ca3d424252a023aa743ed9bb5dfa54f0891e335f842e604b6ddc3ecbde474416bcc87656bea12a54426da54c624543ce3db26b18f2cb18a6794fd37f391b031a8826fe4005fb137e3833baca2519efb7564255d3786cac41a7bcfe6977986f12173788849afced0946b3ddd8c97e2ac117bc31930970dcc964fadb9cdfa1544c4d2c6d0b3a471e63ccaf81fa34dfa6b1f0dbcbc1b9f1a362426e55ad40ac33b420d4dc76e783147198bc5cbdde5c05836cc2dd4df241463866c5cb00e8842d72db494d22708a14da98d6ae3578f6e15095e3101f6613a1c0c8f9aecd63bd2326c7c378f340ca8a1ee6d18f83bce3e195a8b4c6b334d8f132a60da71b9b4c663467e3d812dc0a0fda770bd81c4eb51425e77a280b001c2b131ca099cd00731555032b2fa7409f478f59aac676f6dd26d1c99b42aa7932ba379f87cd5512c2659f0682bbc01e354c3d3466c82b1986a58ebe84106e804f29b1d9a13c76bb3f15eb8ebdee0a85ed64a3676a615a8ad8e14899f71d6dd76bdb4165ffb571bb9cae2b485dc8de2b73b702717198601c4d0b76258a5616347cd2eda35debf3c7ea3f611e5e5352ad333f9673184122f65abda5700dac4af1bca690d94ab62942744361aa1065a9f1c68bf036c57d8e89e08270abb91b9d0a81e1b58c5c7df60ce22919f55e421cc897df135b5d522915550977b8b8466aeae89e4cf0b3cc21d058663a5c60ac69d520117a4db42d8a21ff6025228e81b84c987a19b1fe855bbaeebfe8243c6e58792ac5ea98101ea6c1f368199c21a7414b3fa75058db94e6bb04f3c2d5313e46c554c1f81d3aa152cc64c1c27c1a8993c967263ae145e869f7ad480dd169940a3b1cc6007ea13f6a97f7b30016d6dc8e1f50d5d357ac49d10ee36f152fdaffcbaad1755247b0186bca7d882641c3ea558196860a9f6e6a02f6d4d0ccf5c98e2a87eee9fd9dc3a07e536f171238f2477c1f7f07fe1aaa8dadf80325a011fd88ef7f4690b87d2cf161726def971c4cb102d48befff5cb4f359989602dc385b5a82aa61c642097d87266074f4908a9faa1f10b33f898dec56308b342302b9226bd39da02e01e86260812d3d75d3db687c68531c53c9714f5bcc11861dfd013f95b5698bdb8c0c46cf4fae84977f7cd613cc77da7fb6aeaa59d15007d3210027d1690d1a413c40fbe7c2baf52f7e5732214da4288352341a0ba5b360f104ac935b8d18feb26bf2222635774c072812fba2fd40c1d21a553e3d5abc68a3318ea505bae1c7c618dc95d3fe6d3bbc22c599ca8a9022911b2d14d62b50897d91c1c9a290edbf23ddd69beac7b8e50a55589d16be1d991735ac7a00198cc7dd55bdb89a11cb022d062acf1895251ce0a5ac6284119b533da0ee19a8e666b3ceb1c797d6e8345c01127b4586d8f267d5d631312defe89adb6b4e5f29aca57731554bd9c03a2c4b79084509c359a7d2a5d9c0b3746ae54b79e1b92474f8f0b30b4dc8d77f1036f5f98e35118820f628123e901131442b058c03f21dd2007091cac14e2b6d0009fcf4d7acc44038095c88e6cb8fdfa415ae94e414663a8b2e30d61c0193611ecdc155f89603ab6fc54e3f6218d2a126108f4a84367eb2a4d13fdfc18547ca07be11b0e36804349ebdf07f9e288c314c27ee32d6a478cb42898b618562251c89a6fcf5211c3da631a26f63c20eb19a284ec14ba204a794fa94f7fdeede128ddc2a1022f6386eee7566c432be2bc30ea7c753b28763780476c7b860e5114cf51eb5aa177231977136d9b78703da2f1eacccc54c6a1d6915d1d9a2000e52e23743f67f38fb196293bb2d8bb40d54f427da1b4a0aa63790292ac04a48fd490967249a57e8c7dbfb28575d061570de7edbb4ad1e2be507e5dbefeb4c165d7df194ca17f7dd4691a8df822f2980ab0401c0f1d1ea440400716fee392811ba3030c670e6c1367754b8d1b8e99ce791f750ee57098223cb65dbb05182913796eb17d938765c8f372193a2a5ac5c1fdaa2d9cb63e58deb0587190cae7cb7788e2f2edc80e1e72dcaf84340953a92a898bb643c874a89985bfc0c1bdc1362930816393105e6f94c090a88b5ca64113a44eb952c54eafa9ade274ce89fe2e7060b362905d470a3abb5040fde8f34dd56332386655639c1b70d5f53428022736e5648e812a048d2beab10951f86757e9941f53a748c79004a47547eba5fb6cb0f499b51e95fcc19e2ea229d6ad193e1d0f3616096b1caf5f25f21ff1a37af1293f2448b3538f49f8b1da0a36d8633605567b06ab0746604820da235366757fe0a9ada3d44bb0408f3e91e31fcac218b139f4ff57f351bfba57fd25e53da6a330e62732a4942fe31edb3dfdbc9fd9a43fcfdb25da49356661bd2d231539fd6752b87bfe0982ca0d4a529279b14f04c85d3388060cec2b316f7d6ed95e4ecde197bc7040c9f7c3771c1c4cb9a9811a148c52235dc66e6de14d98a1ad5d3393f043429042d0fa0625dbe75286bc335130a5a6021c079a5c0494f54c5b12de4cdb53b4d85fa837077058ec5d7f36fc68854aae5d08500545a2426e5481eb0bc90641477769e4c65710cbca4400598c89a64ab0782b47825330ca19968409be0fe25b2d6bdb20967da2afdcb05e3d84064f528790b1efb9af74698819a6a0764a9b41ffb4f20d354576d44ff71c965de3fcec50e0097b484d46c5d04826ee7d683c225fdddd0ca1c82c7649b72aecb7302d73c50a55440445269aec64be9e8b08bb3390d74b8ff5634489cea973ac111f357999866a19ca5ce98dcd15de38d7e0b455f7c42919830715175f137c46fbb5d8459d6ae274128875fae79ed0de0dcb85c7afcf2ebac0691a643854cb7157dc1fd90cf134e4a21325b6b59984a9061572bf186643cae039b037f7129ac1c411efb22e56b5651f1dde9cb00b7b82242835bb87f491851739c5b3d0d798427826b07020f8d94707e139164e09c49ae41fbe16995df3b4cf76098e151b991ec4e68d3d6b831aea2f86a4143538e2c72276ea34d053a61faaf9b6048a899cfd5bd8e8dc4f39fdd2a7e419948a61a012549ac642c3e7eaacaf9f1aec4873c3d4ea9b15b017d41460a9535893648c9192fe008faec2852d796af41c1742ee297f15910ffd0bc6362c403c6aa85bcbee3841dd19baf943c2208358002ace4b44af301c939c9d7d1d0469397d8e75ae0b3a4c2c53789e688fc7df8aebeeef4202a688ad079137210b75d45722a3343e16e5d32f476916af39b10620cd3a3cf2dbc7bfdb09e80f8b47b56838815c370ed83c312bf07a06dbf24e5bab3429bc139f01747881d0b0bb4059cb61293ee080be8fc1d2435c364cdd98342d5e99375d07a1ec80f94ed86e40b8c97ab18fc9764eeecfe049b87f45e944919481292ceaf74a79d9b97a9e64eea592cd8676470709f021dc8af418b7e780f9e27250ada49932749ad052feb95946cf0e4e7e67ca9054330e886bcdc6bef25e27a37e4183377823321c8e0ec29254046010650a3dfaf9e36d8e831666fdea23b489b99745944b2ba77c144aefb68b18;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4d767d2a370003c79866a92b8125ef9eaae852d0d3cb826cd41867ee7eaa229a85a08276c9cf7b749831f24a71185015483106982230203c9257c9dd7d4a4736b7bc5df2b9ac0eb2d4494a3974b375b085a37e4cffc5d5751d56868c104b8d33a7658ce85b87b2281c807dc3fe538280f6e6d9b510f5d80b2273563bad8a74196f0e1f97ae86a2a16e8b30e972e6b01761004b7feae197c5d701726fcffafb3263f9a1bb43ba75e29d3cc0a459030e19aecd0e6cd92860359bf993af93c246da40d4e05008868363c94d6db37764927c2f921293afb26daa67096e4ad46841accadfa1dfb26958b1a255f09b2744b59d0dc036a592d2fbd735243303b7a9957130c035c23a609d612dbe34cca201e2751cd8eb928b3c0abf3ce1a0268a74f14e93c8e26f14c3391c26db6da081b7b00457879e175bb7a899b90e28a53f9533b51dd26eed65ca8cc6b3260b4f30011a675e1310a42afec47481be45f5e0addd3d1f5b4ecb61a70a9002e07c8d3fd3d809618ce9b97b25e6553efe0c97bb7fa26e180d20b28f818b0096ae398c47c77d89f5bf8ac342532808cf461a4c11cc2910f39d513dd904000c26443e614ecbadc08a3b85b9d350e52fc8de8c0207ac22aaa4a69ec5409bd591cbc33010a77e0cdf6a4792b9954d4d15d38ccc9f6bab0b38a73a3af4fccaf9bfa463ad27e6f74f23701c8cde56d3584532d2399660f0961a81b84048a07e127eb59693436dc58075d55c49f2a680c2d0f37a1ff48b90a5ed95190da548e1ad9ade3c90eca9b3ce16edbebda74b141c7487f71f2039736cc23f02d62f98c3d3dc5067db03f71514f65c53169006426132e2ff83e8e2d282fa6ba3925f401b3e8cad79cefbfa6cd9e7ef2548a4a35af1f536cb40a5b6c96b20e9b08faca54d822bdc85aaa8301b791c2c1c47e796b244d7024fe73a4f98cf9daaf404e59f5939db75aacdc6550554008587913b5d7e648641cb3b41024b40277ccfb78c7774e12f27f79208a69e3394ac4970deb52a5e607ed7125e743d910d63b5a5524c9bd266ad20683ffa0ea335cb38aec1452bdf7c7abd5e7101141c8da480951d49ac6093170aa1e7512a595fccc9df61eb8f3df47261136bfadd83224503517b29320a77df5e68f1de49f71482293c9460afc639c4b792a93cc8214f4480063b90b8d88f801e7e7a99e6774bafcd4380943c1cd96439681e255b009b66a6318ee91411aa88b47ee7b2cf858518162018613c045902d82d44083cf2aa1099e88937748a8da35a20f9cdd3627d7da85feef9c7c81a94d49a25ee422b5afaadd0e0de9173ae16925a3fa97daff67da75939f7cec9ca837eba6ee3fc861992c162181bccdbbe0b8e96476b8d93f191dc96763da8ec79e82d835c524435dfec7d7e1ae7824142d0efef242018c832d77137e306b30c4359034492085ee3c826e5b608fd266f758d4557bfb5c92dda7ef4415f9b8262a18671b7b85b5f9ed490857b22e39786c5d0cf15073eeb67f1c4fc383bfd7b20f92bc4112f099723d9b0f7d7b4199e27db32ab61d2b1b176ca0e8fcebc5afc784329204a80ffeb8d0a7a480578c89400c50a3b088408eb2f20db63097cd92584d768b02edd9c2fce43f9830cc613073aa83e11872b4cb6570ed4b5594fbf38ac653d8bc2240b2e4be4ec3c980904cccdff83b03c546589d3c9c559959238b2e3878b4557051759202e956dd1056f0a1417a9f1bee5f16dd417031d21f98fdbfead069a8329fca7617cb020659e7b600f355cb7482f9035cf24e3bb01008a4a684d92117ce8ae9df82240cb024388c1a2709de51d8ad98f9a2ee2e8b7a61e6a45b88c32cd5cda78ca925acd1ea38dc15651bfc93f9b852ca8bacb146ddaef0cc899b2b29748b405cb21e2d26a9d1b8507ee44ff675df6dd8ddf62fe255f0669a7f650554fde60f3ecde9d13441f7ee16550392ee75e1788a2a53ef1954b7f59c927ee1e5f31bd6f421c882be9afb1a50209a65f9a0f84e521a82d517d3063f67dc1384133e4fa96939c7587c34bc41ebba4e77a4ed3a135ddf693aaabfd230950d3f556af063a4c691bfa9c9aeb0a40ef90ffedfbbb39152ea52cf9d6135e97bc7477702160a90cb9a0c7e1b4a5d3ffe9b964a0509dae21f94ee99032c7b2851b1c4102d7703a786a3b42ee2269cc4bd4e9a66196dc77e30c95a60a4f2cc32df881c0edc2468631d0fc95912503fc5302363d6840b9a0b3c67b5f2882f0bd29602c3c1d2f9909bd20fb65e0616d4c6abf01ee3efbd986da21480a5a1898496ce81264eda89e431d4a12f48c1aa9a15d6401118a415c9d447f83f12a863a2227fd61dec6b0c989d99ea196d94a5543b56c6643437cec21466b5605e6a234313bfd65a7bb7545e3b42e5193438d51505def641389a1d9eafa8cfea8a1bd440028153672736345a5de6ee26830d2bba83636248196b63ef4136eaeaf591e8961189783ee5a88ba6eff0f674467b90e4c4ebba10114c673093fd5c96e815ccdc9299dbbd3552370ea11848805734ceea3155cd3a1bec4ee4b94d961f72949786a786e819f3e5cd2b4114bab00e2dfa4d6c7c6c1b4ac29a4eb7166268cd32d6b5376deb137326e7c20363aec6eb0063d431f27a279811f86dbf735a97f83e9517ef5c55f9ebc1efe6a115c76d5a448ea18e35849090c7ac785b18769b7a211f85cd7652216e849a3d6414a0d6b20cfb5641308d98f7030c1d79a0711d021da115e6a5a56a3f54be38652523c357022ef46cec47f3c7b0009f3320938a056803d1b71c6f353fb0bff2c20228046f001484f3975f68159641984c258b947ae8e9da33e79663c20c2da16e95a6629db2c651835cef1adbc71abd76098ce7880be288c51f7b6bc6b7ac4f4d5c3e30afc340f197309f7e80ef7e3af3f79b957383ba1f67ce31996c56d5ab2c0069ec0b07410334029116fa67b156d48ed477575753044a6ce049eb8e089e171703823a5546b4115c9a51a9dcfb72d4b277b8f4e1193d963a71808bff759ab06c343a4333fe08a04732d86222c47387e8db8406a6fccfb7153575bb35bd41cbdca851e6a49b770ae4c134c099bebb552574c49d97d492c053ad4a7b38bd9d2b722ca90740d45efee0fec416d826b0845214711b8b29bb83cac7506bf2788b51c0e34f784d3550044f308150f685e9ef805ebc36f72f8c8995d3c86344d8ca1ed4493e2ae3ecb53200b3b713eee9d01836331aa76159fdcf6883546e4bc862317bea5b33df7062e767de30dfeb092dc13f6d186a0f3914d11d86e3db27859c3b7507704dc7ebd3eed2df5e4bfd779d28ee4a2fd91d0079e021f62d14cbbff7a152b50d2f93ea59e3c929d52b58be7d862385e6aa815c2166083ea82e63a901d71bca6d35f6c2ca111b6d6f98499a5bcc66976bb216058bb0f9d0873037ea931ba35b171724fd6e0c781c48cc3fdd9ae336d35f258a34ca12419e071076225c987feb63a3de707796a9465354791cc951150138626e67ffc18498a0b4497c93b600aa51271f908bebe041dbbf7ef604d8301b268fb9987c514fe81f369b11ef5eb20860da1ad549b109dbbb12c009c57f9331ace2d94a8483190940d8d5a62e46a23172a1a94a46c2c78e9a6b3c13ab753d81323d556f7aea041cc1ce1fad6414e5b595c8ba84f0d0ee55b01971d687e0124356792dd6b3e3009bae02e7e21f0c6cd4871043296e628ed1f3b50f1c0cdf3bd0463b78690f0c3c42ed7171e3509dcc978861392067b04c54a691c1e490f858b34bb89870e9957660e46845d05c269269d63da594c3c5e752f5e51604e26115d0b57ac063258c59773c32916a1351f03a3ffcaa3ecba806b01bd650723b8a0ed0173a0e5710e94a0e303a7331360bfd11fc7b6b6491f2577d9bcd213d3a017689263f41f029c78323bfa434b46686353e6779ea7241b5f2cad3d1dfd3d22303d83384dd354cf2df13f86925a255cef45101b95e570e0a0f700be7feece97f86695f165eb62a2ad50d744057529981a31fccd3d95f348c9f6f5dd5139f77e3be323f7218193eb235418de0319854dbe9d8499fa9186c1fb6ee632f720ed1c9e3067e540d0485ea175c36420691ca72e290f8942a275d38b17b63053f6aa19ae17c42ae0bc8e1a3a21e956c77f6565f296f53e792cb1f32dfdd3fa4beb176c42280572c7f098173cf3f49fe995f5bb6adc3330cbadd56d9d17e828ce0663cc2a31a4bd0210fb1e4b10847d24de3506af9057f16d464231dfa0c2473dac2f056e59f138743ea964d22035e1b5d8655851f4a405813219ea1db6e2e4327cdfaf62ca4b65bd351426b3f797e847ad2cfe762511c6c421b29c4aa5843ca74ca5be7de8d0014ad3bf0ae45f1a95acda0f75c458939209a2422bf5b64cdaa03e30f7f2daedc97ef7ae998af8a95cc4550f1d1f671dee89728f0c21881c843bcc41257fe2fe277ad367cde78d6f374ad17052e67c35c62194e6c75dc4c2f18ea4dd692bf5573397b06e38bc4bed5469775d95cbb471966510e0b6ed35516a22bcb7ba74b5af7548141297c89f884a63b86114ec45734602d7e0aaa55c97169efa3b4e09e9a0075513fe0ca4aa83db694421308788d4a805b8eade38979295cbdf1d4c158d5ab2efe397985d4f172b51f29ba7593ea15bb1eb42b5e2a3cd85cf84cdd56089cf84fa2df5641c2c4ec38f62afc855e964333a06211ee67f5bcae08f16b7299c8f11c005e12abd1b6a48f29558c8708f4d65fb21e8756223bcf67430291528c7fa1f396795b8ca7dfac740291970079ac5567e7348aec78043a40d0eb97388fbb458f836518332d80c4108f9499f1973a442f336051c1f5fe9db2763fb22c6d0d37a7606de4d00fb7aa76834c9d4c3255a21a2a7904407ac1fb876ee88c18ac997a84d8733e4ebd57641290a4c5fa9d16b41462b3516ea3cb9218eda2ad5e10f2f8f8263d73359625af17f1b5a601e2398094cbc0a343c5dca6b1a6f2b5a76068830714a6a4e327c5c62ea65814d7bd6a39c2d6008da740cb8e34a9cc717d4cced3b37a078338c152fb63a9568c53b35cfebfcee783029473a228035da275f6fd0c690cbfbe38c7b98af38a8348869b7e23425c0d9f02a4ac837603c50f86fceffadb9093275a8315f038d82a041580177369b4c386fa57d295959a4d56155bfded670caa19b929778c4f2319a776e24fd62c770f3a81adfbeb93abd560c657a596b74b29c32c56458d9566496a37808a27a7c7434415b21f766197ae11d6b2ea3d2b4f3d0c4085757a95417e0d09a72571b0902a7f97052cf59e9cb58ca399a06cba1aa9ec46e71325d93aaafa439734ec5db1488449225e9f6c73ad3ba31e77ab5a5e28ebedc3b2ab7a5aa032a621e14f3f36bd5598ec2566b01976c40cfe37964fdab7147879a89ac6ee772e038a077b1c882ab0a904854beec1dfbbd6a854ae4f371a50bb2b29c247956ec32d96530cdd331b311283170aa844651b0cd050e32374d6ff08cd1323f9e7ba02ed70cc737f32c4e270929b50fda4c3fa8d6fdc99316a3a956b5f3ca743b13c32a88bd75be8d47b157cd823e34b7099103ead46d7059d1909e87cbb1276659cf4ec34da4430adf80f7188b23c2bd6f2e4201ed3d0858ad5126ed67e77051b449f051a0a1065897a8273187b1abeb60a40a9f7b4cc1ef2806f299e33fdaac69200d500082839671a7a5435d8a4f872761bc10e1e59b52a7d1496ca05ee6548b4f1964dc39056c476157a9efa6af00165e91f4a6612574fd2b22fd55f484de0db7dc74a193;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h512ea8b7ad4dcf578243c1c556d5752b54e4a776020187ea7d2464131f3ea34702fdb18761d5a2335ce4d25efff24d531bf304dc1ac44cde6a9f01caf875edc188346333cf81ca7200adc806369aeb8781ada65b8f218e4725d8882cc206c97690bac4421d5ebfeac5f52b50b597df2281fd2ba55b8e2657b435039070d36288dd8d97dc6b844ad2b43158c02e96a8c3affc056c2c6b9545598d7b6eed3a646d2f63c38058095352257d6f8e10b3bb4dabb7ab492928f4dbe0cd44663d6b37ae2b5f08c1e12149eddf92d6cb31909b661a0a2a86bb1a14367c2c95cd484f6cc1bb1d5db091d662dbdbd7799469e3e8376cece949000d1fbbefe82b9077c147b896f338c05e132842a6b55befee07e319663f50e1bfeb7dabfc3dca4cf55128295f35355cc7eb2284ded5411c453df3cd30a3ccc9fa5bb48195deb31790ecace3ad44a4441da6d7f0addd46c130ce07cb58893d4cd42fde4c5dbc42db801af44a58561db8d04c23d122802b7d388fe72bc2025d43f10a81f4f8605ebdd150c5f38f3643cf937e6fc8c94b4588444ac7174634f8419ccf88e61f9161edb62de14f0cf8e1db969ec9bed6dbb489dfb2d0b1eb7c46592e7b521bfeac98a22dd5d128f601cb2b44fb20cec7a742791e4462e14e421a3ad289f5f2ff6a7946082528c198e8363cb504e3562c73cb2e780e95486975465336d698b01fdd7572208b5dfba33a7860fc3ee8026262096a3ec1a34b862db62ca2a7d383530232764a8d1612a044244a6ae082e6d78c892a6925e7cd417a17476c3b520ff8180f86c1788e0769c2c2befa599bacf6c9e3266fc088936b346c424b9196662777738c50ebecd82165ae8b939876497846946bfb728e9739f35ff94b6bad0063ac176ebf0f244b8a8117ea01d39b8e2a654e13e9782fcfe2a318612eab82dfbbc6eadc02b0868a2f5d85cc6d53e907a3f1c514fa318182ca70a77ebc47bb9938fae4f12541671a4ab58940feb107c86a2cfed03e87990127eb03f21ee35c3525f4ce80262de6e7adcbb2c9a56def8608d91294f980dcf8657204649d048e245891c73272d9e639d225f18e5e248f0def2612bb11fe906db1643026e8de4578631e545f792aaa20cc04c1f0617a4e10fd7178d2e364fee2029901c22b70905093e5956502ed114737af5a7c96c4d48ddc7c9f563060b61afc0d486ab23528231088b781ddf61b41ea405e9b5170e7b67493f1b4ab9f0acb57c81e10b9d69fc7b2c1aa993429e65f738c4808a5aab98e78e7a7f69aac2a0cd11f3b34bdfa1d4b832fc58083b3eaa6580ad11cf832b51d9e915e44585c2f750cc132b295127ffe427d9b9cf899d62eb78bdac1e2411b032c307fe67a1d2165422207fa8c2a56e8a6e33a2b10303729b42b914bf4e1fd3db043c06b1e23ef7213d4dd5fbd93576549ef8830b7c60a26adbf8da7d2c610a0a4682f74fa8674e387fcd827407855cb55eb2246c52d64f69de2adfeb671868bccf31f5e94cba31f9383b3e03221800849bda56f6fba4e7dbd1d1c24fe3ded92ed6fb5f920bc391ba8ad3214efa15fb80c920f9e8bb0a2370b3ac5a8bc1c25e4f7f32baae5657d8a477e8cec2cbf0e199a5f81631d51288e48ab1b8eb5ce5a58b9e841a7eb80d167e75e2e64108f10d830e77d51634b10a0123ef53bd0e1a33b76c7093de538217f16b7d66a541d7646c3c45ecdfe7eafe5260d9421c3ea726a1fa7edd23c3ac08732011cac0ba09695eb3c66ceb09093f714450e18824cda188e1efd10b509300f6bdbbd69e894cb9d276a1e5524c15c234ab0aec3c5e1839077d8bc50f6caf0e360d4d102b561ffd6cc08f29a358c95cb42238a51f64fef3b2f189626a0789c7e69190b127624c8df819e50c629f4aeee3fbd2c3b78135e7caa329f6adc6cccf25fd8ee2d0d6d3ff9df675f4b53409579f3c5d6b9cdd80d2b833fdaec0eb06ce0dd0f895bcbf492fe60a4ea33185f1c51e702add241ed669321743558b913770b37693b39147bfc730fc666ba10d97cb8e03d754d059a2642897303098be59081d79f03ccae829cd09bfde7b52046ea8ba069f6bc2dbc07fc12e582d3b7432dd82cfd81be1b79e7a77ad6fddeed2722653597b7b616019650d8b29498669d069dfdadf52206096cf73698f11cc97bff2a3b8f20524f66b6605781352e70fcbaa1e5b4146d721584b9b4e0b135b6ceee81fc6918c3829fef207b7f285c285820d71af86edb851329c71430d45cbcf3f651f78aeb5df8183c09cfcfa445ea84ceb2437f3261468cc2db96e404246aecdcbef74a053ea104fe1b0780fd00fe4e53740513dfded34678eb834f6a4e30fb6d02d45e6899d49b8a9b1be097415b60b16d8b6ec0790048c0729b8a9af343aac9785181678cb06301f8ae7408dc60b89a3c18b9393f7d26df06f02b63772cfc9a9185a138b4b6666d45e20eda8e15ab9032e813b28b81727ee3d71ba1728f14ac311c8395cb6fccf238ed2e34e2e7dc174fef6254285cc685fb0fde837c85b00eb9f517919203d18504afe2cbc09e04053aa6dfe4c76cdbd80cd15c0203b5ba8fbbba1033d819ea460bf7f076839f25ac253e0c74f299e3c8355069199825520b9fa7a369bd65f951637afe4c9dafe8fafe7d272bc368ed8f3a269723fcf801231e417338656691ef2f5a53fc3320395a4cefdf400d2c7b9e494b1112a8588fd7a2b2f5b06eaa5f9cf820449de3694110ae11e00da1eae287ab2dcfe63acfc8bad82ee54a8f323c822511327dd03558da7b00402c379bee61cdfc2cfc87f889d156a828341f7099b4a7f0dc88ff35f063442ce7e3f3c635cb3862185d595158afa99385544571e0e1f1b633d003b39754af2a3556e2e0f5a3c1a10a8c270c7b1b2f1bc032643cbdf53765363d63818426bf3a8b03c7f0e7b37c423fadf9c1b6d5fe409503d1f323e7546216df5131e1b28fb8b9d0a1b7b8f96fc0d7a627396fb490322ffc00fc5e755490a78c1ffbba659e45ed2e75b3c20d19c2ea4a484a235d64db92112c930cde81ff978fbac292f248bd07c1e66d87912b3f10bfb27b7b289f8c8c554b09fc3b1289c0100c3b106b1f5aef4df439bd25fa16ada1776a6e893a662d4fd937858811adc73849ae8188e953c18d83b37940ddb85c53d75da54d49e01092712eb579bd640c38ed23b7c11bc9a6fa913263976bb6f47189766202918013bf5566aa7c39ad89394f66ae0ace6993ab060d97e97824766b64cd143fc93633308653f54bed839af9b6872519e0afb86a7ea8489b56f4a615b693d5e778aa406fbe6fa48a76a113fbd628ed5ef7e6e2c7eef4c1abb592f7e84df040b3d7a456e8fbefd83f55355ea76b4b424732ffc6703faa22607dbeb6760e3c484c9cb27c7fa06935b474ff1aa74079a5711f82eb8837da6937be12ef4510f6e6ec945a35f82f934d36efd3075215bed9dac56b2aae53fe9facc3cbf7c97894ff4d09834e27b4b60823ee75831d934b747479eab3fbfa5cd9c6164ed174596e1cc322bfe069054cd4b6e62b215062ddb9257737f19e86d7247dcd3057dec53baa274d92de90ad01c2055808d43aff68f9e6efc94063dbea35d26206fd7d52137a21e77684437209f532e3f8d567517ccfe419a5ada3e4e0ac61951392a77df197dcdb74b64c03d657ba5fdedcef2e0b39b0c7f76b69a380fabda7ddf3774ae91cf5ae7fa8442f397ef76d62f16a89c16b8f15d86d25bad804c32698d562a4b984438b0d45f770ee493e30f0cccd70d47a4de2682d73ef137e73ddbd98725805a445acf8d11492024a927f0efeefdc8edf2188bf7746f14aa1b3e237af3f71c6c4fe78b16ae1f229424d7ffab2aeda1a2315592fb35c4652a81b288d513a6d685d8ce1196aa731cc3ba46f7b46de2284e4bb805efc5266ff7fd8cda34b3923af8d9d318e659bebcf6f9399c10ef02c2164b26f246817f1783d47efb6d3e8e04ef00a845a8fa6c9dc058f168d6cf5a9c91c412e0b0cebcdd01bd178bf3102e88f1d8d140024daa0e04e1eca056dffd4b841ec227f1f2666008f6d389f2765d830a8e61e4505358050310ea4881c143d7d409d98aba0487167fe322fa52aab026163d741244059991cc125704251c76c5b8137ca73cb5a43ea9b054427938e815e2b2c1d527e4cda3075c36a6410e0415d8784e662e456087963cdc9071ca80211dab063a24f201f20be794d4d435360c2fb973d469de31b544f97da628211183b751f8dd8267c47e2ddf289abb86a9d6d116c979f4d23034c2282adc3889bab2952b680330ba1a9f277717d12cab7af6578b2ca09630e975aeeff1cf52f9dbf49f602e22ca26fdfedc82d29b440c5008ad0def20ea8ae08c00de20186f0c791512aec08ae69f8561835431337a786995f323cbc9407ec56f74e3239d07e209383fbd75696e5b24d4550792bd57dbe672425b57e61bdedb61c5bd951463f51c5ea71a9a951b271922cd84972f268baa7c33bc1425908212ceff52afc0786698bae580eeba082c794a2518640ab889e8b539705ff3af229ffb2322c431446aa8812c4d59bbbd9be6be436183d3698bf3e3ec194ab294f88049519b082f410d968f6a84acebd119a9a7718bef1ffbd8ffa6bf29bb4706826dd2921d32ad127b19e466df04e373804f1a72b67c996cd553fa222a08efe540a26f2c0fda25277827fcb97fc7be70cf9246f2b04a72ad0e559fb68b5f321a9e561ee84e771c30066eab2aa8a4deb2f18ffe0c09e0568961b78cf46c83ece06e84bc80b0f22720ae3586183c7d3ff5977ed32d8885ca2522ef3236df116c3dbe43791a1541c03b0d0144c1878e2124d8453363d0b5447a9fbb8209aa7b4791b238b62e0e79716e15becd860d9d7e0148f3727b2c229a0395b6b73bd032404cf8217a29dfa97629529204d642fcd8f932f1a064cdb4a6db03bd2e2dfc0f271ab07cecbe329a37512bb9c026c09e446c3e133e31ed42e6e39de19655a0a33f31b35921f8de64ee96da00aceaea3fdc7d06c87055a877fd65a9f5560c3fb4a2f833fca4acc2cb1d3844e44c1505163b0560abb2de513c598f2a4ea3edb883684ab9b50a9177ba24632bb24ea236c51d71a105f4507a094c60a217c124d0c16122ba6dd937b149491cec39b92f323da2e13d60b77c42753660da6f3ff169896cb09d44ee5e99c1348fd2ff2ad28764d347b3594e5d4537c0159bf91d1ccee6b3f3be2db1c79d772c29e08be778e2154f4345c31926e02ad86ecd3dfae005400b0957ace3b30e2d87da1ebe2246ffb506f9e1bbfd4fac505d889d7d5d0a8ae040292bc17be1a9042124f425e9d0124a937bffd205c09b064e972e0c7ea817e1e6266aab370e59f7bdf97b044a734caedc882fe96207188dad01907c7cb78d436fdce6235ff31683cf169cfa0b737db08289cf834f756f0ffdfd9214cbab4521ab54f193410f9fc2f8e838429fddc073e2ebacd422e4e11ef3d58a43cf117c9ec0007b3924a9942b2933ed37122a5ebdf4365653a72bdc5ace65a0ab75e539748a036f01930a135804d5e3efde6fe80a3f3e3fc1c2ba6d6dbceab25a9b683b67862826f9cc764b0186d222804535742dce42866b0d905b4fe8b74ba0acbf52be3cece762c0b27a9ffe2c2f27680f1aaf77528b2714c30a7bef670913fa1711d8737fb59d1ab6a16445e3e83dcf9ff4bfb548817620d43ce04209c2911c2d088d83eca8996f7f69b2c8b4be4d181a65b12da3b193fe24cb747ea0a885bb5e98cfad9fcd0838c6ec99c84d006a9bec667ee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9f4a0929a0b0c7a03656967a9d807aa65acc7da1ee8e9e10451b2afb409c058bd8f38d9b0070093153fe1e0fcff902eafab90df7a20e2a9164daa93f8814af31d6249ff59ea5aa516c67ad1332fb7d0f2d8484030e8cb5616bfb07cd0b9aaa26846e5d98b2010f430bffbbfd4c7862fe6ebdec21a1edd4855678cbdde25ac9bd9cbac68665777777a7cd4e52e440293e85c303494376ab05ef007efc23a996834e996c9f8d82849ff6ca4ad50e29747a24e219517d4a49d2beff61525be0e618dfd37dbcf5430bfe8ac213918ec71b4c8052aafca342937535756ced9bc3a1556b8366925c6adc603c6f256fda6fb0233d1276f72f29e33efdde84315192e6c1bde3da126bfd5a9055ce03cba70f77f8a3576610e03f64175f65116e5377878407693a375022215479eb61b288a5c691f868a1ed6381a90f51c020eb35a693401512752f95d2674643a431e1d424b47515aa7353a84d3cb79687e4ba54e5ae0505ee4cfd94ea284882606567af4e580d47efcf96b260ab9ae06b250fc1bce3f07fcffe10de047c3da2f15c7e39ecb7c395c52a9e218d62ebb7ae1561c261ad8e87ea49e490406848a0891d7421711e0c5dec18d4466211c73bc507d0cdc37274ab33489af78abdae313c3ee24860232d58da104dd2997994182d8c8bf2660bc37885c9b0a533729e39bcb69c14be50fe6d440b50c02453410e29d848130a9cae0b5d4e31c9a7f3a59beca0dfcf34daa21731e84b395aa51c5405685155b7052c8fbf361e46f42d351056d67624eeff4766178eae21aef2cca304db54ea6e8ba7e4486479f1e5130aec473bdda1637d987e66c3229a5a86be8468f0c8e336074c0d56e0ad1d5257389805893617fc331815c1bf3e6e8cfaa90db4231a8cd5bdb9aa65d4582743c9d4790f89e68d1dccda0779038686b36fb9b12aeac38e7241f3624ba421dd3812c8379e943f2a23115d075ce2341f0244383efd2e88ff9895195595b4931183d7f7a8d8119fefc16c835944e92b6a7b8cab0d68879619118dc6e28a5d61e9e966f9ab48f9c7c83ef3b98e25d23e2010ccbf1e70a98d1be13daedcd4af914159bac37ba7724a18032045c6efec45487affb72f4f005d413ffe66050839e82b0853744b133c63d080ca7f87f3843f0141b35e57fdd39e6bbd8b77883368e6290c7325751b4c80cc032b9db1af292bb40af3f25895562d532f8149d60b03a1215fe4843dd8dafaace4994a5c836fbd991d318b3669b52b87a21b174446dee01a4ecc2c48d3b45c51b2cfbe0c304cd06fd60c52afa6a22ef589d89ab02ad9a710b71dfabd35b9a10a963f284cccb22bf67eab1a2b8689e40bc69e741020103403bbdbff73f52803ca6a9f30726dbaebf85678288556dd66df71f95b5348e87887017850b36611dfff7b2749b47ec9c6434e1672b984fee3d5a9e9430bd9eaef9634d61b5e4cefcd5bed933da4351775e4938a13fd5ee9ec68df4c5482b62518c77cd3bc6ebbec3b74a87337fc6a1105c935692567984fea3e48c9010bbc8c074d51d0052253c1fed684a5e616a98694682878d0653b8ee2b0aed9947bc5d97348f1699757eaec25806c3242ae85e2399348b96003e29ed4ef69159edcb2beaa92984f2bc0dcb2229be38b399083028b7aed7eeb76d7523b4334a511e4ce401d99446b1acc5eb3783ea0e7efa5fdb60b9945e1fee0263cb4975f68a854a2a9ffe867faa1e6b1dc165b7cce22191b977dcafad2f770048dd34f3e3287fc495dcbfb57666026aa73032c50a63b5a8b906ff412c7010a269a8f71f2a3bc8bacffb9a408eea0766cc159c9b138662b156de644627a8241dd9dc2b26e257fef1221eadc756f476bfa12549d95bd4a3ff3c45b5a78d085a80157b792b041b5aaa560d9a43ef241d0c352893cca7baddaebe63b58c05b0552d1849564b620647340eaf1440777e2ce01c8cd25550530cee5fbd1d13a36fc46b8f5fd606264961e7eaffaf11118dabb53e39c5c68cbd095ee18bb6d2fea1ce0b1a4c8df893b6d3f519ac9dbe6db1a624d9799452e1afaecc988dd140d491125b99a9d787fe2b32e1eefb6f3be12635dc6941300993ed2742089f2cc011247dc29b072e559aed405179f3c340b4f8460709075778f9f5c4fb1e9cf6a7fdc56a93e8eb7d4b738c7dbaee6a10e60e6137aae92f149a7ed3870dd36fe6ce47934a2e515deb8cfbb41d61f9d6f9f89ba3e02790d8c7c1a664734e2cb493a492dadb7d360675a9b14df7e662d1c9b523abecd692ccc017f4b3f466030e3a9273236d9d80014f589347aa9ecf15431a5a82ae10bec74f4b552b452f3657b652eaf2a4498d85f341dd855e7e75755f3e0c7ec4844ac9c62740233950665849563682a1def4678878fbb8c6e4f6f4a8af26c5ff757df4d61ec0cb7b309c37596b2dd8b5ba62af17fbf63f864d9d0946f25d55ba216313717f125790dd0abe47548a87a2af8bb706f82b5ca0dcb3f99e4e6fdedb22878e0b935e442764ce4b591e762760905e47f883ed65f5a7b16e642e93da72ab4dbfa7df353a309a10f5f69e118efeacf16468ccafc07ddfb778edb2bb69db5350c105f721f2b4ed12e028d276a618552823fa464fbb3305d3d94f25a93a273411a06423f2af8bb006b71739fbc731f36f880330a048df9766e3c649f14caf56ad00f09fdf2898be883d3f1d4d4f07ace2a158248868e3d8d469c0b8de4fb89074b5b5ee7afa80d412fa8ea712608db4a65d9ac4176012398468135391f3f5c0b7c0b8c6080fe117c9428df13514208b0164e15a5083adc7c9592a669e3ed5c7742857378f1940ba139e2fe273ec46bc71acf0a9ba18687fe2d005a7002106f655ce7dfa3829150ec71dc120d6c624e8cd972b12b041e9901f32565b492a84b93d64d01c595a0ca53e0dc943cb1bed087eb102feae5585603be7cd08487482ff82b8837ca1aca25dda2273c5e5d3869695dc27196da8c67ed9ce983c4f972b41f740da47e7031b4b88227b54f696fe07ed927180bd3786668b92f51ec33e8e0fb646dbabf33a80fccdb87c59edf873b15d09641916eee91ff077969fb5644625b2d1e3e55f7b30a54794c536e6f8f0a60e925b1580ddbc1b8b88799fa217f3f11f102c27d0fe45b9632b6ebb4d2b1b5e7bb95ba662f8d2e861b10631e62a8c1a9b3e59293b4141a6408da91fd2318db81021e301c9eac26f1828dc4ba3a5803faddaaed6ae44397281063850273a70f43bcc09340174d6593ac1cff7d83ccb655c4bf6115f968997311667aebacec7e90d6a57bb23895764347f68e0e238eff6c333fb67c725cc1adcfede3b369a428c5db1c33112c05f2efdc5589c590c3359f7a4cef3735d96fb18a4f0040037fc2590a22261fc192545ce0654c635af86618b72c3f2808461fc29849102d1bc8c867629e67543f183ce2c36a1f1b8462082843c539aa3a10131ba2c6941328cadcaf6a4ab978b3c6241a443b81ccdd7b4e703bc7a2df750c52c0bf953f4c43740dad183a47ae312bd3c6474215ee36f8107e4e0e1ed1f0e1a8e1f3960e262d5d72435a910a26474ff93ebc3697228f313f1ffae52bd78d4d511612986149b5f0a11af2407f2da17415ecda6bf8360ef1a5ead3ec48cd93ea3b94f2355a62bc5f06afe8a673f9a7c50802f5270dd55f33cecb13f7d59a412843ae5a25822c2aa0b25baceea873eb52136195eed94c6eed96e9b990e7428be5fd79aa051743906edcaf7f414f3211050d76938e9f14f4db9ab9fec4ee5f6ce25d06ac03af0588b987ffbb79c8c66ebdbf46b763fcbd804b9dbacb5e1a0e2b2dc9f869b102d6af830ecfe6549f93332003cce7378a398f83480ab3ab96879addcd4483344103fad6d60b07f179ce8425903f4a94a57e2c0ebb975f9c976b4ae803d47899cb0e5d3b86b75653217a66984a640d5b9a48d64fba100c9da973074c4ba953082df94038b62baa3e7dafdc474ae85e3a7eca3f23935eaf0acb0b0eb27c576dfc24ff9063c3a8c1527dd1f7a7ba4d02ed33cf8907a41a45a563d6f2afebc8ded39405a36f2168cf61eca6e669c488731cf27e5a2f839ac1fc058c8675e10c7b0f9661572ba088d8c8e1a80e9a57fd61800e0f2c199552919a7d9a780a93e77835ef397410921f31eebe6a4b89e3a9b3e2039067553e035d29e35917a19711c063dd046f9412ee6c86c746152a2254f6f2a94afc42f988bcf4b1119d49786921c16049beaa6941f30b13d06fbfafabdb733f3012abc3a0d07f3beaa77870a0b3862d1519a292d8b233aa8135b2b6add0e4dd8499900e14c31a9b32f2c24ac1de0e551a55e6d42e0bb74b5ccee93a77700ee5c512f52a6e7479575559b4472ebc69fb702be6f0e5bb68b7502c5ae939a5510b2d4824845b9e28746eb1c152c355a2e1e14b801e53932b2733f97e8781bd7a7a183e4486bf7e5b482716dca7f19d0600d6671e5f59533fd6122ff2f8e0e94489ea57a700a6ee245f562d73b43436f71041c4b936eced7a66103d3ad41c5bccc56bc7e50f2533f8ef1ad611ad24abfc57645f46a46026f124972482f210268d121fddfd9a251f0456843d6b670ddeed8b536a4c23d158c3545f1b030bcf86d2d3cf45420e19ec988254be365fdc368584f24267caf379cd681943d9eb40b4c1c2471d915168304682d9431e3ffb3134547277fa35493706708d406f345c3fe8ca6a725581f2c2c996927a63137d5b6811efd5c3ad03401164a2aa639fb27d87eead1f2c104a6509a0441b19586feae199aec6a1304173c155753901409717b4e16869362aea24e793396c1c329c710982bdc01d054aca8a63cbb8c7f89ff4771e861bbbcc8fecef883277e90ec62caef35cd5b5297a8e6ac473c518a673b45d9968071cbd7ae911e892be4992ef339199ad1f5634e3fb0eb6726da52ec8a0529454ee81686990eac25b970f79dcda4a3e8f9b054c4ca9e73470a58d0e56b45a0c5100013e608811f6b3716d3123a6e85c72371a78c20ee47a1b81203c87989b3a83bf86a79e2698d6b23bb517c4f4a97dcebf969856e891961d23d0f80f15b5db3b0501a91bf3b4b95a746a3dff11a7fd8719210e8004b1dd95ca0189d535feb7c1358ce36a62d959967eee9240e6bf78c33ff1cd098f19488f9a1fa6c07829f3d4b13ceae82fdb91e85e7bb3767096780184ce248388f5257ec7731b2e32ee7841fa11a1792ce0bd5a85edfd7be0b6d828d5651c04deeb47f6c09db0eda14ac0389211e2f40a37e81310143b8f14891b35abce25970b40f6717bb248503185b2f1cd2e91a6ba91616048c533193d41f204cf6ba0b817adc89608cd27f4e9998363fdf40501f1af72803bfcc85707f3fbb8f895ae7e84491f2a9ce1d83e479c4f48432d55852cf42ba9ac0d96a7227c5bd1a2d644454ebcaa6d5f9a269a49afe5a543c6ad464a9353f0ba29fdc0d0ead2e2b20528215b32b26846ea12a78baf52de8ef0aa6adee228fb8cd43bcec874e07dab0d796b95935b3dafcd8a33c6d7bc0acb3edc7a5709cc643deade29d0e8c6e761ea2fa383ac5ab23a03ed46fe1a38bbf02b246c4730acff27e28b4ae03916efe52a36b47a314f14051dea128c485d66fd50272322da1e43b65de5c8438ae42a5f29b1491590ef581aae83ae42869ca1a2fde57ac6bc83c173ad25f407ca4b7204e5f0fa05f5cadaa9c5b878a289188cf6180086175246afae8813d86a968e3a2b439c30974db037152a0b6a1628f71decbec41ee527627de4fd04e54bb37fe99048363196ce063b5a2e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h694476c7d4d2fd2ad7e77f561dff141eace3033fd46172a4ad3edfa2acbb54b9368dfa3364cb532a73d0163fc7468eed42e3f2ab095705444f677a8785a609c3d0ebeb031713a99a2e77cae3ccec8f4ff870d25c176820ce74751f85af3eba71a4bdc54b9e0cdbbfe47c3567a4b42ef9b2f557747482a14a70a517c524ed1bc47e66ed11f9a5dc59b738e06f3b28a4bb2a7147c5824c33851e74386b3b9468d099a4e31585a14d86221236846ddd6efca0bc1019fab44df44f7c94f9385fd10f4f1bea3fb31f9d48e18f9783b262d59fd1ef5be551f2931f2c0a87d238b118663392f3969ac6046e213ae601377739445be75800a376dcbab6a7a15a39dee8c34d1ec2d8a9b4864b81749ad9c312c849d0326830f1d1a10ebdb7e5d8ed6404f0ba079e730e1d13229359946aa4fa23e391d0b3da9ddf97fe31e774ab96b38562589954bf9bc2dc7643932de21be62fff59a59b93737df2c5777c20dd65a0594821d0d543926392b6843fcb587db3a749fcbe18fbce140033fda1f47da4ff7e7592ba5492dbe6619a2bc5220a977c92254cec67599048072a399a1c75f5a671468c5eaf7aa9d3ec06c0840603791d3fcc96fb0b7906769deaf2afe77ae3dfbfb84fe44a6dd9a4bccc0aabbec55da682c4ddf8c21d2e2a15aced8c8bf85267f0390785daad68172355d57597f27a7971fd40d7384cf2fdb7d8b5b09ec8628a2de014fb6b9feac1eebca6a2ef24fd530aa5dfd47dfc2931c925516cd1e15838f628fe46f9b402ad16954368853c73b7b28171e10b859376ec0591a6898d609ae6f29f91f24a0c616204a03394596cd9b616c327ea346909ee29f2359f2d4e8a34218a6413bd8e1269a229b15ec0a64a24016e3712d0f058729ba10a722118f80460f90a60d761eb07e046877f6a24bec09bdcba57a255b935c2f185c52ff8b3dbc7ba3f37b3d69518ed7cf52e4587846dbd68b928de54cc7095b8a8466c7f6081d1b0d0db94e2a1175802bfbd341d4f572a38ac126f13fb7af19cf24c62ac7393ab24842beef4386b591d929132a9a7d8fabfa60a7e98332578d778d18498977809d2f8d142976ea344bf940df0b915260ce10f9bcaad23e7cb3767bbbbc43ada3d5923897d1a9b829f7fb86da4462f17b3aa88e0f8f5b247e430b3028709e3c1bf89bfcbad37f0dc09d88c26dcaf007946cc11aecaa1a6b0a0f01597643095d6a3f8061c475856bc65f885f7b440027b3fa6707563573688acc34f6762b8d32d02bce81ca3e0ebb25373e207d5e62c367103461c7f2f1d80deff0efb23d21a2cdec820245eaf4e11a73a0ee0f9cc346799b3be83d46b145a1fd0838a853fb7d921127db9edc2ada88314e97b093b2878eb1d3d8d5215b65fd4a0072410fd1bae0c43be00ab752079430f3e3fefa375e9a3b5be3036180a0720e1528e35fd6c9f050bb083af15a215b399f9f9182565ca178ebe6e643827f03d5c3c399289172af79c8a4707d268be9f98aa8964ca62976da1242abe8a7a141dbec1858ecc3ee6d7fb581dbc9439a3503bc584d1f94023e103753a5bb52b47b7dd40d2176f1239e148796c33ceb515cc25c63fea2885719b8eb962ba04d66fb80a45696bcfe6f6cf0c7ea749ceb71c9b1bfd1e4eb15f349bcd74330ae20c177c48dbfd4114817c03434a1965d28fc07f3445a7c511c5253246db8fab6e9df76cfed714347760aa3df9e925862f24f7366c05c87a371a16860b0acee9fdce6ab96004435430fcba938ad74a1dbe939e306f3c173522f6f47a25d08933febab85b324b55c9196610ec7b7a79a980e24ac4703d150f771f4c54355f2582c79652ac8e85c084b1c27643b2434c5b19d05ade2d8f6f1d0d42c143292885ab596214d67bfec8e1b5658eee602d05e71d4226048b333bc62979188904da0a3da2709ee327a0e18b9fda5de09fd7fd2e64e894144ff651caafa94d3a56a7ca284235b1a3f85eb2e21b29777432dfd420b004e7002ba1f0553acefb0d2b708815965179a453675d82c9683fd084ab9e57a53596281e793bc6a8d8375ffdf4e61f6b609fd747ed1a820ac4849993adc953aaacea3dcf622aa3f48c4dc5d12dc28075340c34313309b20fb145a4dc7d869f4d6c38933d8ec37f7beed2030d7b6a19d937c2154b8bc6127e1a9a36640a164dde3f8ade366da9af546898f6df7262484b10857e180b44ce00aaea0aadeda91e5a4a9ab404ffd9fe6e6be0db929e5af2d433844f85e7b46c6a60103710cf3fc7ee384d30d81ec34b9f71e9b8092f2819d1a25aeafb06f995c2da7600aeed50cff6180fafbee7cca18d800304fdc54176d12eb07fce6c64e931902eb9f564cd60e094840db7679efa46ea3ac1be88e4fa19ff435561f8d7ee73215e3659a52b0a950e3e4b1b042aec17bbf8a79e96ceebd2bc9cdf7ab8198d85941373f768198a7bdcd938ec1ac3aaff8c135f361fde022bc543148dff4e1ab25a21f14e54ad1e7f12c1e15731acf8a3f85bad2255b0d9b648641805f2d5bafef377d426074eaa55fe3a07bf95d1e4b03823675b6a2c597e6e41710865b388dc75e9a8637ce9226190f61ba3eb63b9675c1d587723c3911a6625ea3b96f711c8da0a0c7f7c198765a82e99879b5df7df4e558475eea91941383082a713789255f3420d05307ed69c12f5da5d5778db2284a717adba5974f0546059006966511240964dcba3c79960ff939ca4229071646070abb4f7eb58c9d510da72f14c1557384e2f98c9d1ee35913c3bd3330dccfaba633641dac90c9ae09fbf47e36672d076afb658220ff015547c8bf026afa052ac6b795efa07f3d7f76e912fca7316d55869cfb1dc865bc7d0fa0e91aa76388bc14c1f8e9e70895a7db44c2a2c0809b7ac8f073b3249f4daf585ad99487a19f194feb7b0236baac81af7f4fe3c31828582150cdfaba0359e2363c1e35b6ae01071a5c7cfdd57cf80730d498739efe97c9bf3c7151be581d575440775f0b602cc8532efe8d27c503abe05d9aceafd426d23cf64a620e472509ff19a1152835fd63bfc276a11a79ae654afbaf2e1d6106175e88783c971a579ed6bcc21682e626bba07d94875a8338dbfca5c60940834add5706edb426b331855f68a4685c7b743c315867948f114366fc551a86c2c8b3e5e0babe169e4d424dd8bceffcf9cd6fb50bec647fed23a29262297388b62993379cc2a248b34ca4cc750f18b051dca6d9c58da7646001f35334f0a56e36877162fb4931d6ac8f54b5130762b439fde3732849b71c6e42a7291253f69a97c9250de02b312a55dd4bd9cf4d5472322f8a8e17d52d950c7ea4162dedab3c75e8c60ac553b7861eeb925b078dd932e14143fce84b88eca94155ec030e40c8d07c748c8fb677dd019d12e3d3af40ac4f7fd93fe5d75fc3890413bc5216704ebb683a86c63a5c460cafe752522c41238e4662c54725157c3e9d285ca43bc0450a70082448f732cc669d8867ead260bd5b0b509c091664871875366d32742305d6e4c14bcab76736d053a1210567a5ec0da20af1c90f8ca2b18cc0a8ee582b01005cd7e035909e0ea326f73bf7ade224612226d4229eeeb40ce0522f798d01fa1d048f8eb748b53ba9be9c94146de0ad0e06d361b9e81b53f747d0cebbe0f073bc073201d2b2035724d0473e65ccc958a149aa1a18cc7809cf375b83bc8f2d2a1b61b4674b090e8dd1ec1a38e5ec98871c3456be1993d422e45ed8f2858be8f0429242160c04a28b24f1effa54e7d1cfd89559c7f16c374ad6ddf19311f2eb52cbfba4d78f05c2ceef7bbc52641e140006880fd309f3a8f399b52c69f55449ff954ce73c0bef2acb7c429ac7c8b88af051514069d5db88e8032c272c11a3a99e35b729c5166b22535a0afb5cc9f964fd8c683699ccb59d4ef55a18ad8b764c1dbe38c4fa26299f385991002a928d61b361c758639c98a027ac467deb8f566c98ce4094a2d9b2a919f032eb52157420ed157804cc0379cb05393f1d16edce5fc727ca8c87c81ff3679eb5f97db3f201c9fbf5a33408f935eaf9cbbf38c75a33c799a18cdf45b2383546db916b420c98bcfb35e38a88309cc63a46c6e0cbf7075e29cda8172c6218583c255c7a4f0b1b463d3b36d29712bce692b2de69caebe230df5c825e85cfcf7f39421deb6338dad661ac56a3696f54473e1e68acb0bcb19d558daaa21c9b07f32e0fcaca74e38ca8a041c0cd990abd0f3004e3198dc2cb47aaaf38452efb8ba01a198bceba2c30fa5332fa249c706c740d9f85e1cb9391ad9c4cb3796906efb4c9bf9609c50742841d13a6b7c0be702822ae1d9229eacf41bd958db433440050f7d6c8180312bfc0cd72d8b5e492fcf72d30a59080d006f40b4fdbf6d0c63c762961a87caf38825f63ba8abd35aaf43f65179d8eaa9cc5141328480097ff0536c8ac74268706b703772fddcdae97df405311260f69a6c4b152182e4b26744d9da09cdbe5394e2d31b4f54731cb77994b7a89afbdf9895acfb5f2682c5f02ab2ede6ecf3f7034e3f1b881dad490f24b751bfb00046417e9ef6bbe3dd617a9cbada2e97846a675fce847af111d1237285a46d615c6db6ec901b75990de39d7670ada7370e9b154a16e4b018cb4860ae377d0e1f68f92a6b3190fb4bbf1c933fc00b7a7e61e0f51f9ff0becae415819d73fc794f37cfff3b170c989446da82598cce5752586bdd3d75bf62baef5b3305f49233a0a99de3fc0a2a776f419b40deed4a27abfb45a5efb7492ba12b775361d49aa820b89e9634f5cc178f6d949285858ac9a5948eedad22cefcf75e5e6bb2ed454d0b1cc2498f99db785340830f817d941dad2c091891cb966b36225da714c3615ccfe4f21a02d0025ba9e7f326b668ec08afbd78e921f227e2f581d5f22cec4db14668568f19981a781c1fb4e99b4947cc60fea897f388cddd59854eddc95d024ff5d99bec7041b9e2b2117646ae1e0673eeb8f19cae125c234aac162d51ab90d1b5a1abb67c492ac32ed83f17e77c0d21ee564cf080e32a04a65c1e1e2dc15a9521226b4f5a12031af0aba02b196f51a4f2e28eb1a9e71741fde2b06f13a66ff939138860988ec230df7662fe1cfa5b7c9a6ec818b0b2c98550bdb0730efd285da1fe980761d591fe1f3957204e9dbf05547d0966c405026dc2e4b1894962982b74a0682775a1b38cd40b1b3a1e6842b84a445e7c06a53af414a6bc34d675a36e63ea3db7ab98ba0418539a120314536b22d25c6e9eb3a98e9a9a8095ae858d218294f8d37c541936dadd39f44cc61ea2120c41673b7e53bbd836f6f50600f10f7855d3c7bfccf05ba71f47d0c3e5ca29c59a0036f5e7a35bff602a35176235ac4b54ee884f05ecdb22eb1fab2f3b0d811b51e5fd90c76cd84fa62167324743add08e80e9efd4a1c51fccf1f2c01b3eb1fe31eddc41b7ccb92b413e9f23ab824d5cdc2d43ccee814b8950d544f9f1bade3db2edbecb85fdef52870f8663bd5af3540eb98c00a0563266d6da56b710aa381f3394cbbab86a29048972a0d56f60d8424e3b5f5c42bcd75abd276c67d040f2a66c19243335eda0408ba7788cd68f17ec1d963a7400847ddcda2088ef96687af85c19a34b6864f01d6b37dce26fd0ec4c805f2b8f158b63eb3beef7fc67c8706e644e3795a54d7dc2cd820b135803d0ee17064928d8dbc795e7065ed7d67a44f9abf23e9ae6bbf5cc2b5f8c3b901b1d21ff2f52212759ba05b4d8fcd0d3baefbd8bef5d958dc468561efecc358738b11883c2a735029b3559dd297d5d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h943acfc474bdf1b76bb6c5b5ca2963ee7e290a65251d22a77e9f04ac4ebc0336da8f0fbbbf0389aff25e25c93a0b78374062a15f863a16c0b18e1eedd700f33d1e0ce93b795098131259ef8ac6e06a2146dc0c54d15cc7e7b0a01c01bddb50fbc917677e635bfa857cfa7835d20d1a257569c0f31f09f879c5ccf2b30a3e130c1b1e2fe2513468c0e09cb9eedddf9dce8f4e6bab6765f2db8d2857f54ed6812c92aabd39d93580eef6cbb7176f1eeed653e9c1517d2e29118320a31ee7ff68bf1ef89a935c37b472f4559dfe585d1750225c780d61507ac8ea4a177e30a77116c2c0f8d7fb75a5f48c9aec952e452642d522ab7a29b6c7608bfd7ba3a68c7cae847053fc1150cf676d6661b5b088343553d82327e450e028c112ffe99d935078dfee8010a0ac130456b1486892e3f0b81d78ab413d3c300eaf287896be837fbf7ba92ec5da53636dcb9b6eff5d6fd0764d7068c729a96263c898ebf6fdc68742ccc0995aa793a348ba2a579c3914c584ca563a7523cb98c19065294846db6f6101da5e3b558e6e3db0f96fc5fdbc14296b92dc516f49e154a110c5aca8c99c9166bf71d1414994f5e7895e43b206c7245144a9ad179433518e92f95c8b0fcf528b73a2eff320c155f83ed99496274445e9fc3f47cf5b3a98f3f4d08d82ab1bd0d0601f92ec4cd6f63a57495f12fb4a41775c9e9932f11997a0359317b8a89212dbad3fdf37688bcbcd3e75500e182c1acc6b25774dcb41017e58ec1b33aad9f3dc9a3a460fd33da98e700af4edf44a571ce941f7b5aa1b613787064822a648174d0e21e8dca78f161ccbe6009e8809e73eec5e7251eb516b5dccd17f902a2b49813ad5b4c296b3469c912be6c8e5e79efdcfe82f58534c6a41b29a374696f137c9c0c6ea67bc7ae71a94488be4786a725029adef46cc1871f4bd4aa94687d52660c78befb54bd3a9e1d34d305cd69f610afaadeb2dd7b68972f1a8a2d3587b3f7128ebcb729cea25ad5797a5ae70ae57408b4674102445c80b9d7ff92234ff66311d2afcb8db719bfb75f278422ae74d5528a287a75817fe2b7d9efbff8a1ed368da70abf252057fc43f6015b8238c5341cdb130a5dbbe60b98a4e1b3dca876b1f661fd2683ad634e459fff2782319211edaa2f7e617d19e2e2b7f977aa280b745da40cc27eaa61a2bc5d667d2572f6cd73a573489b27ce5c0acdada4dbbfefd59d063dee97c481f718caf356d32fb61aff73b44ca7a609170a3731e6f4b25b05eda1fff18970175fe1847460233c8ebdc825a7ad79d509ce5a1f3583aa4efe6af56759ad1d68fdd3c80f721c17bd33c0f6a020b067007a2fafa149ed3d5c0a870065b2ddb26d801f93e08eaa28fb4eb2ad2e2f957c8d9d018bd991d4e731b8b7a63d686c0802b7e14235ef2ac48e34fb5e2874d0d6d95b644255c358bf8c69d0ce505df8d24484b0cb6dd422bd00cdc6bbbdc0d5478348b6177ca8935cf0a8d278084d370ccf6b4f413228044f7c309761358284be4fe9c4036c00c1ac4cd337c2d9a585c5b0536741fd55a73217c4aebeb967354fb6ad2b97055410ae2a6cf47ad0697c8e044441a8b796f97c6da0d948fa249c546cd87e03b02a4a5c7f66bef4b0b795478b3f9199a2144b791270c1873631df0b8c13b7049f62403c81c3734e89380b498ca02928d9529595d1767825ab2501d28151d5d94b963242827ad7aa3824a5f43b3c4a6ab9cd3a1ef2c07158f1275e46a83e20a8c0ceca7f2b6693baccf4df63448d026ee69d690f18f9d1073dc9036cea6cbc99ab8732e1f51e3d30d20b587644784705a090b845f2a33eb8456481fedb4fe477b36639427ac28cbdffecf534e48cd77f67b0361675398062a6afa1484757a8e5d85695d5d5f837dc8fa9c84d7595011a4d015aa11fda68b3a837506fa23e7821d1d879ae910f758cd0643c92cc6ca5ece5176198ed56a1c7312ca5540cba4a669382f942618a4536c6ce371325871c310338a0c6fbebf71e2a14203a5f237930e87bc68c108a358e37d75f77dec1291829b1329b9711297a04034b63cdadb199b339b8e13c8f0c33e77c0a0d7e57933dde4286f61b30a768dccdc3bedf6b56ec493eaac1a178ab1f1f76e0d19cedf095025a2c7d37e8e09af75d3d125ff0723c175286408f45f8f0b7e9b843e51048674b1b90617ae70d7659b651c66006399950ed7633635102de4923e731a2f4f84fad4c98aede167bda649b9b0ef7f25eefc47a089d14877b11759a62d834ec890c05a064defd994cee0185d9dab89dcbd82d354283d12a273fd7b5f3558f66d63058e6d30b7dc603764f43b9500dd94cb11f512e19b1d5a7c3f3900716b296218e3aaced892a7670e533296f2d58ac8d1676aecd3eae8c9380ded59fcef7a83972628651e9ac65ce8885363ef2974fdd4d6989c2ed5972fec2bccc4e71cb56d9da45cc7529d611620798394a10e9f178fcfde7a81700e9614b359b8f3005cee4c9dd50a2a45a5fda92ce87f78b39b6fafabe2f6fccd743b102686154b536456b26b48ade7911d3a0954a941c827f2f7f6f159f1eacd6b2a147c217c91642fc4b1fd5eca1146965b1c744789e5d6399dfd745b4312667001e7872c95994870b69942631a3893c0f46b2a5dde35d120e101e59c451fc49df8cc90b7fb62785c08f2bce272983c4ac6faf9cb50f2992fc1e32a90c1b361853a96fc4e9bb045b7b73e0f52b5a2d5ee7b8a8bd2ff63cd35dd79588f2e46223380458cffe740eb789ea3cb5fe97d96b3f095bd02d9607987f9626835979ff87b382a227df070a479c8a9b41092d1e9d2810dfdfd0b05c2b4c72f107993dcacf87f05377ea3ce03bcbbd95741c3ec2b663d2de83eec2028b62c0fc823f22c8afd7d79441a78c1566b5f8df11665fa1aa51f2c32e045e0d38cf74320edbb8b62790c9d6926e8003e65aa5e3739530d8f089eb05829a37a41054aa1b556e25a9e91450f1ddec7fbaa584abf73c99a6f17a7e921110dcc8847d9b50aad609987affb79cf604a0fb5760dd29acea217c0df229876db8767642db0b6bee3ee78bd041f62ad9b0b255cfb39a439d435cee7429b0e99f9548bf76b49d59123246f3e13a3311046f9702df3ebe9e3525924c5fc00fb8cac360bd29e25088243e33650f673f6e709fe5039d5b4811e6702914d8a54497cc28ba944363e6b4d5b06791fe656204ea9b1dfada3b10b3b37c214b3afe162f402039a81aec511cdf75d80c837a7c7ce93580bb9f184c7a142cf0dd070d9773854c06cea9d25ce6be6840d88b99988f4bfb931309524be903536cb9c2c5b75a3bf943f1c87df35203e1325ece091b37e0fe33007fd56435029e796b5ac96a2f942313dca5aad829d8cbef2948a50409e47e773f29b4ab2b71ba3c725ed60c32c65dde95d4f3540b4234fb352b1dfc0b0e868353aa4a9a919bcb0cbdb4d92383a11830c2ca497c5d2e2bf55a9f726cea60243ac0703cb7aadb20da67b6adb9d81d7d3c739b1b07cebaf94440fee6f20b4da8fa10eb5d4ebebf63f467ed83564843ce1d07c861e742445402106b7cfd88aa9d7d6f0af01f894c1ee88a134b879fbfddf2860a0813640a6cb0b2a761f7d2289bd24a1185c3a1031a6dbe6ad81d1a650f449a7e28c169aa1fed47ab946e309c793ae3f5d0e1be57e646b010cb9d75d253cf3dce3a4bce3594f0e2393bc6c6d210515c7a5295107ac18313344115cc46e4c79412677ab1ca4e7810e28b74501440e5c1f9d69745cc32e03c135c60cd1fbdb6c4452a3eb7bfad656cfbe802324aee4c7b8db1338da2498bce5f5f9a73a39665d3b042960b3fdb808171112e12822f10f6fefffa3e8c38ed16e61d25add7a0d01a7a1ed1f81750c91d2fecc2e94614b7c156573ab72843af0861067ac48c17c2f4df84bed537b0b73b7dd1bc0eda662a83143e365ae9cddab1afdbbcf219d6c2173efba6bb180e73ecb3a89681826e8d754a0da788b72b10bde9896280ee57b6675062ec98ba8abc43a0b2507fd27d81aac20864607eb31419b8203e827aea372a96ef443292c175ef4751ddcc5926d0b03a07886ddf3369996c949891c16d0f89368d6a4691400ecaef934528896cd19b240f9e51e6c462d8bbc832d4b008d6739c031d888aa38f032e750884d6289149a280c9c7c6c6e0291dab31dbe722761c97072be0087a34c228899b7302a2cfe46611965f4c9aa34f113228223cc4154daf96b7142a07f57ff46a5e252eac9ec0c2448191b1c1f93a2e9b855b57e6523376a09db412eae1e5b2ee2f32f26bdcbc281b459c418eb292b0d683071af9df12c35e7c7eff0e92db5a483095a6484195cb73ec64504246ecfbf4b763d54d340a88d4f1ab6144d6e78a3eb28647e493b7796796f1700cdac6a898c32c5769c1331cecb415a01267eef206697a45061eea9f4e8d509b42fd1f3804f836c913baf613378c0b1ca3e13c70693c54be2ea3c8f5235e117ef26ec24a6b217f64f362c65202bb6149e3d186b43691f232f51057efa79b3b0bdc743f2e6da4facb1e5fd10e8ca63ea775881fa332160dbd5b16b0bb9f89ee196c9477af74ade6cbbeb7390517ead48154a8bbd08616cdd9e4f3486946f7809f311a0359de4158fd483eca73e234d7b4d24b9b1ce8d824adfa34111d42741323cba9c72b0349b8eac4d01203aa973ca4eabe2e293982007eb403d53f401791305b8218067eb6a5369eaf3ee3016216362f525157972d2107677e6e57da7e74092f3c7b203c9f1eb8c6ad629a089006cc07e1b5cd73e892eb313a5fee616d6c6af43ff7e28258d8c69dab84647bbcb46adcc5f1aa55fa2a5ce84990ab6f96c5d5761adec477b90d7173a42b9a774f2cb3aa072da37dd7502258b31a29e2e46c6d441dc5e5cb39eb29ba74f2c3c7f5407d5666140090a2db1d74115cb4fd97b1d51f6ebadd47fdb007cd11f198b31d730f8cc87d6cafe70fd36b161a5570e5617b218de73d9bea14b6d1df9db59323692f8a4f5f90edf8e25d04105c357d313bc200b69c59869b23341a3ea11a6ecba16ba7d473d530396a19ec35d3bc01f2429451d69c185cdc8243d681856d1df7992ebe278b482723729a9042c5799fdb1c85575ed8d0d133a470cf82e0fba602f9b9f71600c26047e358e3c3fcb4374125b2e81eeb32163f0c7f288a1c0de5f02cd50cce38619c8890b96b555d1e930dacc9d944aa7cc233a641a37bba79879383167fc1a6416921834c9d60af750f96efd59da584a55099d97cb082d31809161a2b8afcc8fcc6ff24210240e62d75b151ad4337778f687f1de759aeb282948958f28bb743d10a986ca95d0672cb7b81aeb3aafc88cd4d81e30b593777fbeda2de74bb970c3881008b2da844bb08370912f6c9b06ac32097a7af3382efa0a0c9648db321cead25d2db9f46c963eec809c04ee6fb39e7cc6c9935c6f1d1a2cc8df313a0a756aeabb5b137468f8bd6f5325fd20d732a6c53108c54d806482f83f3032c949d3dbafcf4d1add52be2b6bf287c4d544869bbeb356bc0002010267f7d01f68d670f758a0b0c52c7271de1b79dabf6cbdf693b00ad0165312c8d27c319c4228c9dbb003170dfc0c7952c753f6d0b1688ddc01b7d1d6bf78f6076ae24e3505ff6de47d57d0013a24d1da0f0d0a9b49b36bfdccaef99008a8bebb693014efc3a4fe9a51083635cc4ea887934f96d1ac927b953e6ca396ffaeb7c6b9e6817a7c3df9b395fffe6ca15513a2fe44cbde8522082f894ebd45bf70a65c2f98e7470d9107864eed7f4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h59077467aeded1ed0c29ef6b4ea09c892845f41af6aee71042166d2224a8182f65fb23cc1320de4c177f2e722388666fe2b2615cc8b9c1825a93917a2054af4c74684c0eab0cc68ebedfc32a2cde224bb08434ef62b6d834e85cc84caa96eb9be15d772d59dde7081df3d9bdac249bb2e23948ec7537ddae58f1b9396265316d5f13af8e49d090a8d148b1ef4b855e1f4052a48e97172cfa6bf59445ec89fcc50fc64c033076b72fe686de185709e9ef1079c97a3007c62f1b7d7ee5c2468fd7f8808edd5cdc4335e70f42b616ca0353396c8a551ca37134b70426d46a4b1e0cc077f394a41449b0052ab6e29e4594304e86ce01cf9424b9781de952a5a6ded8655389044974e0ccd3285c782b3a76803a0a82f9ced5c0438e070b655851280dfb3e2aa2bb0628d29a4bdf5e737348f4f82c4755b3f238f2ce78841dc6b5e508ecc8e1126840adad5024d1f81f351da1bff7341dde878c2c5b38bff14b366622f447ac605ebdbc6ae8bbd66d90c1647dc50c9f89099a8fac040a07c48c525b044bbb2f8fb3ec255cd47f6a6378b14f4b24cfda86307723d84f57e7ae34227c59a03c3444780c835d1fef8a9c85b6c18ebb9ed43e5c20ecd90683ce7575ac0ceec579eb0ac9e8bcc6a3243ccf32d2ec2fd7a9eaa8869cd9a7f4efe3c66a78246df3a7c459c145b1d52e30f984c6c4bb6db5da1291360d7dd413c00073c7c39bad26426bc198b120b256331c3f6691220e53a1896c479c49225b93835659caed680ec6e843c1aeec0958116c5aed9f88330d575b00d83612fe6e1b61d490e744569df081fe6a7537045dfdc85d703e5a52006f13730b2969cc94cebb47e9e0b6233027d18e07aba8ea68b54e9780425ef3949eefd959105bd6cf1105919ef313628c5c4060ec6859248557bfd788460dee6cca441e16cfa3499c46c91d9bc90c8a75faf0d22bd5abc3079c055bf5bfa13567dc3a81a869c0e6607a74167fc1cf86ef4280c88cc9ca063877eac2f51c0c3e66fb515f5bfa1c44c13339997094a7e7a055134b08fcde6b49a90c92d74d5edd9d46dbf04dbb2e6da7afa9c2318ae8003d73da0228012379abbe9b3375ca478cf4842b7685e2ac9f681450662859f0496d0233b0095f57ac2418d443b7cbb3573d93d864799b4e08f7a9c27503457c1ffe9c1a774741b0b24452eb946824d07dede7cb9e39d1450af8fa62dd4feeaf93bae8fe1cbde73f40ba24f3e0e198c555dc08017ec8f85325d20549c1302490462c0caad515611386a9f029d05fd65f3a17a4603d2bba1dccd8c2b6026a1f926e5f730a11f27fc02b58040a3d3010bc8d3e55f97878d7ebc8e7913ad7ed1c11a55b61867e4d96275b73dfc1ba4cf512b7b9e8bc98f88b48a8ecec98ff9c46d59d47c721f38c12d644ce1804297694f00f36cd2a68442dd29f52754d519263932c5ae23e4d948bc09a9e52132ab8400be18b8342deed9910a2569b188bc037acd5e3d9616fecb1ab4bb9cca42e5ae28e3a9fe88e69c7ec2dfaaac3aebb6ba922606ed8ccc6d88bda8268652626ede25a9c81849f3c282d55bcc72cbd5157fa0ef7d9d99a2e0e1be0df3ee923cc025e7a04cc6b17518614f38993e6232bbbd1d49396f32d7d7df83e90ce23d41fae43c7ee2c5b74c8cc371e6e00f89581ef98df1ef7415fa88975e71a4181c3b7b96340524864579b6ba5f58e8556021028ab8fc715ddcbec63ee3578dcab1ba5d6aaac09b1fd7c1266b816c18f1f64b0c0131e33f794bc91a9b04d903d6df8c0541348150b6f16c618b663168fff0ec6b6bca7be36a1ce64ed585b315de672005ed83c306fdbe67e27bd606f269c830b63f8c6b1d8325abc7c6b50cd93c7c5b4264062080a6c8af9ff2ebb55a727a18c986ad3414198c5c74e8fc5916aaa7b975e1a64b242eca3c9fb6fa0e9533870ea907d2a447513b492395bdfe3caf72ed190a290d4e8576b73e4acb2edd2eba0c5a54c09db8b52ed202ec80f99d082f5bbc1ef02f7d7e3a3a8510708a551d7b17a7f1f3f4fd34c0da9e8d24a4061eb8be46728bfca406e6cdd3ff1748520bb404e46636e09b7190e1d49939e2ebd5281c7a792f73a5b3fb8a4f171bd71a9d27354ada6be8801ef487b4a5e1ae13ea4d8e5e2935da1a98f62b05a1230f30791e2861483569d7ef9a9cccae2113feb3367d205b4d6f306923685f623050872cca7cd7b7d76028035e248489820e36e37dbe409c867deb0dea90df4d843742b48c99427356df18a7c985bde86545160c6ccf202d0718adfa376fa445f5177e77806c8421bff19781c64755d1bb44d659af0f15276ac99a1944af7c79a51a2e5f3b7b022128c418c56589e90c0a0b9671ed72cbb20a0092bf82f511d840037a08bf6aa65544e706cd3c0173178536638b0b1c39182f28fcd88605133a895fd94e526dee0a38e5b790e1da6c0717b51185e1d7b73bed7d4d453fbd168ddc769d66f21c4f57e5a93233a3e8d5e3b8c649e142ae282510c762ab7fd8d8fbbe5503bbe91a5f850decee31e07f8d4a28f5a12640d8d51feb70b1288716a493cf342851256c12883e61ac10186f062358e7acd224e97b9a83fa894b16ab2d3812757ace504585015b1a0c8d87a0c59a721fabf43d667a792e468816085baf717822ca141b466cbf5143845cb43d8a07c11a8fa9ddcdb16e1c8a8fb65653def411b39c63398b7e91a741164af5d2bb1817895ac8d913b6de54e64f1592dc9196448ad57c1068c366950a4032769052255509b684abbe552b22b2864f298a3268aaa948c4d3c40c58c29ad6a60bfde4fc8ceb3681b6de3531c99088489b5713e2def0bdd423339bb785418f464ae68f3bf16d77b6a51f1560a52a9461bd857aeda106308a5d0f6cad8804954051cdd8a6557e70492d8ffc04fe378d72eb1cc344a5a79fe639d50c1199834c795ed9151f23fdce63653c2aed5118b19552d0bde9e05974ee62ff8da71c8028ee61d64c0ab4f0199f333a2f0ba0aef5c5fad75b03ddc1b71be0f5742184317aa092b572de0f62c6e7964d67992043a5592f1e90b5d31fd27ff3a9dacda024048ed0ef41d20f8c190101b149ca6f3d80cbafa695b1bc311657b18a89812da4f42a956e2d38337d3e8d17336b7c44453304bbaa08d2507bf411a35a541378871faa551a6dca127c586c98f6ca8db1e1174149549fa3bb87a143e5a89598272634870d9821d5b1fb6095e59c83da1d43edc6fdc2e59d45681b741cb9f48b19345b06112a328365c29a11cffe91445fe3384a34aad49506a35b939b60f659603520e69de869bc00054ad8f7e2ce1b5e17b1d7e276022cf8aae46359f2c45237c3156faf3802c5fac1ded2f99e013aa18ac58cffe13e78ccc56d71f2c90078c22252204e0d3cd202a5b32de2d8c8424f318bfca43564463b0d8c8a185f58ae8e521b3b6e33d53375eeaddad173752a3078e512db2c00a33e71183adffe220ebac9687209274be4cd41ad07eb9bc166a08c469aad2167e0f47b0eae18f2e881e1e54a508ff4d19d533f3e1e5d6cd5f8218a5d71aaa39a811bb22b1808f12ed5994a11b52b7066305f4e064af1b4422899f95ac69841dd9ccd221b091ab9e277432609622f3d6f73b9a6144cedfd176f78bb8725de62027169c72dff9cbdc4ee386998ec24d6ae98fb2da30f64ec083041effd72e9475946889e1e0c32b36d83d3679c6d516711c4ba2613deedf5c20e81a3fb48e2e6fbd4249eeea801bd49e1df9e6c9bc362d9e5e0bf46eb6c9602cdb0aea8743227f5a10c6a3378bf291d0590f24fd0f327cdf85dff7c003df77264cd78e34529a8f51b4efe6e58fe321907d4c2b9e4337fe4a5879dec306c8b56e08178d81a165c01db6f208cbbf53b00bbdb321a2c5f92f3b0db772f1659e3aa63198180477a801a953d29374cb0cae5cef63e66c048d23541613d21be201a3394ea7265728d2f3c93d064fade4923e7f169bc3de1f28272e670424579e3450482e2aa5c59a3d156097c6a345e76791421a8b55d77af1fc490778303cbfc6554c6d623f78d7e3ab5840fa52d3e0e72a38a723f4ec8578fe1d4bf1388495dd3266d39b533f5a783c1ee2bb72f09b0c8f191eba605c2f66e1ec1e51742b00798c06ee9c3e97040921217d3b82c8706bed19e73438e7d5ebfbbd870b09e0b869c259c24ed099eb34c511d73177ef570679c7e582f321674b9dc606089c187f7b4afa5188d8cafe0d6b18ebcc79e8e02fb4f896c61ecd1cbbc8f1bec540f659215d490560d8aa4ed2ed2cb50220bf327e45109a6dc24b06901b8c12824aa839ec6652abf8b079063890d729c17b90734165e0a89013ab60bcae882576044140d7aada1b329432092b9d2c772598fd0a1a6c56bc85b8d34cc76678a2b23390631e9bd0e9c53db0445843731786f3ad475bc2a379288d26995b0a6bdf54f367c13173108a1ac00eb992c33b65feca211d4de4549266b69d89046935b602102e01ceaba1d8ece27bc1e59315e0e28833da341df480e8fe29101b9a791c0fab4752e60aeaeb0ec739a027f87598f148dedc421d6e0947368db79c6043a9360000bc6ab84e6fe0c1ee823e312b6dc0090f633c58b2dfe39a6303b0fe1da8836d0885784c2af2fad983912e7fc5f5a3d84a614aeb8c0c272ec6f6f4ac848198165d1b6fc253d22593bde4836f9420fdbf5c507ad195ef93ada175b70035749860a20d3fd541b995b96a993a4e0eac67aa5a5bff096e17a38c4cbe270e514b13efd81768e41bf709304fd88f3f01fedf899d5bd661b201e8d7ada0ff444529f5892ce23fac9e11ded9bdb29d5b6a8d153a784dc6fe293c99d072e3506d178011f64a44a652c62bbc09f0a904258258e957596f61f1ed0bc805e716a1ef61171e1e0b96e28eb2dde7f95af47e7cce5497e19ee6f6d8916bccff056c9f81f0a45024647de2afdc650f93a3f6d4c68f3080beb5949e3d37d17d37b0f404e11d12b9516e1d1c8e6f4702c259d7f9f734ed67efa0b79a602b3e5f74413da8ac5785cf24a29b7604e082e0082a4cd88f5c08ef96caee47e44af1ffd18541c02491bcc583c91f934ef023ac3edc320f12a9f6a62a6076925953f252095edba9b51af00afab23c5704d463a8f15bd4124648dd3cfdb7fad28656c06bf7db451403ad18d12c47463ebd082a66414c1001b877bffa5032db22d8207afa136ca95e99107ac7421b9469f29f57496c98d93fc33b57bf1a1b33952b58a1bc1d6c0036d16010d9a045407cf402219ce2df8ff384b71dfa8187bd1b028de45cbf107290edece583da0e2e2c6d1d67f59c7f717f27fabf2bcf39ede5f8ab21de207f326e1e73c5d72c50663078cdf710e82a409d81605673b9e76cbd52f0ea241e6c466b4934f4d6c92bd90e13aea8519704b7c78e8d51ba042896bc2fb8120c1be97cfc22026ce59bfd7ed4ba62ae245ab1914c2feb15605ee1b530f6cb04574030af9a38d10e15f2d504a327b6f465b05e6384e3938218c413d7c8b940bfc8901a1b10484e2cf96c73a663e1049a997af89145d412f1286b1e86af2fe68f91fa3e866437b92d6ddfeb9a4aa41ee37c540681f82e1a54d152ef93bb11563910268d75e21b8619d6584c8395b31608544ac40418ffa8817ad467cbaa467eb0d91c260e12a600b665350e397e3ec5c76760f21cafdae9eda9f18ceca5f9d0912e0db8204f037fa36dee8807433cfdc8727b6dfc56959ac2d4df74cace5ce6353cbbf67e927f3d2f65ffdcfaced88d3db89dcd1daadd381f2306e1fda56f37fe04ee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h97d190514106f30718156fec58c4598bba6f4dc190a69e193554fe7116396890972311ba7334412deef53ead05655468070982f08e628871988331578dbe602f9a62b6c6da7abd133498dbf1e47589d56455f43a7f7137a6fac6ebecc2edcc2c05a74a22d56b50d211e85a9a8697f7f5327a3a44d09134923968f90078e1cb1e24836eb5fbf91fdc6d38d686d3be1cc4c45de4f71fe46d5c049184ef1f75f6a3f4d8e1df97417b5be67d365da0cac8e2aa022f2fb49220ef878a42823a13ee6756c67515fe9ebeb9c2e70aaac2b4081325b29c97f35f83637140c0b7f08bef8322d9f974b4fa9f8b8641912faa3ddcc092ddc3eaa19c4086b370ce32bb2622a13939664f315cafdc1bebc38878fa69a6e939b762d8a7949062b0b6a8e17f843c932292459487c048eb08a8d942078dbcedf9d5b98215e4621032b6ca176355fbbcfb900fc3dcdd398cdabdc63a29667932a6761519c6aa8fe70ed1bd5d8d7969b3378a6bd0e30600560af7c3d843b91b9c942a3ec0b382f82530b00f44c25dce01dd403b850d124c1b5a17715e9f3579171fd511f2d26f9a357456718e2d0e209daf18a73b6281b131e0dd6501f47a06b9b6ba68d63144d73d969d441d9533e2a1386464b02d2b8cda602e2298340143e730a3ee45ef21d0a0b7cc458ab7d07a8634f80503445686762bf3d68a63f850f7a6399f0327b4ba1a257749e0e8a3ddc5cbf331b8fc59943b3094ad0b9732489f03c0d7e85cb6a6e27a0b2ed937e5c1af1320b39631432cb2f3c0fa09d63d3ddd9ddaaf3eae4194484124637ad5da1a490159d8472eb337e71c1a8d10fc6e348fb6fd695750223720b35da7d687d1ced95942f30671ca4bf9b2fce2f28ebb4aefcf06f536fe888d4d87cdb9e9be50f3885aec37d8f6c5162ef015996199392a86dd36bf34a324baa38788cbdcbb162b9dcb782973c6c67b73295cd816418ff4de329652fdc0b6652be3cb3673a4098703a784e660565bc9b7623aa9e7dd4dec65b5dc4a6bc36108a9fb8f08c2e23dbaf707a79e50759a80d6891627b46e5f6dc8010c435266dfbbd54a905b178dcaf8e6eec6513834405d8c5427f35edd1ec74d0d9240db1a7acaf793a90eb8beca30cf727fa307685f1bfd527becdbf5095178782d827f74e9401c9e6095b7f197b1ce3dc9273ed00f0e3603220a578d31e21259a3dfa20a338d3e014ef5e58582246449d1cc2a44f27095c2ee6345b9397f20e9fe0ef829c1813ea8f5feb26f6fb29fb7dc01131755c9b53a16782bfeeb544623ff0cba2ad496ffadc27f7d0448f7c8cc823c0cd9585dd740ea2550f9561cbb0c27b1d1ccd58d84480e35f722c0b5e2cda33db4a44bd0ee24985808665d0ff4f4f04e7ab313fc45bbcca057d7acdbead178e719606fc50b57bed296cc417291e3fb82745c9eca901736e72d2da9cca6d8b5e2d3aafb454afad22983370ba9c31cc2a0643935169d5a27f9b2b2309d845d8a66e431b6a5839e1af6f6f5827aa29e00686fb932406a8c98dc411de12f53d345b2a8d7183fdfe13c56f4abc22cea65309341eefe6e6c112f94c74e9c35247259881c0a699c496301ea649f7d55c3da4deeed2cf91f2603411cc1ce64a647bc43d1d72222ff087152f92a9d3c3a6f89d66f264e7530d920e0caa3c5473b1671a9d853c9525ff6e7c55fa290e9d2a39db98b1682fb1ae80bdeed6dde887e90e17e4938f32efc406c17073ab3e931192195f680973ea0fc8393c84a6491cd6c6a3afeb27242662b54fec3318f3301f4b2e0a81e73ce426ae8b4211b28d54172a09ab5eda1e6626f3d0f254717d3edf80b4fa235f8f96790637d6913510800277cb613f92cf1c263fbc850e145c0d9b9258d83b59b2c06ba00e2b43523fe06dc7f53738e1a143c1a5a3094128fd9769534bf5493a486705d9e8174fda174e74d42537bf4472a42b433f28a4bb1dc99c9a4fcdce9aeb8eff26355aff568bb497ddb13f0e9a2a06f5ec49d8987f8f1f2fc7887974a957e43d60268d4218de7549670e59dd8a6483fb040e70f2b04c4d8fbfbd29ca5d9257cbcca8c7dfc413768f8d849fc120f1abb89bceb94445b4314918be3776a2d107e3f73ae527d21be03739dcbf0ef2a416182b4ba7f9fdafb489d8e1a66e2e9bb442dbb3d202625d3b7f3afb802ba0d15002186b81548855d1e09456334d9db1773501b82cf68e2230d67e3f59b68a1b6172520907af4764a1ace19ba1527749d30500d1ecb0f10e01b36fb50ff4fd418aa28584a086e9c7cdc2eae797b67bb6e09f3297608fe910e4f2124fe1fcf916fb2cb4b5c4d07069d208a452816d381c340167ae1687738805d59d35cd1875d187ab9384c9ff9360b9984eb6433bf240380769823ba5b804909113db8991f849229d033acc8bb69b146f6df2af428aa5aaf782fad1a40545abfe193994d1bf1696697a64a4018436cb311f55164fc986b42fc056514b73e2ace6a5ded1f6f17116d033e462bc7635c4849a5d323f510ecbb514a01ec4cd07b2477b444cb94b7d5cf81c39baf43aafc85b76615509b7c3def30d377be7ef0ec0780d6afef81c1ca125ec6b25c06beef3dd43d953861d6e1b3c53215bf29ab6f624f676f37c423626a57dde445c6d511fe108beb1e2fa6fb9fe8bcdb83dfeaf13621cc941c7c4edebb84bf820f98e3a2d595fd6409288f920c269544a81a20cbf198f59037aae7aa0d571c9e4d1de28b057e77d2add52a705e593519d922c6f14db2215be4141b65305d4da239a57cd89c80c5e10bd6a30a90a1eb3e625ef69e14d3170a78813340930832ec37d6cc032b90867b859241397e404e383a1ccb660efe209ff0fd503f9b1bef68286547b02eb09d7df0bf9585fa6ef5701f26384e5418beeb960972494c977be3918dd017c174b623479a4e378094ec2df04e4ca6a5640a6d6471a47ca8b0b0687b663dc0f3b088ba393c1a7576ecf3938062a1816a8403c688139518a225e456cf4b2120fa2c1df60a954a6411f255785d023a30f8c0f05bde3ce8574fd4b71198e924d3196b32ce1e75803318ac770f4001c7fb50c12f9ba78c599b097ce612398b9a341043757cfad523aad8bb69bb55a8d14bb12f6daf91349291a4e20f306c12d518acc1587b7f22ea41973a556b399c1f0bc5223bf5c4263e3f91b7bbe83e2acc4399c0576136c301265f6687ad48a9c10fc6cf0c404632661e9f71f931d01b03f7e03a8c214f46cd175c3f1ba68beb5360c338717a125c38e5b3bb05861e91a54348367188877f89dff1fa028b7ba5e178ec52fa87fdb50663bc72a12edcdb18dc78a2ba56bdbadf150233670097065a9a1cfcb155e5e4ab0b3c19482f6397410c082187579295a1f15b3207154a221737cca3d5967be6a158754042632b71c0175e5c54a36096aa6b7fafc6fe3f666044078aaf457d74079da1565d688cd32bd062285b8202c1d6c55006aa8b9bcf14f836464f58790a7943e335be884298048130826379f8240faa4312a7409b6c04b91dee0ce286db5803aed64a18dd5549f79977fdd1131b02fe4d3a0d0055bd9093c463d140c396fe65f13a8f8b9c964b719e874bc10f8ed729ba4d95c3c62c51dd05b2e138570885b62f42fac8b2b5d004f7654b07139f8efdf17b936c56c21b86819ec44246b1a12f936c4720f46377e9e6ba32965b4bc3710977e2071be7bcd18c24fc0d27db632578f51f8f5c4e4fd131f4636e3144526751f7be2322a0c3a7fe543dda9495f001a41962e806e02ef196710aacd942a4d87d25be75e6967adb4804b707843445a71dfdb76ea3b754c46e877fdf1e2a8ef44212031727706ee468e22eedc2c093dd60a93c67fafd4bd042f11971eb70facd1edd81e4e857a753433d6bb24542fb329de26c033dfadb19fbbd644ba3474fe90005e48973f279cb7b94772f857f4784808fcd6144f0740d0076efb21649265756f8234865d2cc2d6a2e39e4fc574be4b9ee8f28142d1e730548a4718f664af708f85871bcfb71cd542d2c0f2094eb0a170c91b317f5ca734175795edfd8da37a446beb187a7722e0757c2bbae143f74f224e1b6f4b17cf5484a8c4a748a752a56ab59515d5326b9d3accf32e7d92b6fb0a0538f8a5f67715ce95aa338c2a3609e88b94537790625ac3e9ecd09ca3be549d3a98fd18effa9e5c68d33317af820db15ac8ec9a6651c706264a84e7cd57d966baf0694c3eab6a245fe7207c7eda5f4e386405f7ca8f035aaf8f5e955fdfbf09075e57d771c2d871c5c2e77344957ccea9b7b128c75c3401e70b38a2c9ee02d9358fccba57a31acbefb4ec65d85efe4699650cd6dfab24a20e2aaea1ccc6f4d7c38ea965f63c0d486eb1052ba465050958ee119cbf9f9c8cb2e6e7cbf41bea228894aedb9add81b208b3306a6585b33c43d6cdf8df13bc1333962527bd523a653f17a773f3189a52cb292dd56d89c1d2d32abb07ab1750726c55511b671ffe36072d257489417a6ad84b05b4918f577891b9b3451e0c1838d6b2a51c127007693f763dd42d652bfd732e783f0028d5338fed0840208b77f9f8c5645d0c53dfa307da11fb753ba74bb1e4d5bd7cccfa89551b4c01a58cbf9ba22e13a615e62094d55769e55414284e8966282549b5671e357f9f17852b940093c13cafb8fcc8acb2d12b1c99d9118ca7d4ee4a775729eb70c05997373b74bcaccba74c3bf4ea14174fc75e5b331fc1859dc18a2b0e616f87487cd6f6f1bc6d36c6c8d9f1f990c3fab3c2665c0662bba2429c03e8bcb5c146b0677a65b6602eda58a7079ae5c67653cef1e0f8be10e883968918b8eff8e168c5987803c8435a912e76e286d966e0a85fd1025c3c89700e4490a7f95457c4964404656d1233ec9df607c3831e9d01c38a3e8dfe21b076a7183636b1b231919de386b8f98770899841c366d3f180c0d29fbc10fa346fde10363fdeef34d9113cedf68265fe3575fc36a5cb677251ade308e6ccc7a3fa9b8c78b4b19c9bd539511ac73b4b749db42c9fd066fa2b8ba253462615be336b5ac7df5ab9ab8207ce098d5014e44062d969854fa83044c411f01021fc42ed5679de331b15878a521d293034f12859cf62ad6bda677f624b4fa90f18594e692bd656b4c9315fe8ae67175a3e83922c85e2f23e361e86c4b7642943e09db64fcafa4ef1aa2a4bf86a92556476ff4a0efd9149116485bb981c2f2b8253a4bd1ca3ab1102c208fe6193b9daf8515fa722d1a1945f4cb6d712f70557d82f55d0b98d2fe9f557a313ffc75b60303c3428d31cb844a1ed02ea7d575647e94e0eff934a7393d9bb91e76aa147ea0ca2c6b0c33068355eb8f55941a036d7a979151349586cb5f2262e827c06a0791d10040f3061734fda4fe9ea117aeaad2536eee9a4e249a2bf4de81e49dbfdcada385411008c89132f0ff11ed3fd3ecdbb25de1b60fa1a1eaf1d015759cf6784473d2f6cab7b7a96860a53f21541a4b3ce4bf93e9af3f572211cf22f9b5aa5545e3da790eea0da2be0e9700e35cfcf0a5e755de781f36096bdc9152c41a62752807df97c9289f180fe49be35173017845493e8a6a25cbb336a2ca4bb88ace2919e2c7e9d3f7436439b28b63d588f76e93a62557b2de47c24ba364d2d00401c9d7e695d7845780a5400d7e7deb34f5407872fe3a5536b2d412b6c6eee4df760245ef5a85e820f8110f706da29310941ab2e5a3c281f70d1621dc45c6764de60836012ed76b926d8ed8711b387c087a1e12d06f6ec4472edef844ef47dede97fcf1329d3aa898ad;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1cb1e1cf75e12edfad165d8903adef73108a1ae152b377d0d4b0b4506dfbbfe6d57947a5b6855153a08284ad5f5020a1c038f6ddde980d095ddeff49ae1b7540fbd282f0c3c1447aab398430952830ba5f05c98db414aa942527081475f249c2f647fe2aeb39ce2f65003553d3e02c82532939eb0643311e2be416c9d47a892bfca0444b8f77a8835687b514d8e5e4be302d85ca4c4499ea95ddfe65398a9a05e9bfba5800c5ca85f95ca181c3eaef138a259192e0b8806403d35b0816d3f128112c1a360c229192eae6e736325d2cd75051c29b0fd61a93c746ccbdad49cea0e672c65a0c09ee95c064b35086390846622237d57430a1c32186ca0eddc164989fee694a5d3577dad1841726962173d0c0207686a359a477ba99f9860fc8eadeae827d3e6b0d34fa1f35dda2cd1235d1a1f2f087025ae7940fdbc70c28262e72464639777675d7661228f7a8e97a33f5c4edf6712b03976e7b80d47d2ac228601368c1844ee341d27be5d28e564ae73cfb635b79e13ead2d91ec2cfcfc4fb0dd2ddf77fd41d23e3021a3bf3080cd3af44efacf4e7ed5d44be4244a8b1b7071eb144f708e0f3184d92598448df5d597126150d3c5e0c530756eafc2b4157c99ebaba4c8e91e47e5238e19b171f6d2de3e58e690248737d12bb3adbfd9efc5843ff931bd3a8ce77ee57cee44bb2ea6383ff40a96acbb4a04540472ea39fb119878271678d417688944f83222a2fe0a2dca31f905203ff86659b5df4174597402d787f234dee1636722a515c4fa7035ac5012211ecf52905a51a9516b8b2b0431975ffd3bba454765076ad8507303433732d05da834d6d6bc55379d98c3fca1f5ef674583e4660edd8f876ef1934b2a73c46ddfe6ab9af0c77e4d2808a580a6b0273fe6d2eb01809af39b3a446e406c4c19b3396819f26aa605267a49481c7189c64e20264a3a9ee4be9f27eb460a7975630a4931ed25dbaccaf349725ae4ce52847dea2da5672bd0f0ecce5a335dda13459fe45847f50cda671cf3f8cb97c5779dcf5fd213b55b026a30b2abf8b3f92c7b99f0ce5ffe6875cb94f9db042f6fe8e5282e1a73f2eb8c103f4ec2d933da578afa39b1ee1c9b1ee04ca1d3de65d1ba1195cc9e291d48770fc9738e2495cf75b8b409de81eabdfbd6068d54df1a79d5c74efbbd88450143d727f3efde2efbea6d18241b188c1672e6d132e866dd7ef0ed54060b6137aa2f0429213d47a65ce4dac6c0dbbafcd0eebb81d9e96a50995ef5a76e88f4d4cb606415f0f3e950a401b8eeddd609533d285250bf32ff602748b0a8cfd427a4758e27672287fc8a1c9d454fc07671ec8d8a35f776de69a0b42f29d746dc04f0541d64f147eccf142c7453b384c2fade9a14364ef06f5282803f8b5d81131e0482150ad1ab1f6c041db2aaaabf41d94cd2785df2d2760c20da21f3846399805e8de3736867835a6f82a35d15fe6f4bbdf8b75dce210d30762d8a98065db76e01e6b8d77867d3db35ab941d586a09cdb17855db4c637b76e2dba26ffa2c512292497363d337f77eac317071dc50e26c8968364696fa50d3c3fc709c53c5a972ff6ffa5a376b6a55d1a65a1c91e175fa3410a47fe31ef1fa6aba6239ab816d0274df9d3d43ec7706d75b8d01c12e6fb3f87260b46d15c34d4ed6295ed288b9928b40bbb1a59a218bf029fd92d2958b85a67828e95542017fa84d25f75a5a519c4ecb20a87d81c508ce686556b98809c6bdf56fc0c7887fc002420458c3be1d0b0069c696fd020c87da9db1d5570b77a45885ba2f3028c05514676c2bb6d98b1d6cedcbeb328ead4818bcee6e069211a5153c51d4b4ed9002a346a2a768c0f0b38e5bcb3a23518686360039244cf4eef33ab593f8cbd57d2e600b550e438111a97e3467567f5682e1dc7ff85eb6731448f99a23cdc34b5266e90e16d24159c6a3fed8175c544ff39631757ad1057735a4977b76cfa55ebb929e4ec32977f7fb97c5b761c2e5379baed1687f0c7289567b1bf79a47be9fa209c0b1d8a1effe41982e6fa3dc26e91a87d6b889cbe55d0826b6ca17be8cc40294b3acaa2f066c3a1a66cc6ffe2b5af3cda7848948398b7686de5022d31f716461371a1ee5bc31b6f7fa812bba0d9924e48344cee8aaad87bc9bb76f888faccc0fd1832c0dac6148661105a015bf66086fb2c219c73418d76d2a13016ad9bad7cc010f3f311a209a498ef9bf736cf96a1a123103293bbe2441a6c68c42b230b9efc906faae19d8bed203d9d9a1a68ea466224871fb0b318428cc7daf0c0c788cf3a87c27777e14dd7cd1b70f7482d3ab03d881e567a10da6892fd322ef91961d0401530c6afd8862f0c035d11a87d2a5d57de68dde6687d15c54b462cf381df566d369db200bd0927ec1d1ff8d4736031aeda4df9da219e49c74a5347ab31ba5e0e3922339d28843e212f5c0bbf3d53092b1f128b3084fc2e0062fad1d57a10cb18e247ed19c56a08376ddc665aa42a006e4a29b591bb83ff76c1e23f1393aebb9df4b2107b5e12c72c691760c7c67abda1206115af8f02be674fc575abe1f676f5ae6a3147db14b8aea6230bdbbfc291f4d5252538c47007d9b0e9e3a21653f8d08d81349a1665e353d60781462b919b8cd4b5b26af2168a8777d8a32a3470dd7ffe8af990529a22a8b04f902709c0f70124605068aa3ca12f250a09b5df72390d7f5ce51eb849c33dfd057eae4c4155ade42c9aa8a2459dda2859698421474f4ca605f92ca3344570316ef5e4dac6de85b3f03a50be9219eb3970ca6148c0120326feeaf9fe3d687879e1e6361d698e97c0e80d9ac9674c05f76a33de6636a9499fea15f43c824475e11957c23a8e8cd2b4b14b19c26306974c7b8d0210ea01ec2f4396060a9c563cfa8d7080dbc1611305b083afa2d598a897a8329b420e0d72ddb35e9a3085faf189ec6944a0f06a1de5c20311459392946c32be5c403237c1ca7b23b82ecefecc55a56ada1de174882ee8d149853d58abfe0a21da855f2ea2c56bbc98cb86b65cb2f36ebfc2f50b1ce6a0d19c648a178d3cf88a3eaf0836a725ce7be7b6b786de2fb8ee339dff00d34daf4cc32d648bcdb637d79ececaa1cc8399b445548b594b8e3b39effed44000bd853b38a91fee9509d0ef3e187fe3b3991e7c2cae548a098969fe37659485eea392a91749ef592e5a0c638c76b79e72571cf5d59175579724b34c144a0bbf4259453b419a56236f9224613b94b4fb096ace619178af08627de5be52ad0527d0898a7faf30ba746cc54f8b70b1342717ec44d4e6fbb5fcc18cf683ac2b6e32628cc7e7b82a6228fde90da2f4d859527718cbe2fa0fe92cdee8e7421c89b510ed1650dcd3ae94fba5f602d8d3453f69e32ce7e159f9ac58b4a6ef0a43e739d2758a78bd8a5afe46459d2d513a9397ee250d59c9d7c478e608cfaedc3702db2bfa5aec0f1f001d54072fa994e983d85fc3287d10bf091552647021c902dc99c3e991781326648936ff7f02a040dd71c1724499d774c0655a1b3d669d6a839f09ec150d6a0665628d7650b745cc0798e555713363728efa84f028420976699f1a5cc7c80230e14bc623e9b56b91ee14308f7f5ff45f91b1a64ef5d4b8aba7985b155c974bc7f02108cb73b97b23f2d2ba8ff21ae7612cb281dd249a3f49bc122e68ea2cae12b03086d07f330bd7cbb4450edac05c4152dad9f243b89314c84134c5ba19a5f2af3132ae3ed249092bdd5f682cf31206f895224771861732f42044c1869f48daa1885534fac82707432d852ddd9de6561151692648f99843c860cfad2f49276bb34659547be0935d489c859f89c4d524fd2994ce19a5e834fefa311eadd3c30627824d74172759641498aea8dbace30466be7d6c8f1c1f1749a329567bf633662320aae84911f347e559d9605512d5883fd9bcdcbc79cc1c1feaf0b6d024dec187d4e8e52051bc071f97358a9819f27f5513c6b63e20754d73cb3ddeb1d3f42650533d5b246a5325ea5c5159e41e85a29fc6267a48b73c37a30126ed7ce3f549832089e0cc1609ed266c9d3f2ea3dbe7283c239c56ad64ea37b9d222c6e24174b86a91b64f105600ff310b703523b273d93c2c1cae24ad71c8e17488188574ba6e3d1b142f0f0a69ca3c73b02a5f83869dcada8c0e8159163ca431c85fdfce669cda6c74130dc6e8a3d388bc7544332ff272f905c0d74325e5386327ecc919b58c4047bd3f5c9e951c6c7cf355ebad981156fcb488b020a599aa8b94b7382fb74fb992c1f92acfef1ec009445d0e3684b9645729169b83c08bfd95ed16a6dce3d2bf630c34ccdf7ee8615a9954cb79898de8d53b456109061fe6b40c77c4c4d83409b6797c07c1e8e225b11d99db5ed5d5f3d724e7f88c548f0867af6eaa4cb0cc8dd59a8a16edfafb9fc1ff24e6ecb818b3a00e43ca112636ea0885c9cc16d71ce4acf052a416f366b0866c867d6450993b00a7e19d6ec92ed7b067f081bf1e71e1bf7504c03be2700d4375a06336cbfc9095d1fd16ed2461bdcbb3ef55b02166f743277641d1639a3e6de9aa923bf4dcfa21e3849580d9759d50d70bf4d949e064b075300831b9780705f8aa81f86536a37f58b2edc895273cda6396936fc038b5afb553a8050b3bdfd8b079a143b0815b98b8690c360d5928cad8b09a87e8593f416b1bf749b4003947cf0a91059aedd6f7f031f46bc85cb5ae7c63b1b8ed21569ee22619c7be47c83d6134a8e62e7411e2d89f6440e57559d3307fda3c08314e3dc6a72d4e76bd9f657ba02d4fa3bdd64fc308ae6d180590076140345b494a60e5e74b95656cec927131bddebd1d1336ee05447721978b11c81d55a26aa39ddfa83ca65e3e88afb5f083b3c4f9e79bd28dfc5052fb4dc7ba6b18257c776d467c4f9ed11dc1e4670716432e10d794177797d340fea11b336015ea18bd3d6e790fa009726d2046f81d92ed4541a5166478618bc59787021c21afb3891594ba8ff0fcf6cad1aec923367ac33803b54c4a6afae3b55d456531b5e2e660ae2571b39ed3ac3f075a9576d83c3fff72c9af6195ebd4a834c94d8d3b444bfb7b0cf9f4b2c93aac4b709c6c9313a976d829a5de4b029aab0a7e26109bc12de133fa89be39f0ef8d63e0ae4e48b6a541d3b095ca831ae5080702777299cc935ef4f2798e35720ff6f563f044a15806aabbd07b4593daa9fdefa8732e228e239814b9663cac7a1f8e76a82032f59ef992eb1126f311ac49f0a81d80cfdacd89de571892a6f8ae511bbf179764fda644ecdb5ef3614c3c8ddea58c61159ba8c1221fd1647f6de1d3394fa604b6974cb738273c3a7ef59c853b58af8d7d2a5b9c90ee84774e64f1135f257c3025c891fbbf4f8e311876f3110cfaf3f732103b577d25da5406ef5115588034b78f4ef34c2d5238b0c0b49de39ccaabb9ad6335e1006c9b873dcb2d965d2ef3bbd7289d5c2df087e4d7ebbb4aa76ae320d66470477ea5b7fca178fee8ec3f19f929baf40983b70f086507fd1b7c15de0ba745ada828832eeb0c50580cdb4b4b13c2c7b07c919e60b36d4dbe526c546dd4698c6e0da7fa9e5c980aa0e2bd516299b470588c735c775e545fdd84b9cbde9ff9b49b3bc7f1a881a08a144c68ad33453cf8f424e26119dc42a73b20394cb3c4dac14d37f0a6f3d5316d7fec840e92275f5294e58788044e2fbd185944b239e08fbafb7281d2717fd2812135ab05e5bf0f356c1761cd8eb6ac165c37fdd695c24e9182605453746147310ba3dcdeff33407b16d2d04e7e1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd2b814b3bb9ec779ccfe54c655c4da25aec6c0b5c17609cb39b0d174913810498c175316aa04679eec5a0abfc4354b46d5c287cb624cbb5034e83041984f3a6c4be7838f974f30029cd5e6d04ecbd0540db397cf24c3c0e36e275844674a274f227b54f3a6c6b01b5a7698e72c6e1c814fefeaa21970210474b3db9e777c757ea8cddd65050618386d534d7d5d2d0ab6be049d57f065c2c66d25ae9a00c97d963beeb6284d25f8afc6fc28cfe09b08adee71313480290af2880f18e1057b89a66433b4e51d3a5baf623523ed89ce7395b4cd11ad9faca4f0d5643cf2625b405fc591beabcf429cc5d9a50bbf05213c913effa2fdb95a0787f34c3a1841e6c028f880c9b7e77d6b63a62bec9f2c9767d381b19c6a51730e643c01671a8793cc9ef27cae9d4934190d040deadceffd2ee2c58347b2ad198818e47cb34e174f691462711e37741dc0fd85e07ede888c6f980016592237c81d91a6b564806f537455ccda69c72cf065724de31de70dcf53ff914bb916b09f577ed3d5ca26d4d976d6d8f933e5e72d99982935bb5ced06e4d1dba2468a8d9571fec855e238e90f7373cf964831d8e3eccfe976bde7502d558bec2852b457b8f6a933c85c84691c76c82fad64e94aebd00f846462345a366b719ba8dfc75d8d708d0a1d935c1724b7ca3199266df2b860f4ba3bda20f8f8c3d6bb35e25d9025a1ea6247a6f874559bc6baac4f513114739ded02a868395190625cbf959954e65567b48dc472148e171d1eabbc6fd5efcd06a4463dc7e7022f2c133d6152eb9801548b296658a48cf00ce8ce9e5df0b74bd038c22fdd92daa6b05b4bdc8781abf3c8ff36bdbc89f7d9f333e4ee476740464a4cc6524e60a906b14033e576edc5af432583d9553f21b3348093972ef2a790a08e49b628f4fe31a63c348e3320e8f822a82b4ea7523aad3519eaa1cbc9c6bcb371156911f9faf921984dd0e3ae6d36e54e76791cd5ccc3304d455a29c42ddc1c047609c816e4d6bd3ae5915e91f3fdcc3a15138b8fe41c9e6a7ef56a96197d9804d448ffa3b5c3ab22043c95fd431d66b3743a6767fdf4be67f5b3bbd416f93a2f81cedb768aac052f9040659a1f9a0754aa9d1495cd8995695b4a0ad61445ce8d46a69dac3569fb2a61e5222f529508a9a0266c2dc048e1502eaaa45da9555e099a940f102a960c3bb32b7f1f175fa732102cfbd09bc9406369c6170f356451fe87c227b16855bdcbcb037aa6dc8bae728b8347c765c9783fcdad50047f2f97474f332bf47602c92c72cb64981f1357cb385e07469fc2c5be8788818f507ad7a76a2dc7322a6715ba9e325870e8d5d99fdc585161f7a6c1dfe596efb6367db6fd99dba219fdc29f27f04e0d93c8e64d5191c5981cf6dd42452a0d32a078cdfce62d8b911767f3c2a27e54bbf7d0e320ef7777d309ddfcfd6ce418c5868bdd431343dd6e8ec3eb92beff15a822d33037c51f1badc3b115c5818070be945e57c4c8c0bc96eb83a701bac0fff8563ba544015ed73649cc5d0b6174486d41b5ebc9410b95585397c31bfe2b96feaba06f032a04febaaf6ecc93743d549717ff8395c060f6132b7cefa1e3dcd3875396798f568eac44e78f9bc2b3ba6856d4391ac91841133e824d285bc5ee126eae266c1e52d0ad3278008b37b71631a5a54fd349f0721fcccbd6857ef16ab2f27e9c6636f68b295aabf2d24282c39159e169820fe9076c87a7ce62087704a21aa31fee2bd8bc7d054d71cab755dbbfc796f79d4f95d2c61c57b689da934ddf0c2d508ba951c14da3a377752e399b64b1e30c26ee11e740414f562a767ecd3259720261ea71d2b7e07a524764e92e1799ef3d31e9d3475c145bf60489aad8a8f9a0cfc9c5e66cf737ac902db742d96ec3804acab55ea25ab6b9f70a613c3e2c440b42121ecb69308b8881cb294d1131fd65fa182b93cae586197f26321621f60fa144c407fa3e8577d4b1068828b803cb1d66795991fbe88030bb84fd6dd65f16f52e6162f9280a08c03ffad94b75fa3568c0641806033ff43fae7ae949337591168a527e9fd215cca10ec65b739aced79652e199145f7518751f10704ae26d31f8591fad8ddc3bf845f1a561f12b5602aea47f98efe91f16dbbcde522fe450c4f8b1706d98ba8787b889051988d6bd4e1608615204e6d005db107b8ef1383194a14752d34f80c20ce1d103d0203aec9fd871fa562f7a740c6b743c297b2797909bc61a6dd4ef65d5341c7cca4a43d94c8a66878bf197da79e58e8bf0d75d3dfca65bc8eabe375189755bcbd95855fe7f178b34c01f4fd6fb56c49d45f8dfe21bbc23a5d145c0f16014634ed0f98eced433e3166e4c8fb8c385487f6e16701394872b07e0bfb16c4edcee4ab175f0014031480a4ebea1836aaae4219b5d2b21cbde0faba7903f0ef90cc5ca4f78132c48a24b70ae2317479dff643d37e7ad897fde48c4e7fa8ef45dfb5c04980884706843bc6a6aec017fab7d30d8985c47c96083abf3530821a7e7efb5f79d1e39ef25c819b171d0cdf3fc4bb508c8f3b77726e5d8900bb1851264fab822e69e93dc408fe02c03f5735e553fa25bc377b2aaede8793b14740a2ec4fdb1cc988e0d7aa63b8490fb1f4aefbd5294fcdb85dba3bbd3c3badba0cc386514a5b414cbce6315dde0e5c24febcc0714698d74f133272546961d28c071463df526146bc39b8dcf8e73180f6785c9ab470115de863b0dc556c16948083bf02d77fe89b864ea50fa47c5af8cb0fb3d0e9edbe333107a4b367bc1d597a351d28dd0536b143825667d34a31aa4449fdc721fed69068302dc2742743e597ae7902f68677da418b84b3246b59f5bde8037118ccbaa8dc9b33fb9ac0a6a5ad3be5bacffd3ee573853b91a39844b4068b08a72b637c72e705ca8341b8e4295c40c443a1f528e03e23dd87b65c544c200f77bf463df6c06beccc347d2f501dd36622a47ca0331b5d7c0254a3aaf42e737557c254acf69f9f56986a673118c5f04da2fe05cd8fdf740b615804398273a1ed58bf89fe16b05dc65d8454c1f1dd2211da96d97dafec4efa1192e1877a6fd190bc54b5e15e39d8d147de8291f6d473e6475bbe188222be03e93979265e8f21a1414eb7e1140845d977381669de489630ffa4247c6813fbeec63b8ec3bd0b4e1c61945bbd90fc5f5ad10cb35727abfd9e94cd8adb1bc89c8b0e773f6e975d0c4e07c1419ec3fbbcd7b9c8aefc1e509c1d3dc2aecc342bdb6dc7975b0cb9136a726e47a3db3f5d369e8f550823f491786e394aaa5690e04c66a8cf408057b4364dbc79dbecf5a7a0ecd236973c3a8e947ab885aa6b82c218334e878f74dd8001855c897ebf2496cc7c247a0ec679de21d1722328889d9f3076c251f47a401351ea6ec2e3480320858b1b4ce102c6e762e62c00ed3484cf50cde985bef09a4ad21cbb64042e87234586cd497eecc2ad847ef8587c3f703e611e9066c30f13f0e57a420e488e803ed8dadceccce4e6dd67a3c85b07f446943e65deb48b05ea0c4b9e213514c6762c6a9f5a5902c1b9c30557d0cf9af669440d9c316a3260bb3973efd0ef7284bf28e7a6529a1279893665043de66f57204f17e2e9bcb38833106af5d767149c257c8d319b49052b2906020ee7126ebfc7f00c0ac12a5265202c85b8552da07a25d4e2d5ce21fb9c289d6366697355e8f7ad9df3b7801f22a4bde41c2eddfe5e16d0788d89ca6fb44d3438a96a533a4fc515b9753991ae146b2360fe1262c88891a911b963bf43a67ce15e5a6c02cb61d293b5dd7ed5f8b80d4774f7d0165e1e23e46fbb1a86ba2b376afba31d189fe9db8d635b864256d6a02220b05303c55918b30f9680d09477128d7ffd54e8a25d64fd856cadfe0fc09b887eb9be0069c35a77c4b7525ff248d2d23093e568971bc5efc3ef5ecec459a1c683ccb0e6a514c0319c63627e3b7ad2ef02030fd8fa03ae22f65251f18d7b14d7802537fa57793d4fd30e2c80e516fa464d8cb46e0f98f71efc8586b2745960cb2f982f7dee11ce93ae7f1f3f3239d339a6474cead1c66076897090731fe523ff0afdcc3ff2e82ca84bc697b1a3b4f31c5fcc76ec866070953136a0daa105a808eeb9b0cbec788463996c52dd5f9f51adfe98c68c081faac42a3951198a9ceeeb5b316fa1e9fa54433c4090b3e0bd1a969747e08705a6903c4c6db370cc7059ba3abc8b6d24fdabe8df1da45e8378f6431296754107d640799866a6d6d5a6a6a8b27d32d9d37e79eab7b05fd2c67f4ad9d2fc77a76c89deca949fd8d3fc8c6be251923fcf34b10675cb7a7fd6e12791ea0cc20225bdcb8df8f5d5d14aca1647af5a6667619235cbc47942fbcdfbb86a1725f3bcb0a3d2298cfbc696647c213776a4e415f75ad1635d485bafefcf6b335e7360d75910077b41c0b7a716b5e929246ae396064cbe5dd4c198b4563e5470b9f9a594344a1fdeb74c7bf464bb00d14014d586ea6b33b9b35bdfc432825e7855f9a9fbe0aef29a71c8c99d15ee5e7c3aafc74068fbd20d5194685cb87f9a32d23c75a45dab3c063f2d86c6fed973d306846e855971de62040341ba98508263251dec7f861595184a0fd0f38ac191232f44b97776e1916e153304496fbe66464ce70883ceb3720c1b552d330b2fb8ee5337c93acb68b2cafc2e3e7f1d90629f2e9be667f0b2a86d0300029454aa78cfb5a87b30b0f7271983761c8e724b20663756d892179c3c9f8d398be5fe69305a0accd3ce0cd38626e7a9b3f62398a7289b892cd53fd153495522626008ece18469f0ad133849bc1ae904f5d3e3e0a35957bb237a7dad6f558ab5444a887fef0a692d09c5d95c4a564be816ea0c42add714e41acee4cbd19b60431c95b1f7badc32680753b7131d329ece681c6129ae062b5ca6cbb9f32c1361db42ddb9cdf663ae4a3d4711395f68d71493aacb45e17822d3223f21b313b8218787f154b8884493ff900cb429f272be87e675d8d16d45c09bc2cdeb8eedaab92b3454fb56d31b2dd738c6b9370c82bb185732aa1ce80b8e8f1ccf23ae07d6f96e3a8f5ed4426ff27e40b8040a441fd034b45132c4c39cc06efc2ee119e88677ebdf060903313d1e31d59aa2ca85b6fa344cbc57b0194587b42908fdbc11694e1bbcbf93a1a259f2a3381e511fc4ba896f036f2d803781a2691c5030cac22ebabe5eb9d3430fdf24cefce28c9dbbc57473b5677026a181b6f390156dc399bb8a1a8dc00e4d0f56187a23728c4e015eba386d366b7c7995919585e1f5b1c4d838bc68957ed3033eef79209a4ab8e3568c5e7eaa51ec88f73c485e3e68cf6d74b2b142004087b6b03b96203fd91027c4c58f12f63afcbd4860b83754e7352eb408c08857eb65ad83573ea53aa7eccac17291b044f38ba6f1525b74a411d6516e5c98dee4d664bab7d821381608f7d82bfae8fc6da41b6de0240fb77d7165826d97a7e5020046d8e2d795a685eefd87c4b187911ffedf045aafa1d7e0be31839babafcf454fba8af0266faa367b8de652bf0a16b29d4e9e9c3e83f50de2e3746f5013c0c40662fba952712ca0c4477d3e8c259f5c1afc552961038d8d502b2862d715b3ac867208236db5c6007988d78107c98e0d7c673c5bc446cb43e19b812e445d23ae93bde5ebbb5ac42c646f47661299507269a39b7d2734aaad22a0e3eeaf7b2e13881176035e4a9adaa07f48d6233339b0e5c948d3a9fc78566215204bf1ead04011ac73d02733ddc5cf214cad2b7b581326736ab0c51dba84f227f1c8bd2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf01546effc7cc2336ff44efdc797ca718aaa5af1f47ca5772b8caecf52d80aa46f12b2dc26bd5d76810ecc8eab7f7f896624bd10a432777cd438834ff0f033858845bb5c9d59959c50ea81f18f8061fc07955ee5e61c8703624b1766da13517691d8fe82ad6bfd4100d72d57ee7e2cd5a92e02ef754d0d00976229505f50cfc0c8185fc518764aaf378e5503ad0a46177ee7915e4e2544dcb211bec2f8ada2d7c497910b0d183170926f2a0b74b95e42965f9735a30938ec0002b6be3d1ad135d1d8f36b5fd37e941f63f3f2e9b03569b1e33fb275fe0a1b06c71d3ab0c7ac1245dab38496b5469cef079cf7a36dc0c61d1568f8ca0a4ffbd55d180bf71ac70ea8f37bcec4760868872f11d226228e5bfcf74c884343a2533926e2e590049a97721a0ace3870a7abc8cd472e89086e73cbc011286badac6b5298832aeff090d6c97baca8c11147e984ebaaef6bc5d9993b5c3e8fc9532871392c9c0be1b126d4d3cb15d0c8293e0bf09ef1864bb44c4e077868146ea5dfba9084187f9328e2e2e88d54fb9c6696747d4e33387bf3a1f6321139cc398dcacf8823577acbcd9f61edf4460c60a667243e125ca5b6e9a08e99726ce008ac18b9d3572633b183e92929cb2de16c1784c4420bd64c4afeeb31274ed55685ded98ddcf74fed4fe275c65096309cfa7641b56c17afb13622b1b805d7d2322a3078f13af8f60e32d882174f66ec33b49c1e0fe79bd33e6be4b9d877848dde11daa40bb0f9131fca08673d874b6bb99a1a837cc833047c523948c41e435473a4e7e2f69b29e2a1ef91370b40fdb0730b5953bb9e96f84794d053950efe3e4b1699a97f88daced6de828b4b69b121104b179558700a3fafe436cec5a70162857e76ab6cd58dcae0e1e3eb36235ad103ad2ce0355a332467e06aa40d353eecab6ae38a05d7e30e399d53f24627b65eb3362bd752364a25041130259d1d845079857dabe11307a4eb2ef703b527e355b3da3cc4acf80962d04a2b9fa7710864f60c562ccdb21a77f5d934e7b3ed8db422fddbbff6ccc30ff884948d8c100c0ccc383a2759057e89388e4b399d29dc3b37863e1f1839d8a1541768c68e4db6bb29e7e5bf66ad806dd7e07bf543fcc3444ba99715f083ce9fd1d0159a476b384314d0c0906d884e0db648b1ac73c8281c4357b2dd3d135d5413f3d064b105bca96d49f68ae08993f12c3f1700804e11a5cd80caf579fe84815b349727410d3fc03c6a391778f7c1bb3084d6282a5d2896208014f85bfef89b27c170ae78e62f64ce06c50c9b3e39e9b2e5fbce72fb356c4aba7fec21fc935e96ea75a4095ad817a68c2524122309a6fa04486000781388e263883c5f53572a751c39e5f14989dadb34273fdb3ffe61cd1cd53240191323b2ef546c8e1b4da715c1fe1870dca2ea6081e3a7f60526d908c141f8aa60f56d7218623a846ca033cd9f2b1b287c7efd9bf528ae6169f2815154fdd06703d1cd1e96ca3476b6fc5e3c33faf5e60498071da05796433ec2731a6a17e8b0613fbdd86c6dcb8376b4f0605653525e8d99193dd80cb79d8b16912f01854055ba6def1e3ccbfef75061f320a5465d4ccb3914eb8c4804ecccab9c99a2f211cfb5058a9f39aa05e2cca04927b3034b34d79f6c9db9e657165c9e14da22c2b2dd120714548b7d40f8f853398f5921f154d4602757aea58ed27867dd856f4caa29e23dd8ab1d94776851ac08d49b70003621764b3bb8c99cb8f42fc7d9a6a2415156e266b047a02b850b38a2a2e5f2908d519a614a728fcd0fca9e51c04097691e297b45f593625d578dad7992539681f9ff7db38f89145845aac660c27948284884a0aaaa5e223a0cbfd59ec60063360ca8cf1c31923639f52ea1b4fb222c0282a621fbe0b988be2025dcdffbc6597dea6f2369a4df23d93dce7e02700446b3ed00c102b4dc6e618749540182b5423278547c3defe27bc54adc658a9b8991b8fb4ca1fb707bdd13085678857670e899c6743cb909221650fffcc645b5c379fa58d5fd4f30cec782ece177dd839ff58aedaf440e5dfd983dbdb275841633f55b48d5c15976042ae759249d8e4f1b17f0bae4a5f797bf8972b97dae3495c3848568eb64b3bce397a25ee96b62b817bf681cf2c48edb9ba0d90c2b57988468f7ed3232ead09c93f3b4a86d0c1e014f62fd26bdae1f1596424baf7918179249bfe89713ac7f0084c864b4ce500c25dad1c50b0bc1839a5fa7ab471b6338ac63de1088f15c1ea1286ffc5635b1d15c5bfa587051e249954b28a1e1c31a627a77502d8bdf72490fe2e4b68d38659ae016a7bd55d280f498890aa8411391538383c0e556a27ad953e18d792284c6980e7ec2cb2ab447df9d325b32d116047a49f82bf82689a42be17c1ad7300ba653ed35c00f9d67cc229e1fbc064f92f2c61d14f20329b357f928095c532aa09eb5d3fdeb096bcba931d2a48ece4fc124497429ed5dd914cc19b5134d54bb6bc1bc946ea34a26f21a5d835c48f17396d065d2aed590962b77f2d0b0a0aecc6fd0b307fba9eb377fd3aa416242d3cb6cbadf2b47bbc4b62e14208d69bd5397f23181d89ac1e02ffadcd8c363e22f10da5d50db25970803bc7ea243ca031b57be3007916067044e9e78c7b57ab11aa7c0409b05f930898beaca593240d462884c3441c776ed80ea820a5e4e7530b386f110cfdb39a420a0f7146ab52182d4997995daf0f967018cef5a89f83dc2886d89cdb5a813948f1df2a8c00c6d5d20b496dbceadd41318934359a5d109d048c9e4c78256b6a5942501ebdc64a8e32487af600843f481144339cf1038aee65a7ca5d14cf6cb737b0dbe2f5e36459b47c27fdbf2d56077ed3fac5adb861538e29d038db24b0c5cc4ec69dedf773f6b63e813ee5138d80cee9151845986ea576dc801888467c80bffca81d2f7688a6178c8ecd0ccfde6ea40df8675c1ae0c5db76404ad04a681cf2808ecd7e6e8d9fcb2fb3f779183ba5c87aacde6079a8697f2c17c060757a0ab035d72fda5e8c4d850a9db8c70eac454312c952366d6542ffd816450d269c3d42093c1568aaefdbfc9401ececde874d5ba18866e78e848b4fc9bd1ef23582907ef78e2c8c185f5d295468e1a9065fb6167d7a98bd1582b90a2a15eecbb3d309d14629212793d95dd2137ffaef873dc443792bf4ba14df1f05886d0e429d764bdaea19631a0c664cca7e47747fbdd163b37d748c2fa032978ea3f72d17d3e618e65fffab7f17b74407fe773878dd3d605af45ec971fe78591864d64e7ca8fff7a3441479f787bea5ec10b06059b7713ff0e5968d08aacd5a824a4dac0eaf1a05280fe599485e917b1b8780268d8ba3f30c633f0a06503d8d5b544c9011e1ff68539a6386b66d38a93384d11eb49ad9d2d96b1780f26c71253b3f421d1e2a264258cdeca9bbf2ce7e41a0e7c49d99f55732996f7ce74d23c88062ed1c42b5dab629da5b59916631c56e51846d6a4c8a901821f6cf37d02fea3eacc10e882690646619f571bbc14c66cab4e2ba3faab9835eba3901ddad9eb6706eeabf2753dffb6d8f54ff5927c7cc2790e8183bc3dc903b2565cb677931d3dda36b0e2d78bf19a7983fc5238f20c23d4bbeb312b02f2c77a48ceea144da047d15c245ed66cbfa3b19fadf78d494015ad5c119c72625606ecaf0118d27eae87389afde6cc88d71155146f7775302c34b40911d99086735dd3baaad047d92912ecd250fe52d2fc88bf4e49a8f3f135e4cde64080ad2dd312a66b9295765674f8f3f3ea72e7612d623ae5f5ed439fd94d0e28fcf72d62bd82729c86148e54d5d4c67b041137a05454b0591d4c9d7b83348a4e128621fd23c46fec442ae4d6162dfbb17c403e0ca67124836fcb33ff73c0fc9dd89477eb752756f9275c7c68ea2d2c9d03f498f44757a37dac1da4f77564bc864307261a540b134649741f941afdc8bdc0ea2d829bcc2d59f4d37c302daaa255ca4d9875238bfbb378de656db552b71d2a27a721625639a1646d2152f90deccbd6208e8112f937cee746f5b22908d06186382abea3471f591b9ec51c11c920b75d6467393c5738a2faa7e9e6d0e714c6fcf427febafe5975fceb453798d06307c9c5d62d5a2ca6603d156430b8bf8be617d9006ff83de1c2a491db7edffedc08ef76290c82f8054cba01a07c84fd56b49173c59df1bf395ea4eb3d99367f9c4c383bdcf87a905595b014daddfe467d9d3f7f995e6e3efd2238bc69e15f39d00b32959eeff2d1d354920da2e77ed218de03f8e22f5ec722c6cd5822a9fb1b1f027e9ad4375c9d2e98ce5256949fcd3811159b11684ef56fc8c4883e97c5f30d8f0b6663e67e39f6f51c92f45c00d75490ae3b6a1d4331d54069a761158b7a30de358dbc422e705a9a307ded238fadccd70630c687a32d8e8e3735fb4c4d0119fb2b8401746ce95690585af128d007689c28a5fceedd3b1f8c8e21457e6e930b5581623e930b953cb9cf884861afa107358095b0d4415517ccfc60c916ebfb9c0c8ff78d5e813eda99dbc61fe77c3b768088742b92e40b0cea174d5f3191de61f2fe9261aa47416202e368707c45a5a125b03b5a6ee9472be50a9e620346c7d2fa78a1ff104252a4c5b8f2c00125f115ff84d4a3156c93191b5d598534c564adcf2718f381ea4ece8c3ab92efdd44c10a3def05bead63d3ead37bbf33cb638894cc1840a9125d756b479af8d5d310a4911e9baaabe4224ff95747c5c9076f1d49946acc72e5353d7673d779f2aaf716087ba2185507d73e6215564a50e5cb569ba8d143607ab42c0f979c470b4479aed7d2b2fa568f5066ee3cb7cb14b8ee8d50e943d0cbfd2cc465f2475de1271681b97937e3dc11a9e415712407caf4ad52ff0f4bc44fbf748b92e09d8f2d2413941c2018f970e4cb822f271b93f53f50548cb1b8d2142d4add3a8bb16162a85109034b272dfc3fc6a30af29d0c682e64afd71cf61dc2b591fdf2d0b0fb74bcf96dbeb4d1def53ef2902b1298100676fc1309fe203246dfedd73d9c5b3de6e77b26847f456575a4b39fba70624acbda6bd19bfed38375fdeea5aae16b5466a31c6ef7f355bc478877508016845aa29223c62d86ef4c4c4e8b523918ca47f474db6f6fd0a4c6b72e57a8f471f710390ef983342c6f787de48d8ea41b328e0bebc72b5c7d2c76c6ba0aa4bcb9aa651921c96ebe637b9d94d10b963d4d18667ac6a99ef04cd52cc9dd7f95ddf6b491a9c025aa733b4238b63e8bd181e1c032aa91033fb173a9fc0d5792b2aba9943c524de7c4453c1cf1e7883f6a0e8a3e74e44774b7fc3a5c32fb0f0880cbc4424a8f1f8c99d2dc67d8e604a082950ba8cf85ffac93b30ceca22534c5fbf0d9fae5305187f25e0cdbaf7d855028ace24c8c9b08daca55e9766cce8c005fe56b05e48ad1dcc720ddb9f6451f83b574b1fdaeb88f18a79809f067ea01d183ffcb8141bc9972b70277be7222f594bb7990e1d0690039f4f0d74f023e7e9d3245fe268d3e01e36290f3ce38a3e34354b3f33c7eeaf257d13eeb6f8fd5ebea8a77841de12fd7edbe79677da2ed5358c163d97cbd4dd36b5df01e0ef3690744b2f617dca7a9192bfd60f948ad2f02a7ac57e765587239898d70834b1a7115a7c7c20dc8f88dd31f0326baaeee663ae2a5d71b0bfc1616115d909d4b9b73986b86be413fb479588527088427f21bac2e8deaf7f1bec20ea86d7009956b8de820b376b3b4af123ec47bfbbeded5b313e7fadd60dd7321f9deb4fb9abd7e20cd54cd0f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h265d5022bed58a6dfef46d8b9ba1e817b1e806a40a0ec611bfa8534b79330109de423885e09d08cc9f60e956307328f8a47997c4751c3395c2209e7299c5eb5a4cf5c8c705643ccb3d97be3a331a4ec5d1f77a86c3881f8e0759752243af63e138826b2622d56a435e2e36e512ef4ba9e7b64c87af746871049443051edce59cc843b1cca3edb6e7ffffcd70da25c53840a8d15c3abdec96dba0ff96101df80322970bd7bb9fbc09edcb1b24a7c3c6008c30fe2a7b6142363df9fbd32a106d13d007a746f1c51de8c3422daa9933704c39f4e081f0f2b8b9ae43fe3f71ba33b6022ebd56e3ca4282f92fd1c5ad86d80afcb2aa4fd753e4b7857157d27d79d0763578def1800983b82e1b9faa92a9591764570fe8ee002d2c031482fabf815a292c119454dc5b284ef91e2ddf81d022515a4b9b6aec4c18c97479cf09814fb1eb5237e8de16bbf445e8e7c73c997539d46ff7774c7214653d0c848cc5fd1f3746828eed442546976a59d062f549230649f3937d02e3b7c75ef326713e409c266a04970b5a33d66b141e06036062671376db6ad33143264aaf428ff38ec71972f82f896524077ecb8c308040f0f9cdf311b198ec3ed5936a1257b7b11ea3e3ad44144fa75070d87919ac460cec0619772879a723394a3d48d666dcb2983013c20de6f8a269745d76d7d70390e494d727a4f8e47be7337b4ad96a8f230c0df203a850d60f0e1580c971e9d3000417b4931dedefe2032f433bfbf33aa7de4dff369bdf77b186b032bf84f4d246e6a25fffac3b6840320dd7f472a276f379d45aab593fc421501750e4392442136aca308a20e79159eb61ba3e42178b07836641da27c07277184ac0903158cfb3011724e34e16a9eb59c357b4daeea72cbaceca86e03b95b0e9ac8b59f981eb906eeaf712935d3282a40a215a2b60f72ec27c7211a848b7620204a5f4ab1dd226bc56fa30b4fe2f1c1bd7f3e1bedb86779ac1fc69a78fc584892259646ef347bc914d2985872178c0290c6dcaad6713175b6df5355355c4f817219702783c1e6884ec4b9a24edcc6d703e7d77aff3ed78af712553665300586e323a492b6ec286974c579d3175dbfc12ca4b0ae401d2d23053b0eb528b17d831c3dd8ba2e19c7c958a53590898e506ec0755ca26b842129272a3fdca32eca12aef8e46c3841d0756fbe089fc1a478ff1c594f861d2328e139ff294a6672e0c018fe33fb240ff5d312adea357cc87ff7e9b865b44966a4e5d4d1a83c6bdff57ff9609205b49c01fc95f8c46c0196d3f95d37fcebac4e0801b0efe9ec2d507f7fb7716b3330e012cac3691be0a1882dfc6a26e2164a7f829d59945cb6d282ec9515ebd382f199391d6a07c2a63fcfcfbf7858153a7ccd0be39f95c98ad085afbebed5959f27a2221e19b9d3ff4d8a0737912714f1f029b3ca8382314957901b8f013cfb879aeaa59bc677874584780b364df59c4a6e179b91529c1a7f2d76bd6f0a05469b827ef8b313bbe49df37dcea075406f5484316ef1ea6449ecb64b6e6d765418a53d5a76f9bee76eea5969e5e606243d6b864624925d0d4f341cd639a5029e75794ecac428ba8a82c2c0c1f3da4b2b5551810792898063a5b7509dc974a86d46cb5eb508685c5532ca2ba0f27e01398018e36e60aac354c5aa4a6cc54969f7ce866862ebb92781b708917f6dcd9ae4cee7304738ea104a5fc682c170e5523dcb4412a267c8802758895024a0ec1bb0fbab61375b7c9888c5615b332513bef2a7014a87d8b328358d27a59bec1641b3e6107e6acf615034f13e230e430454db5caacab552d3ebf9ed13a7b480a0409072ba5d809d430de5b96512cfd3449b85076003d114600809538ec3fef61c4a9d2e11fbc293528f4c37dc0babb18f38b0f76687744b7ba79db709e38aa8d52557e01eb591cb4d786a526414570e9bd1b5e50b3ad425f24b43d5a7ff384109ddaea539aff75b9f2e9cbd52635933ebb7278207034f9b9ca9eaffbaedb5b6cd6525333fbcff0b530721574df663d5ed0ec924f8b9394b7d3225858be1bf5d758f124b690966f1634491f1c5ef39fb48bbac9fb9e6d419d412ea7c9f238e43a753abf942664ff178e361ddacf81d00bbd5132b819ec4901275b0086cdfaf5cfd3bd74e9ea6b659bb69067dcd5c97c68d1bf99807e43383d9c05c2b666e124b5112eb7c1d0f182143aa742e3213c79c0668d46878af929dd2ccd8947d74cf83158e33eecefd5501d180378ff384581c4189ad1e215bd97ddbf6195a6a083dfbe5bda97f5f4c5bd25f28c4f16aafa2a43c2422f48933a8db31365b568603c35ef7d4afa9068d1d01eda2f281a354a14fd2f7d37e8f3618a0cec106096ba4e57d641aa9162e4764d9b80b9d9ae8d373eed813656a68efff9ed99e78f0cc6e8431186c4c25e6cccae76870e6ca007ce9d8a51540e8ebd452d8317789cf6aa0771dfa927b6baba00fdc53319ec868ec1e544a37561db1ddaa08ae2aaf4c67e47c1739d134a71cb9ea6225d0940552f17277dce594e74a34b9a462da40711c074c275c88858fd6199112bc5b98e7f42b580a4d536d737591955963153c06080f5b1e64450bf1c1bd7757882226917b7597e3ef664cce956fd5bf2237e10a4972e27da325f2997088503b7f11de988825adff201d6c988ec70cc98c70e5cecfe3baa8181a3016569e78b9dfdacf8450d5251ba876a5cc41c1955f080a9ffc1a2d11372ea18f5c8a0863d17f9e87cc77ae16bf44648d77df7c6cb260762b67f206e88c8adfd1efbe2e4001035603fe2a7b80f33ae8ad1f093932b68d46f9c5464747881bcf9508189833fde1dd1ddc4695191381eae6e56de09c14ee30cdf324ce9027f1ddfe7c0de86a230bf908efc04cc224e8b46a6c867e2790b48f1be986f3b3ef32fe836a668d900ba59350e4898cc2bb1be6d4bc3b522cdddac9375789bc9b8a4014c4b2961ef2f6104da56ff5b9ccd81f452f6c5c4f2fa69ef1effe90e5965ebc01898122d536bcd5af7a26aadd687e7daed0349896529e77580d9d22c68c7dd6f0e83819cf69808aa21302ac3f6d49f87519b47414828091ec929f1ab63bc280d16536f92fbd94e4f982716bc9776291b44785d72519b7b87b81cfb1b3b5c5ef407ed23d1ae20812af165bc52bc2362f3be43555bc4b66f5d5ffff3ac7f606e4af05daecf82c79c484e715b47244d6d4c1f3044f8a954e65ca199c69ce239d6f74b76814f69ee62d54e077ab76381927b1a0411f8f4f5bb0db3b976d8a5a403459a17b489342164eb0361394d25ac4c78c0d94534b0c87515884c3702c0629c3e3c2b16a611db8dd7606cda9fb3963f728821b064ebcf8e25321dc1f7ba8c9c03f5e9be1f9b354bfa97e67a5ff49dbf3d472d3266523e15d06081cb9fe70adff8c80fd452ee1428f7d81bbd784e024fb93ee644ea3ec20b609c97eff6ff61be3ac18ea706610c19b603a901cc2551c5a32a4455b6cd9acf36c54e68a0d9cb779f0292410fffd318d91f07e77f7ad0578b3f42efe461fa3fc6c9cb7eb5bf0a0b92c4ff4610349884756daa3a0f11d35fef962e39fbad5b4adb27cd2fad7c0d4c929d355f3838d7c11405b65372ce0f9b37bcc65393d838c1801ea7562aa561957a640465201b9c7da0b57d27e7fa4c52ddb902929a16c4fb08973bea330124b162d08d6377b6d6d75ddaead31db1a2cd58c48249de2b961590bf01653b3e99fd127ccc3e079ade11aa1214ce8080bcd092354516ee3d64840fd68499d810283131f20a595f243df15734df195bd00fb9acda51c2b11b8dd00b366cd60a5e2d2682065b5393ac74ff6c4c145c21d99b8fd36e18ef62c267e64331090b72b944fc6cfd64c2c45f096b23afdf6ec4f6b1319f4a57701db3e2712902dfebb01bc3bbf157c60cfd902b2baa99bb9ed0b2f4bb563e5ab8f4cc1fb03789c79991c29cf7328449bec2ff2bc9b871c94cd7748b5ad32157c9a63aa94e9070934db8e7c6fa6f4aa0c3cfa44e3058fae1e8bc7db0bd0cf300d3d367d1958af4dda80bae39e7106d7101b185b0e0a18cc20be666292ff7eb4182c9fe96d68d0b9dc1acd6758cae2643c6e2511e7a32a1924f7a7a4b3e4ab93f1a39378de3e2635cd29419491c1723aad3c8830f4f7e7814cfc173b46050202bc40a82a6d1472878c76ed950a83724ef38ad47a8ff03af6dd195ce1d67ec9a34c5961cb8d741c861ed8dfdf80c4f562ade8943d43b279eb993d26663a4ba822de22726d4114ca6200a5e0e989dcf9a1ca1ea6eb1a4892e2e377e9252094fd4435c06a8f21007cb7ec23d297a1f88d0d182b7c49f38094e5a53f0c15ad9863bde1f830a90940c5cbfbaa146a7087000e00f43e3842af6c43d169c7e9493fa6286deab39fa29ae780689fe0164dfc939d37462af1278567ef01709a9e9d6fd84a35f68b34d3fa9802807b95fdc00526a847d7b4c811a054791e1c3ed0817180346609302125808681eb3f88ffa1b8ac65283b2f4020a96ca7c386475caca48933033ee357959fe20e25a3618f59540d759f84aff58e17816ceb576dfb90a34818a58db9c6ba82a41670433b8999b126c3cf5c83039f95f1a2ed1801ffc950e7821574719a6a586134dbffee140d3b234b62412d57a37ec5f02ba7168ff78b903d2fda89cce6b53e628950b61207d427406086a7272c0e01c0ff6289ef8d30775e65666e346d4c1a2862a0a5ec9b60e98cc058706476c23efee237b4df24c32d72fb5f666d5519d9a2853d95954bf90573dd7b2eccb78a4f1d71e65a0c530e1f83f5112d56c2e9e4d28a915b06978286606260cea29daab73e5bbecf1640d643b045870598af912d5fa90fbf7f54e4293b0ede2ac37c18c54374f8c968f62d51f2059285f6777c26b3abc2f6829c7e8c677e1a9b04e628efaefe080a94dbacdc3d176e6c00542196f654c0ec0756b3d542fd180c8d5a2a56bd30abc153eb2955ca2062d3bca49126d9ba63642fb65f479a5ca7b811084b8657d3390e0abbfefff685885f56f03423a690fb80d907b3ef851fe7e7158c9cd4cb98a5d85417c011fb20520b41bf3c1a91b6475ce60c6ae96d76456125e134a7afbdd58d09ab546e8e647a52ed0b4965257591cfbcf670d12d7a6a4a56a528182df985f2342ea03081b11fc8a8e09ef51bd560cd66fe22365aa379decb8b5eda3d08932d47d37a038a524fd1a1c2e07e21ef3d2051707185cb90934c538127d63c6cd2097ec0ca54a42dc05fc70148d7e35dcb2f2add9255286ad891ac79b2260e80d724468eb8821bbbc5fabd5053485694ad31a7814f8dda717dad71e848dea84bf09ba063cd452e4a6e2a99b562f0838a94934c465759ed9218bb8d79079270ad4846f2ddb377686a1fc01958f329971ca34e040c6a2048fca6331feb1fefdd791690581910130372d78201e5e364192c7b0f22fd5cf488e12f978d48be49bbff2ca89d4a8dda1a866b57ffcdac2f15cfc42de8ab0c7d8e1461530fbdde58aa898f9780992959143f2b3229ce2781894d00fe835e567ec2d169770a1e4c1eebcd5b2cd7d8bcc1fc6eb57da6cef9a0c05e7d1182b7e96b9d84de358a84b26ab0cb87ae5051d4a3b0474296dfa4eb5112a391f2b862846692b3b61b0d1131afcc1bd5da119348bd099eceea5b7d49377bcf9cf3d44d3df8cecec50e494ba0e50ac8a032e6d4efdfc8ff84dd62b3bcde5f638925a31f28be9c34e99efe31428c6127400a76dd1b7569b193cbee8100b68b3479ce21799bb5229fc7a581bfcba87fc4a13;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h21a281f1c2f2d4c4afcb0b9fd04be698e72ce021a80df529277939166b2634fd5a254834745ae3924cb1aaa27f18996715d42cef876d738caae5c429e587db29458269a6f047d836f2843b08d4c241e032e0577e5bbdf67931a935bdbfff99d47252b081a2c68c7323ef6aaff86855c2e5d59e8b1df1a79f300c860134eea36c439ff670764f8d13c51c80038257385f502de5fad8dd7134aa45ab58ff6fcca318275e0150c57213cad9fd03fa30726a9e421045ae0d4d77fcb56d34937c531009f853b2c6bb38548f727b52a30865a515616f6664eb8ec89be3d83d45fdc8bc5ae0b11eece86579b6979296a965100f6f13f0f954dcf27c75777328eed9121f8ed0d255606d5355a20810a2b40149ade493e5c7d1a36d1b8fa58e8ff3e137c5663610f70a61f5f53dd1a4f9bbf819ecd546e1f82f249a318ca3a56585bd70d9f85aef6d276b7cca4aa036c970372285910c65a50b022fa668883aa070e769922eaab703f3aa27166a627954af39536763d45183d83065efab65283831d5637dbdb203bf5451aa224dd13e42af5d0b85cee9403c5089a053a8015825ba0f300e208e863fb4df049fc775aeee5750ba972e1d5f71770a97c1a1548f476aba53565d4a56d1e73e7162269d3ead994e3884e1cc51b54cb30543cd78633ac0959298a9e5487a4c73e7133fffdd332589092f817c0a136515d54d26291e86a53e61e36ac22a40e2e74cdea37e77ce84cf209edae272a8e0af7788bd3dc93b54ae93593a87cca3063d033eecc02247f500e70e378ff8f97e324504abce290af8b26ede897afd418951f5f6361edd34467345624ac1eaf1bd56caabd95030084e9998f11cddeb0033ed12703fb51585b79be1590c7cc3f45f99f797dc697e00b871ac8f7777f2bfed0075c534f8fa6fc0bfbdf9291265bcd5adc6aa643447b36ee4d415014ab29acf944a31432c9ec7f3a94665a0636151b12780e8f1c25f8470d9bd9c85a5fd8084592ef5c1495f51f30ecbf9e3b8326fab4936b9e2154a1d11b87e96b79f68b2219bc4bf662a6900bdc58e56099c6ba6c3a700ccb7663b3e8222fddd216f40e3662b4781312d0a64e89be6bfcf8122c94ca08ccfeefafee02e2618fb33ecb2cd63d6331c1044906daef507ad9a9f252279f97d8116985ea0e0e1239132018338a39ffe2f275f2de2b5f73e9c071a05576be9b4c2059bb76971bcd7150c810451b9d0963b2787c3e7ef11f946734145b093bc89a39fb98353fef281b9b9e6fcf6ce38b6f20669c3dca693d6586ad5181bac01cddb65d39c243ea75854918b80957e999be10dd69e9cad588632beb4ab3983e15a46f04163860ddee43b64dadb311d2df0d4d59d4082f11ce5134bff2927a0888f01867fc680880b0129ebb06e99d96e7ac8b206a6b9420350402ca799ef435b0bda6e0a355c60e6a7e55dcd3205187b5aa17874173b61cf173c97a072c8b1232873265b5e1801773dfa9b9ab4720905edf69fb44ec1f3da1bbed207d342e01d47a276882d566991ab10c8464092840976b4d2f165d93021b3bcce7e09fb6eb0b6e40f872d584a930349e73a33001c7b8e96508662142d91d7f0ce1f90fa751d8c1e1f42eb2f5b47e6e984294cf61e537c7148bccfb17e80e1355144261556535c8c54b4673f9dc92190b1923ddbf24c987cca1c6ab5525cc03d0382e5bc131e58fd9495121f671038b9299ea5eeaa442af539d1c3552e72b96121589a6949d9d606a96a6b97f5e4cc4a3750c40a296b3abd8289ed4f7cb584eac0c4443de383d1bea46675dbd7237979e11abb7099329189b97978b68287b30436686a9bbed51bbeb45a373ed2380a296593b81cf79b601d9bee596a6ca681bbd36071c6cde71adf66fb8881b6e683f2711d5e6a6231d2c68205356df6c4ad71a7e82a8d7a7023ad15af1ab8551d967037c7f4f3402fd6e03843bff31c0ab3577cc300bcc77f921114d3d1b6fa734e14aa578463848d26664f86579f20cf1a38f453f17c4be641993b00a9afdd41bf92ff2909d6ee9123e494965c72003def51e5da180e7a1ce9db39937f97d803aacf438cb755e6c23af370a7b959261e2ac77f24c3074eec0d3457268bf4ea852b9b4624949723c56cd6d1ea227f91016a245d742077d6bf4dbc3ce86372a5f0359fc197d8f0e46c37a6dfe2f601ff0d452feb8917934ccf65a52d7e1629d76a7adba866f1892a1c3d372bc469982e20f52fec732e60500617a6cd87d66feaf96cac91567fb3f526f6877fed3d726e1dec9d9ea86c8de91fe1e49b54e25a980640d0c96d8f4cfb470a67b94dd96d4175eb2a9531ef6b9b58e4290e938b77ed6b5e391dc01ccc836713a7511373202ed7bbac8d88ec7d7aec497eba58ab6a933e4f11bfa18eeae49e8ba7e5d3bbde19f80abfc1445e4fea6a64fa9c9cdad4cff77504d37615011d9fd11e7efcd14c06299b58c51a84b36abb0eca63ff98bde17cab378caa027da68e78207de23ba801aad9ba146eacd8d7709c757d8798d48676c9bee10cbee39bece49907a0086deb86922ba0ecf53c73bfd07aa2da7780cda60fbc498ec36eb5e24caeeeb965b1097a23f769837074b98a2a3e939651543a517ea12d13b92fd13fce3914fe6b6806607baf1d298aa84aa62e92e7d25d0874c2cb6225066db2bdf8fc54b337c13e1363dd0904a143214c8e14dce0252161ef057768a4708e78861325c231fff0df3d442f19758672284b84201ea4630f8d8abe9d7627d99e015db9ec38e700d09fbeeedbe26ad812587fc3c1fbe81514824e018fb38077a275200a9e89c92b86cd77a7d83a0b6930a6ee00df4318f9f32cda81041221d3d78906ed6c4197bd09b2968e2f8af59333e8f66f85950404318882fac4e980a61f6333ded71e26ba06600e7337d3deaaa0fbbbd29d2dd73f53d60c2312999383fa03d0af2821d1e55b0bb550cf9059be81f6538579863952b3cf0f5522c1ac43cc6fc719d0320640c61f08ec0abd93c49eaf108d211acb3b62ff1f2766e66cc241dc0bdf7b9f91d659320c4b52522394768b655b362b1af0ed799f8f5e315ad73d138b5a1a078f73d1e141a29c02f495dc963248796ab4eab7d120f643a6e59d5ea4a5383199afc556755b3a613b78250a827b431079f6b3c51d33a6a8126113702a18060d1f3572d58dbd2f7eb0e59a9ae5efefd0d770d53bd390011312e0d3e8aa4edd11431d70b715c25927343aae5b347ea67a455caf533551e042a662bcd8386fa46eec704b3b1d744ff0db87eb066a971db809a1b3ec86550663824838875eef90703b6b4a87f5f3e8a1e5361ce1a380c79b4f4012ae2b74321c93d19c91944464c3ccecad057138f0b0ba81dfce7762c7d207a85d5c6a5c64458a34fe4df4df9e6fac66812d3ec11d896f1a89ae830ff69b9633a901ae2d5de6e4ac5d717ced47c0b1121e770ef8a4067024fd4443db2992acc92e0dba5ce4297196072ca7539d8c1996bc809596f0dd825c800590f85f00c393069cdf7f2171113e8e731ccec30c5d10cd12945fd198da4bb0bc56203b6a91f71d037d7307a2f22d0b8c713416d8f748211366d7a419d7d06f443a92f9feb3f21a59cf261fd82248fbd6c06967d14d391201c9e03aa055fcad356ce4ba93a66f54f072c717b96f87e64df15104be70af65c0473c241dcca44a502bc537a5377b91a106009d0b16a66c65c8be62dd7540abadb12504a0fe3a59b6b869fabc037ce77b914e9eada627556b17e9b94a4ea6e1a00ee6c4766196b79d505c1554c9cd97b7a3547cd27d4d538d7b92b30da19f8759cfa2f1ef0918ab0452d5d812ece426f777d837917af7329ea3006e36cf7b879ab31228b3010b39242108fbda8c98da1e4bc4033c7a5e7cef0a717da53c7fa00917a6827fb10f3e5a57de5e2d858d740e43b42625ba40168567c969ee34f3d614a5ba3e76b55b809b8388b0e46d434f3afde5851fffcc9d56f84f134267ebb966f671c64f49103a166d7246dd5bd74864cca8540ec98e0f6f70579192c072e3dcfc6d2853c4486281a15b7c3f0543dfe0244c1d1feb32a10f471e63eff1a4302779f6c1656098ac85b85a4e93ae6a49a338c9adf26407486abe27661661dcd9505c8efc8c57a6c6f0fe8555c0f6486abab3aa78280beaa2779d7144b3a638256f93c6f4f6cd16f651f586250797ccb24f11d789cbcfce3484986a859937f9d8bf7a0df915e55d0d4b2db333a6cc3a91a69298a4185e54608d949713af35130ee8544bb63a5a2445a27c97ca8a08dc620b41595c146ee2855520cc034456b67c2077f75fdcefc8a091477df1c71be45d5092afc46bdd6fb665357f1ad8ad20cebd2703804a841e6345cab32370aca0b140887ceceb0f72350ddc99aa191db4e27c44e30188517eeb8de05c6bd8474528fd9e4b18d0c944c545cafe5a1c8aa034cadfd6ab6e4b9ec1c580b1c997fc24b511a791f934320e011142099f32b0cec90db0caeed78c38a240b580f74a49dbbb93a870755b697eb65625046eab48e2a30dd17d189767689243cf13bea232310ab65c78542342804ed7ef28f2fcc58edc80de095fda81376243eac30d01e2db83f382a936991cecb06a966f9c52b25af1266521dc8e997b11619c63e22dc560008022c3db26184e158878fc51b3add6f6966800c8f2ca1b9c21a156c5f4cea061d82d714a5c07a05134fccdcfe1c2b5832926d8f2035c0a5df7c8a3a40ce2fb874bb50dd39fb787708a45c7f7be316a5d406b3cddaeb12b0cb59a24e7fc1520d1e7345a6023932426427eca9d1f93e20ad00512ebe05f3f38b262e0e21027eb7ecb9ab15e1f79eb2456fdf2393ee4e54dd978bc6fe7d87bd2bd4d84898a637578f7fa59b2359e5aa41bd2788f348c7d12af86be117e11655d4ef722fad1d4b66168a91ce3bc705333f06a52874caeb64036c0d8780252f97f2e0e9ff989dd292ef4b3cb0802be85d8b49ad30c1a714a269bbc1081acd25da9f873b1fdadcf19503436c6f7d63400e47498befe816317105ddb68db7ec5546da781ce48e7fe4aa26a4ecea70d0977fa1ceb83d5e9381eb230e04b4bb26da5819e19d3f112e842dfb84564fa7b7179c51079a3ae6c0f32342ea49d9083300776ad69664e653e819d2d8bab36aa2ac4703b67859d5dfa08d4d8bf9dd9524eb0cc1bd6071ec576d82875ab522b09fd6c616c664886a98bb4bc4e4d9ee7e7a807fcd5e752e410368b971d802b1fcfd9ce6f7d6ed0629f3b8b184cccc128a579bd98e9ccd42d06d3c43159e482798ba29491d22525855c41da1fb71172dcdd8a94023b6211793c6be699cc3fc5cf145965afa41517125365ee9463396ca1bb8ece9c5cb6a30a563c9d8f61b7643cde0637cb8c017466c7e8523f10da6fcadaaa97130d472c3b9e4c70a5080ee966cff580aaba39a716775636554158be91c5fc99add635e9d5c0a9a40356ef81595d9744f424c67b113d5bff0277457ef3bc0b8a9d5e87720d5c0c0d51ccc815c9da1d28cb790a64807953349aa27672454246235ed7a447f21b0edd927d2fd531e0cb0498eafde16f15885fde449482c561ede4ceb76d752a1a94e71a0e7ec40f50f1868d38a4c3a62d65c50e22390aeea4936a87853a3090915a566cfed310544e79d9cfac7f9dc432be4500b700fdcf93c0d7a8091af6b0d9ef6ce6afedab2b43520a55a785039bb34a0f397366b356b32641e45f98369f8eb7e2e4345db2e5a2f6414c5ad21009e5eafc848b5338b3bbf4c38fb541174bd395fab88ec468f018bf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc336782e4ca466eb0edf6f42fbbf931f6aa61cf9a984e8fc345cd9d439130ee8852c734b79370b64d2c3abbcc774b78536a126ef1052eb00d5fa51a97ad0fa8f70ad60dc35d88b2d1786c79af163f461c3a75bc18a1b430d394aae44d4cd64527796d7342e1011a2856e3b7e09037e180658f4e55c3fc5f5baf63fd173ec7a0dd35304513ded099b555f1ed568c74b9a7de268b49e1142b84039ec574a6bf2e661fd8d3f3f16ebd3bc0bbc91f5c6f6ffc53d2e35822915686efc047d8bca66c3a2924a086a2c527846f51eac69cad38b49fa75085f44560e7cabea41adf3716d2dd1d3b14d9c2a05c11f7cdfe38fd9b3c8830336e3777780e0e45c98d338d85b8b45975f781ff4709a9e044d5efbc0eaa5ebca5a4740e10e888831cf6a3a30f6eabb7634c8cedd6df892787c0dbb4f6e41b491a45a67ec3a9084633282ba48210677dce563511a3e46c3366ae1fb06ad631fd42b70746dd77d67bd47c970e2af271ee5f64bab0446dd11bd57539cb288b32c9edb0b0fe2471323e215a5497532e19a28765b64bbc227d72f079120f6533d7122df8148ce2a1b1e7eb43895642a36fa7decff6eec3c79a8ec1f17904756e9f93199baf17fa52fa02b93ff35e06bc00627bc6f2bf817758b4e190c7541c8707890984178295d7c4d3e8f9db24bed2537a8011ca8cc6b7826f230cc0aef00d0f129d655b921b09aa4aa569d866f2e222aa96f5caf370cae4da36439b1f1546be8f87d4ec901099aecea1ebdd562f6c6a8348851abbf39131c71eaa66081d2f0f903ea5d0363b8eb075a2cb2c764cc60b98d7d3826c1d5f3865ed3350da01263f4909b5ceae7402f6d85980ae75beef57edbfd5b29948ad3cdb90f5de9ddface39b925f3d99b6bbcee2dbb15dcebc925c58ec725884f6cb86be925219d89744ee2917da7cc199829accda29dda8eb653a0f79132566dfbc0a3df374df717b2c5a9fa21f57c7118cc819f02368f58c71ab2349820fe4aa7229bf6b64cf93168d442ba85fbf0e2f13563b17c03d67787cbf1f767e3a26e50ad2dc56e8307500fe2e856f6c3610efb9f0044a21c2247fe9a9a4cd37b38ee96ce185769cc0220e516cf89385d9a3fed14e7cbe09894462a6bf6a1bbc48caf9a6788813ed43fb5255a24d82abd253ff765bd149ec532e6496cb469db1a128334e088573c5d5731e835ecdda9e2374cb23e4a752b651cd5ccfb017a7434f4b4a2e6cbd6491c36097989354df9ed67adbe65979dd8b24f38356e0334235238bf17afcf830de3242c1597cb26e4a4fce0319cded9671b2b0de2c5f86717bc7e23f7834e0fea254ed1e3f3ac4345b314b5f6d540cb9de3aa0774614d3694de14a744641d4988548eef2f04bef7d743830283bbf2af04d795e6d041e1cdf634a3b0d0c32498cc30ae8e364e82a3fb7cdc90a5b466fb8a660e07b9c8cb41438acfe6a703c6daf745973ef7ac5a053c704e15d1e7bbe4a5c0c9f4f438fd663aed0b0a7ed9d7f8a27bbcfcb7131d42961e2394be8faeb6adfd2521715737e1e752fba4a8beac6dc60023560a0c04f4c1eee035d5011299839aa66b48fd4fba628eca4070eb2847f4add903d4a293d1a87f302b100301685ed9148961fa33cd0557556d9a66ec3c5cd86c1b0a816e9870615c9d2e7f13fbf9ebd284fc621b292b8cbdb02d39c0b7154bad11f3e800e9517021f3f0d5f71b9f25cabe328b8cf95c603450e91794addcd392fbacb56303511862d4c7bf07857a27c588be9c115e1cd8caaf3cf918a8fb2ee96339bbc8f7818e0220d06879b0d1cb686f15e811bc6f3fa2c745dcd620334dc92c2f25bb92e3ba9fbf48c694004937dc16794a06e6157b6f85c215e30bd4c6713414a6b766a0b91e6e3c043def41ae263e338c953f3a460fa5a1a78a5bd402daa4dbeb82059d4f382a2164c05ae52cdc26d222600e40ae744d1d7cdf6e83e9860960a7c7e82100f3ebb2b3cbf37c9ff5501474d64ebe0ec39662034fb85868449af79de29e80f07d688d08ce836004b05969aaa717075e379d642c6d459476c374e3e608bd6f9224a7924f6fcd88d7c76b97d5b6e86cf4626ea8982cca39b2b15f0cde94696da857072b8788dc4b7a62ab5a0f859f4b4b0e4a388ec2c077a882ed546c35e00802eceb88bcc461362a66e9545b7cb865914b7d44635ebd185d6f374ccb5380530a11179ef4ca8aeb45a9d739f59422efc07278cf34de11b245c2b9989ae1e533b60c5f8b453672b98de130303052e93a8d92ebfd71217211f133a34381d85ce932ac8881bb6f522208ec3988200bc47faacd859e579620620ca5cb5131fbd71d27e2f7b836d78c089fc3ab38eff6cf95ea28d83d58fae6715cf493164e100e09fcf6fe6841ffa0fddb11320a5870a6b8a8494eb8556df8b48586a5651e10f41ca841fbaf223e211b794b482a896ae28e41f05d8693602ec92c0808986ea05b88c7993a737bbbd4ab2c7dd191fb8dcf8661c257fdfc6c6accb27fd7b6ac34ffb7edd3e1f51daa02c377739748956c76b13bebab7e29839fc5936147254ddeb4d0e574d5dac1ca6ed0093c9fe17b95adc2dea3b89318c7fb8c3a954610b86f5b113ff6eade80c1cd188c8c30458f0b1c7c04a2f9f552c74dd3ef64d6a46088ea466762083028ccec7914cbde0799bd02c6afc47c50e398a962d2cfefae87449394897dc024f8e320dc1e6a53ed9990b1fe680fbbe692a6839a6341055542efc5048caf780a3abecdd8fcefebc2949f98a3c21f67a8e4156eadc5b0182d3bd1858f904a848f90448e030b31c082db228993191540bdece9b4b92635298bcd56fbdcae316c619b3c80c5b10a57b7f7e88540c187b941ce14edbe2410c5208eb4b3b5f8c2bc28adf2b55afe1d0c1780683237d03676d48420f9ed4482540339e640bad3f922980f1bbe5c652d097c894a12ca00501e377591b264033102d8b88e1a4e5c1a3ba2ba2afa2a4e7449ff33424c0dedaef8e6295471c06e4863bbc3db2720b40d73f60521710acdf8a6c450c9a79ab3265863e149c36e94459cac867f2dd61cefca2008eb6fece2138e04912e382d3303c06181512f312857125038369fde96e3dfd1a9c0a4a9127604695221bc16890b8c4185524766c2f01e643b6aab79cd5980ffe338a27ea31042f9c5c9891b996beaf96497bf335bc92a4bbf54cd47d13cdb8d51ac7dcc8db2ad230d70da06462f98d05bf2e46693688aff3eaa0d1e6f53cfe62ddb5515ea6ccafe10abe5067ec178cb3c847ff494258b809704fdf362c23a0a471207a4ddf0964b3c0597828297eb9d1530637391f177dd7d48b7d23baf4ca54e2cbd9993eec72564294b37e7f62ee0aff383bcd7f7dfe3a5d94faad0009fbebe7a00f57bdda3a35f2b02e416a3cef55728ff33b9809d80787b74dbdb92e0a12fb1eff5d9eb507e55256de81879d9c494c99d59dc08cb1a69763be4eccce9bcd74ea5f1c85f7398b77b9f9a5d117063d3ced641e80910ccad09d3961e3951abe2a3d33395be261143ba2d46744a4e76b535499fca425060a41a937cefdb20a0574e5b780c32c57f933391502d93df881c3f843619de76c56e5aa8a2a84cb3ade2ffe1d7c86a277edd3ef5091fe0dcdb9245958154d9fc8deb51c35fe76f8b143a54ff4ec83c6b972f3ec526cae32ad6d2352a1b8a113d972ee020bd53cca510bc96c557dce9f907e100a355e1d51fe6f6bdc4ee62de17b007a7c18816a17e62a4253ccdadbadddfb0e5ab36ee901b6fa26f3e99596256dcc68619a3193b89e6eed46f8c3dbfaf20bb4080247581040a6859e3798d1a6568244d6acfd7ac522b451cf49853f31732d8a6bfe66d6eabd30aa4b826216926bf48bdbb871178d782eaebdadf9a6a6fb7cb19adec547349bb133c8b9c0b9df3a42ad218410eb569737779a265816a3ddf9026d79674b08d7ff5ea1abede045312204d3138640116fd470f222e168a11438b92182266e772b329f14a2dacc5f064b0c8ef96da3a502f43dad66adf5eef214eeab417ea528880b6de94765b6392e7e161fd145c263b68f1cbab2cbfe9dbf2a9d8d55ae029cfb1a27cff6268159c0cc4378fc6c88d9e767d5af591b9cb7cd5efe9e8af14536b08eec4f95adcd1b11ced69c0c4a670bb3dda5bfd37f9c9895374470451301649acf68d5c3174ebbcfcd3da10402f3a9df6195e8dbce2afd5b0d7a9525afddb608a9ccea82bffaa68ecad9d57def942a58bec44798af9899c77b015443a601222dd10541342abc39df5a868e5b182498798896c2c4385956b94033ce5b3b147f2bc27111fe5091e73a2b08706d36926a57297dac57b05b7bf8b7f824e5a18ba90b710165d74e9ff8224cf1d5974b1285aa8739c9ad4f4daac9a34d83ebca24fcd1e6ccd113de0dc887a113fd61221182deb0bc465137bf170bec4b8b2ae9c2522c25663d19ed6c02e1d22a355f850a7101da61ae11f2a148ca7f6787ac6b76ee76779386b38c5030246c216e8c58a3bb36af7f0f207991ea4a3b94db2cf90f789db5c01e2cc2edc22e8a4e67958e1d097e72a40fefb2f3e7388806960acc05ef15cba533f72b99008feb9061245e8c1681b315d54a485f7a7c16ca591028010b263d7fef322d36de5d0dcfccff33858cae3fc00a752e18604e55f7b0f0e71f70ea820da82595ea61e0c7e91d5700ef36b3810f1ae1495b3cc2681c658424e88d1352df12a0d143e4936b06f7c2e85747bb4260a00298215463e57746e1605ed729ca30305e87af9f4febb284ec3d854cde6521b9501d7cef74f943164e2d6fe44ccee25b6e76eb79eddeb7e678dfaa3546d33da934e0f758576dee7456e7c6f91ae9c36d4bc98cf54315d97537f09c01e500f4555bbf6ea63ddf92fb993c26c51d445826b6d0b5210cfe1e1fcff76f5688ecd9a878509da1c504e16357e980babed214348a2891ea10c52d42c2422b494c09f4abf5211974a1f2369639fdc01964efb00e59839d9a8d0d1227d56cbfe25a57eb753f07ddadd7fd057831a31f7f97b72bec6baf524cd64edfa8a25dfce499cb4e056dcd0aad7e085e4cbc6cec9dba1a953c24412c9add8a31075f8bd5f0e8a5a2bebbf79997e5fff83025412f3d8717163f1d173f67257f4a36258e6ccae3d3e8c81a007bea5a82c1eee1f578a73e098710c0ae5eb71c346891be1684e973c256d40d95a5f2bf6a8dd8fe97131764f36b079cf879ce39261d484ad3e593e4891b9ecc40cbbd683d76fda2d96ec6330330d78564522363dfb436cac65d7345754fa12d8bc8eecfb43adf9e433bc19220c90d88e1510a9a287f94e813fdea92be47c364b199710391426cdf576d12ceb9194a4ff34b0a1cd8bdca115ad521c999783058b29a1f671d820f1fdc766a941d53c502c06dd18c4639dfa42b4a76261e64ff64aeb2dba15234576231d39cc2765e7486c550345a5049692dd2dc1146cbfc76a8e6e0a50eaaf6fb0a0e86ff317288cb2e782b672464705c51786f52157670d4c297d6684cf509a6f67b02ccafba3eb87f6b5ba5771f6d25785fa9b22e2be6a296e170652df0102ad1389007a4334bc21be2ecd15c658bef5f1559aaee94f5fdd1a548f838f1a4e04ca76101a1d075cf3c0a358147cf6885d03f322a1a10fa9658f66d76e3278c4404d7971944b478abeb91bcedee2d526e3ff54000ca90fbb7530f11d5891c07389d0a50087c06d04a9389265ca895948617c210e302d099d49b6a6b960b4aa05c98f3c2959d8865054f39b7fd6b489781d1e1c2f9538862537aeb5dc9b59;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha0514a5a7616b29ba248fdbe22e2346ea17a2b2a099d6b46b4c0f67e1792d7ed54c5d9b21851f6d8974749b94ae5b06c60152953da0c947b7df2a15e200199802d87b49d53d3c185e4815190780df8a046df51a191dcebe870bc700e8059815203785adc04d1c1aabb1926a8a553efb238f4b0afb9087b6911c75b34c06e3f97443cf1591df310ef169970dfaf9283b4d03b13df60fe91d60c22a2bcf004c27f5082fa30fd7ab13e2916e72c6d5c171481e1d13979a9f0b4c91d117432961a5ccf72fe02acbb5d417c4f93b7a69abd7e5e4611505bc170e09632e0ac646cafa18aadabf54d28e8d3329861233b8a0028dbc847bc5b91ebe065d17a6b1c316fdb8721fdb14fe19498cb37799e61cd85908a7f1aff660d9a982573e2a60bd690f62ffcb15d65cec7734ff19ac367d685bb00d8ee762936a423395240a84cbcf147ecae74b205dfb4e213270eee8125cee97abd257bbb3a9783c4f1bae8e7664a44505f8b20367537d023aa7fb473e5f99c1af07984786268dd7912a73cd014bb733cd052e98f5e21333cac0e5f671e5ee7b95135ec58699f47e11ce21094160844f176a34d25fac3c17f39491a9164c88953d78f09d9c204482b47e63ee781de51dc5b9e7166c2614a7db6d7b4a9f8ce65a16b7c226303d4e20ac1cd977d78522360cd61b942f85764554a8f23ccdac16a83b8cb6707a45547860bb7f6f8dd675f5bc8dcdf3a8bc75b08b31b125872f28cc1ee07432cf86516462e028882389f05e6a6fedb03968dc1dcdfb81fe3339609b534305fe162cb7cdcf4c4b0944781fe96f2a5ffc755a4c9008147d1239404c828401e4dafba5639b5b50cbaa97c493178cf0b1796ac4fc480d207cbcb8e554695540f22c229f27fbe7fc3be5fac380f5c724f92f1108edd487f0048f85ce6c86b780372f56b67bcf1375612ca64dce93989a5c59e0ffa6e732b3693cc41143c3321b909fbe236f84caa0daba687c6aa46449a74298f27dc912263bfcd17656fb1da6e999b4d57198304b1dd5ea04b5b535dbfd2a6aaef443612a877b35aa6f3b1d2e2ac2f3ecfd1c33cc029677620023a40479837d689143efa1dec3df9e5c3df1692b9d9c0a348b1d341c311223d253ddc335bd9d817b8db8d1c31727e1f2eb95182e167acaf2cf617a85dbd87bbd9fea425cee14e0d28528eda25829977f2fb9973e674c9f660e442eaa46c67cf9c58f0f0ba39701ebe9a68c8e993ce2fa2b182b71c268358c58b77685fdf4aeb228c42dd40575f7ff7a92b7029216eb06bacda1eda1127b77032175c8b25f0d2988e73f863020ab2a4fc08be401590865175c66ce61d0e0acbba7189caca5f0c6606dbaabedb768c6799366240c22e030b1ef1cca11669754b858e3c85846102062918aad97f5f1ad5b15c14b42c509253a98f02ba427c26a14c2343efded052dd849a9a26fd45ed3b9b42ae61f3358aaf407634558ca518d07c4a6288a3d2ef9f10390cd6371e096d7d5db78d6caee586c0184c146aa02df09e6ea84ebb44cde6f99ad673a781059ac49c3564f95c9faee65d86ef9dce450b705e712c3f5cfaf34b139ed83ce503e5a8227401e3cab4f73fd50f86384a4dd72ff7c6233c1e6b0ba20b85a73c9097868992faaff5513f63df1344c500f1315c3fd5b49c909ebf16356eb1018e504378f0858d247da2076e1248755563c8b17a53fe63a95572f2f395d0108a5127e2c7e3758eb6d46f14e134e7f0e2c8baa6e2ff110798df9ef74cba7491d132d53a712dcd04814cf534ff3d54d4ba8361d36e8b21a98d7fe4576fe95da8adfdd819e5412b66e08d9015795860aaefd6e79483a3d2f4d1e8989a16f9386601289f0df2b1d8c65720a8a2b497b84ee6cfed4ea7244f6800514aa45140d50a1bd17040d5278d02fe13dadb0dfa42e7fdca5d41db5dc9470bf26fdcb618660031c90660079e04c436b5d1598b87423e66a6b08eb39cbff71aca47051826fd046bcee988a834b114e62418520a0180bb667a761d3e97c0b90ad5b9b38ffa26015a86c07e850983cfe8c54b9b0bdae5fe91d15bad4e92fc992193774f3b577731b0f2a99cef2f592eda036f5d0afa324f270b35142c49bffdd6b7234ab563a17d5b6c237cc31bf27cadd70cc0d467b7ba873866515e4b2da07e34551636b0ecaceca82ab3b5a899552f1850436f193002ab9b65ec02cea692375659cdbb45530d46b816d9c921e9fcaa688b999e47a858ddb2f396a4cc66ac47099997bb071ff120f44458ed9511aa5f5942f9c1019320b85b60e59a973ae1fa09ab3eee9ec6a82fb66442a276a42520362bbe9ebc6c797daee471762a0a84b654dcc4541e143e432276b9d85bdff743e59e4e40d658086bfed9eac1aa3eea7d5e06694015d0c94e49db7908e2de4a28f6b8159d936ef8f6f58edd18aa566a07ce1429c1236f413fc9f5322e9def090e4573749f7dd00ba7a7c816dd2464904bb2340a872a0c9534a256b4762451784f2e6205de9c0c962a685ca8cc8cc99453a50668e8a5fc91a3bb9916a01f7adc5b176b736a4992ebd838fdd692c221bcd549688ecffe6594bf80afa11bce59ea50e718a6636491d47d2f0345300ccf661015c0c6660d70a8df97862f5b365ebd141392ae7834e6dc311e5b1b413b20bc4b892c13268adef9a6523968b9e7b912d876b5d93dd05e7c364cafd44f067f732c2453757f97a6f22c629a1d88a1777ed71b52350683317e144ee6455d15877575ba50534655cfb3fd93f8d6788200ee34f6dc4a2ac06ce3d209e6f6f0c5d301166f6e687a4fc98f1ded4e5a399711425546450a4428948702241ba7fcd42ebeab3491ec63ab71822520b695c08b6050bcf5d2377c680edbc4ec3173dbf02fde59531cad4ad7f3f9fe25cca2c123ce1a7015b340cdc268a8c22d73bc0bfc3e5e21230298ae2670f1372b76c690ccae036607c32060399c1adfac18f9b6bdd9e41cc6af00e172e45c0e68aecb2909289c52261256ee48ace5f30b0443444b1f4915334fc2e0d4a07b7f9d69b8a56c937bcf785bfd37455d03292eaae4b1564c5303458fae6d25f9f6d0b3c9b9c30479fff92b0e501159e2381e099b5426eeed95b0044caa0d561a30f90174e3ac884485a6594d7c364fc52b0de7fdd1218a76c69862c205eaa93dd1b1ee42450c3ac4b9f3b5407bbeb885768129d091009eb15f6d8b6089c237a30d8c05763fb639885d696054294ed82ccae8874d89ac194fc4b83e4e423eebdf3da7f6f5533b85bbb2cc0ae79e28a551a79e6bcef4c752129cec9a4f3d8dd939e93871ec960b01a8489a968c5d7b83fe094196be87c2d3c3b97488f17c1b43c9b9587e5f58e3e4691ac328ea41dd957ae15805772d09ed2eb1bb285e1ea32dcec6a694a3b22da462c99b3e5c5ba4eedbb5b32ca111f6cebb21ebcd996d1742fa1372d9851601b87eb156b0b30937d7de2d29df3cc6775d9e9e6803a790bcffd7c48e8d7ccd224ba7b05756da314369c8ee930b985fe5f097963bb221e2f5e4cbfe572b7a57f4427572bf5f1536e55814ca2bc3b88a3e2cba663948fc3fd297069f64d5e216b8e649520659522a9bf059bc64a3a7da4be510f84dd85b566f065c55ce9be7942826e73e33a1f785fff9fce07fd3832634f22e4fd6166621811b5f1559cbbe1e4f80d2eea47587d1169e3833cbbe38fd42f236e8e4dfe1c883a5137660dc6c2a1bd6eb542e2fed708f8e1f906471034cfd4b517c0ecc6348716340ed277f0a7932a590df5b61ff2d0102ec46ac9f5793d51dedfb1ca5fa5230fc0f3eac86dc471c16dcf6e372d59afea76e96d03cb364551b3fe4283ee3bd1d1d851ab5938038e1a51cdc7c720d1795ab034891a57fe725b0dc371c5bebe0665b111f066c2e5c6d77adb96d7c6388ba7132a34ffa053a2c568451ade22abe50eeab27a55280664fc6da9c14243d12c2a92aee79ea6e5bed05f349e8b534120a453ecb5207f1572aa2617de13eb9025066fff7aefeca3681e9ec292485f52116d63154490878805c71fce03f97b58323e43229e0b4e81aff51b45cc6a4475d82d5cbdad5d4b93f3371bec8f77c588315f816edb34d412ad54f2e9e18f686dc3c4780029da9d4f565648141a60d234c2490bb0511e46d6b56e22149d0669d0f8c12a3548672277a2250151ec1d8bd8f857c72e29ad40beec00d64f7de620b907b3f38d797d2de24eae536941e024cdb01debcff5b3ca237e4773d5d198d86c3b1c40fccee7cf1509482bdd9e9b71317f7b232f47a827de961c723355c0720701f3109ed490f5c1f363510f0f29db23a059b54225421b6677cd3483707f9da74c05679ef71099fd3541d3750e40711a497256659919593d2ce1e75edf03d257c2f2510795d23f3229f18f4df8f516226f0c98894a75a80679c51b6dc3614804fcae9cc4f1df269050391f3746c73939ee6288314db2ed52393ae0abe43edeaf04cc545c2e55361f5dbb27d2efafdfb0455e1eec9a609300db6e90ceae2988ffdd891aeddad26d6324d00f25d138eff57fbb484e29ab7d011a9f5628f2d182ca7294966d85a0985c419d274adbfd98632179c6d042aebb1f938272a310fe4a18de473717665eb647680cf20ac5634fd8345a785fa77d0d870a4245d0f6143a5c0c4842cda5f797cc11e518231a7f188431275d623a1c40f1194762d21118eda7c7f7f40f480f6d694f447ed8f7639c3b1f60a2e8a4167ae54c4d557a4e9a1f25aef670711571e9775678fdc0805b3d9c8ddad43c1a3974b63c86813867cd9f4a4aec870ee376c14b78a39c1ec38873ee9af2b4aa1ec7e7f876277003b05726bad3d91dc21896ae6544f3c7eb2207ead7ba9cf07f4d71ad7b56dd6b238da4b25e273b0b52a5a54231daf9f28c55e1ecb83d37a4f8913a0ceba91c95b6994f3071c4d98737cc8cf51cf5b357f2a364eee085e0abcd94ae65db81641fc1438f2d3ff913defa49e719d71cd6433e761874208e4c703f8af799a7bcce49d120b362e3201b533608abfb0444afac68b3c7d6a333c4c3177e3cb1cb7aab6ed86f7a2786c0df187a7dbe2e3544b9ebfc98f7cb57b406408ee135844462f642d578bf6c721184f0d1274586ce126453c1ee1a7bda01353022b5d154ea18b26ad8c27abb618779e19bfe08eba6417dd72686e3a9d23f84b2aa94f9072ead5161d2b7f17e6977ed30bef79b42db8f3331ca18da452a18fe9e75307f63242b62516c9aa8903047b1b54567922c90def807b9fdc5f3c989e8ffb8dc847e01ead61dc7be4d5d6642eac9dbbc18b84e9a13ff7fc4ada129e46c39f53c4ef94770d8028defb294cd110ce5330ecd80e9d56fe0e7e3d2e772edd6c88b13a95288a634e6e1f14566338df1abbb26e282317e5fc91da807992a0412e50c7c38e9017ba1b2faa5a80991a343212fdd6c3809a211a1a11609be63196cdd0fda5f1ef104c0bbd4622a392b58326e175f2d539094c6d5967ff2d6157fcde31bc93eb73743bf0b4bc6800f5e33605ffd1dc40726672f6e298e210e35c89d5bcbed699028154e7405760328e09343f218acd3739d09627f81f44d3b39373fe06ec642f29141ea54561bd15a7336e87b749f9dcb71e8e87f04d2ce322697750b792454ae33852ecd9ce4bce8ad0a2629f013be658f388b519b1638fa7425e44a2a3bf35761a6590fa25786f60fbd299dea6a6cc687c6b893ea9b443798bba31b3ac3f0a959d7082a9a59f3b477f0cc5c7fd3872f67f89f3adae3dcb597642507f74774879e67702c4f75c21c7e87e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h856420f74617f3afd71607baf043649f89ce016bfc3fbd79232f8d0d250655595624391928d7e8ae8675e461af9ccc2def6ed2db66252bf7d989a450ffd9268e0df9441a21d39d57bf3f31859654b32c5ec11cbe6cc5c0a04e6a78b2411e8302640803fb7e2104364688203048952d14c9499cae5debb40409ce37234207c10b91ab12c15cf6a4ebcbab0158f5109f571164e4d83862fd32a46f9fa138444543db3a8d03746b32fa2eccc14cab7db42c0edd0d6fc50428e029b1077e9155edd98ce521eea49758c1b46664d58bffb35a0df7d739cd9ee565e69f84a900abaea6b6f54dc881e950e25500be9c0766d4ac6f17ddff347a80b1fb78724e48d279104ce09ee1ec861a311447a4052a687d0b676dfd6ada92844798cb47cd9925666df621cb4388a578fc231aa4bafd452354631036dfa3b2be8730ee3d26390d5cede9745e4b08fe6c6ec5ffc21051dabd1d3d146ddf03d53ff98e2d4cdc62bd444f25c9af85c4f51489ab82249f8d57d137c2420644546d35285e58bf75f2e704eb6635a53b2239590b1128c5468ac0ca579ffdcacc0cfa3dae12cd8461b82daf92543d2aadb6932118fff5f5eed8908c39c9c56d2e42402fd8024e13d3a2405fe66da47d8eb7e931c4c52e1fe907126aca30aecef5ca38f9973d990ea8eacc50c280b9646d6d37a5f3a95c974212221fc5c6892f1930d4d0133e460f027e9ecdb210696f475af69ca642bef1ef1470bee31b8d3ebbf08778ccea85db9c0e199d094fa2425e4bb7d95c9835ff6fc482007727203e61125462f03c90da67691a1a7c5b726644adfe3550b5a1be68463cc867b4e0ad6c48629007d65b3071683b6fdb6594b20b397fb3ce771722e4f3faeda11e1249dc39332f5dd44977ff43095bf98c02ce123f12d1e456e70e6244ae0e706d7ae76075fdbdefaec72757b931f3a476018e36816d4d80e049c3b0691a59291b2fe8a82c23de81e9f4219e54aec326b4850551cf8406f8e303b70acd914e9da7a340f34ec608a4be88d1da9acf0e0fbfb36dc2d53e1e4cf1ef0c9ad254ce45da51bd70f129ad3476a463ed1d3f7e514377ff99973f07470032a0a40f0f8c1612ba5432757843fad963fc267d57b9331a04ce4fd713209d02ed8e5a1e00691a2dd13dba93bf87bb3cfce07a3ed780d29ea9d10aa4452dd14595ba4e6d14de9a138bf28426cbc452bec5d542c77c1256ef0ef03900ee4eec3ba6d44fac99492e1bbc52353f3a0bb59c8f5b64730b81818c30d829f1de5d19a6c46c3a879962a2fd8115080eda1034efbc7e65dffdf21cedb1b38fadd7f0b8e8b918ba0dd4fd33d5caee7d1cf387914c28ff728644701cce44874388c9fd0d83c381e2d33c6b1aaef3ea27241ac89d2fdea20e4c9c5b1eaac4a7b231b06d3f462fe26307d52d4d0a926d4756eab16671b599e18ff478f9b4199828b5db635ddf73b252cfc77b24dc7e243d72f7c71c3520f54669ef2fd4ca8f9771427e1a546cb3238c52fca2263d32db70a97b8e80f066fd6a6ca1f589ff6760bf3893ed13819159c327f3b4812005fdddcefb21ccc5975a658b17202042d89c7e53d85ca8d30457dec870ea59cb856af00f558d9c5443cbdea0474ef6d7d512005fe558b4eb03c2bb5d815c500fc670dc29cca1c845aef6097616ab24bb5fe630e44f28b57f1add25b86614f2e4542259fe69e5f7532a00111f14682772c2b2ab0bbae7e1ad1d37d3947d09b09aeaa01c97672273b255d0d693f65c33edde165bbd801d2f5e3dee13b47713b855bf50093c0496f4657bd864417df1d1137b9246f0bfed1ff1114789e04d34669ab1fb9ae606a6c0c000be923c42bae253ea1f482e5cfe6f586edc88466aba7a169e41c20620e378fb3b9a0ee37114d8e3f464920931cb8a00746c5d79d9f6ae59a398fd3b686a5d0e277c8f537b9fea354b04a3877cbb3d54353cb21c07bc02a04b8244668f5a654f25a3dea484bf2729a03ed3d6aef1c034079e10146b078dc633306210f94c1e081af4bd12138663c43f3f97243e556e4187bd4361f0234541e2cef2ae14e7546a1a381a8b89f4fcecbbb5fe4855f45295eeb56109c7a0ebf8cd566ea80bd33ada6b271bc0a454a8abe8df03f8ef7ad5aa8139f3f43b088f7b48b210b77baf4de6fef80f50d8716221b2c94742da0157f2dd6ca2b87f8d2e80e8e75a53da3e09037b088e6553a7aac908eda70da994b89686e803ef14a5e33c81098d6545b0567f7259dfce8113a3c6602174b30f55afb012c6cdc90c7311059a9cd62e4821e94e948364f09607731a3eeb3824eb1095d68d8dfe9cb0ba74f9d9cc5b4c8653f3debdaac28c471455b1473b16031a969f592fd5d45b68fc56078cb0ca32fbd5461a2c01d84616759143f203390a53629996bde29d3d579f66768c35cbc3a3288a5c9bd6f34bbc6dbd8e560d0819d483790b38f7c1c4232a86d67e6f2e96b12494cecc1e8176254e5aa0d3fdde744a20cac9c91b02ef27e5b1e39ccd3f88d92a08fa21ad49b79bbd7e85c5bc35d75319ed3d2a2d588c3e2e64c474ab8496cec33a2b8cc8a167def32878c923d93484c2e05b30ede848763ac9e125fc8d72cd23710cb3d0c669a4170ea1492eaa0f8ac91027c90ad1b3fb8c7a98565897ba7e7e9f2dacf145a95b1b6553ce84e273b4b643812fe38f6008ef25e5bb83b40f71ec7f8e0ff034afc30e9d684317fcc803b0fae5a9011447d07907a59f0c8c27bcf064d580c64c75947dcd8028e681af936a1836d505cc5d0e3c36ecf6eef393c29fa0ca9241608df24012822eb32b7ed82cfdd032f2d759f31ad96d6997d1104f8f2bf1fefcdb3321f9de817d29df2d15326f1876ab8ae8c538d48d7b136232565250b22d651e4f747efca5cf4422d2d9901827c7eef137b80d9e7d5b5a4450aba4dbc13c61c566c4ad8caeea9b2eb84355c2e9732646f226e1229caebeef7286932ae8dbaf0bc62101e9599ca454628ba6aed24e5be7bdc79a198899dd154052e90dd1bf7fa84ce69fad8b1bda035422fb997d115e6e743578a9fd3a80fe8d63d52663cf1159ac3f4f88454464cc8f6be455119787f2db8ba0943e7fbc1f36c8d82c68b533c035653bebaf130a35976711b7746826e0103a61efc29935e8797cb13e6cc371d45f2d7e28721eb47546caf2ff40dbaf044e1937489783d3a52620acf6aed76a079722d16352384e0dbb69df3cbb8749b4d0f9e8ac8c1f5de05ed5103355060a5323ea6b5b4eaf52073ec9a843f277391b793e5833155de30ca76754fa7a8eaf98b7971dffe7e2ab938b375c2ce77a416cba6f814b507e670f93d12ebdf48ace76ab6a28e802fd20277c5e514fde3da82ca44adde853a4f0f4ea7a568184dc2e776afeeb72b2f955f9a5704e004d9d87867c09462b69c3f6d9b9f3711655d8a76f12fc48ec566a6dbf4dcec14bba5c22f5505d255de0dedba9944e26d640862fd8a1c11ffbf339949878b0fc639db7ff3ea88029f99339f2b0fd075b461b52e1c549b47db9f6c88ca43793548ce67a82152c6adeffab9c2ecde82a0d9dc216451c6e540faba91ac9efd3986fc58c9de550c44e2a1a9b8b83ba64080a18edbc4229ac1a2b64ee182a77078fefc0ed30054d609f4e5ad6f3690aba9da2422f79801630a9c2bb9a6974b2b1df4c6ae65a16fff2f44cdfc1a04cc8a22346eca64be2082fe28d04eb618bb11b1b45e0744b533bc3bad3203a7538ff39978787d56b432cb39866cf4d8f3c5a466d0fcae97205dd201531f75400db0feee146f2f467f64f8507f494833d10bf25c3679e2221dcc215558996e58246755dabadca25c981d5ce9c10d41c645f0b1b4e5c7884636e7d96aa5e82e786544666b647961f9a994b89eca5ba9c4c3ae8fd6f6297604f4af539a6ba49d8bac2a725b4305eca5a178abfdb97b6d2c9cd126be504c8bc80e41dfc84c5d39ec027d1c148e9658d2a85bf5fdebf850fdba1991522ced178069cd049c4765847061581f6129fb471de4d9c32d80d806b516a63d00791946c2425b932d29b13bb200b8dcdcbf0c70a629e273fe44eed7670546834731b145f342aa67cfeefbd0de128ae6bafb92deed8a7a212b96eabc186f8d371ff4daad8693132a221762d049a64e9640a4d9cfd8d589d6086dc4ccdfc5ebb340c3849af220b592fa472bcbf1c2104ced72dedb7ac607729aed779eef0fa6c23b6c5583021003dcfc71b0a9055ecae1b6e14b93e228d01cd8d49659a4b4078afef193b9c90fd2d22c3464f2ff06e97a04f0a2a23c0462b5bedabf66297ea415e736ce96cae773c71068f3cdc3fd765dc1d321c4f0e70113139aa4a3810906197cfaa1159940c25c48aca9b94954b7bb1f4276fcc427c1cb3d57aaa7afcef197b58b4201d864d3ebb5f135d33ca95951eddcabc70e600e4086c3d5de35329c617ad2431f997f8e1d9427351020e0f69fc3a5af4cb973b6251d9fc4570eab8d63c988bed247f08550909fe033513660f9d48e9cd1b0cbfcaff20cf0d3ed17767316376bb8d94a287f9b653f77a7032cbbe86d09da8e209e9d8a699d6c376cb13209738d1b89dbb4e74fea76cce0586f3a966007036261a98f776fecc9ab7206e5a45d7a3e615aa895d20f65809271a196164dcac57e48751db3afe3418dacd54954b0bd5e1ddad68afc620c93e5b5d85a6ac3439f8b2a27db02fdcd6b91500b4cd0c9776e3aae323c54e282a93d97d70d38511b794b649df5af3dc2ab9ecb0f71b4458f2359da7747caeb63d2d7182a308b6d8d1c9a79d4a37c0c8fe76f79953c33774c9549e7638182db4e40169d61ad11888429b2c18c4859ab19acf3c84dd27ae6147e3b6cbb54c72b4df1906b879ee999fa197f34932ef384162867438754f09e3e6f67c6e7addda1d3530414696dbe180451eab6950051fb69d97db9be44976e14aecb82d230e4b7f1c72841d537c9d00d8f09480d1705bfe2d6a5f6e04887a5b952594640588fa4f2af5134e03e1f2da8be9b5f0532362550481727cc49fe3d018fef20f9478b7220840d004c8a1f6979ff5bf740958faf2396f9c7c1e34f4901015e2a74b41a1b86ec6e997cce8fdd7788ab50e4937a3b833a1d3d9a3b769effc2b4c9ae110c65e515dfeaa5cb9f3d92e2e740840477e5fd5ae1587a9925e3f836bc3f616f2f6c18e5575eb91a868c0e8be6541ef8b5d23dd77760c8b91d7b53761aaf6542de197b0c584bb5c45f11753f3b6af4046c8d4d5b35a20aed58094e8ab5bef94a50a0f26cb53278bb2fcdb1b8ceeb0f35cca0e228cef4344edbac6aadc8ad23cf3f01e3ed45ee655dc5368ec6b7847ec72bef7f275b0680ceb05b567f32f8ce8b5997a6ec9e89c097d14f12fb61d3916c2163fa2250e393c89121b21de03b588f740e45deb3eaccb7a8dfbaa7cb068d2e89d8976a065370ce550f23b2f8450a78b7ceca36e6304022889f7e233aa563b12142e50df737ed6fb9fb886dbe7efdba1c1c89e53b9192996398bd0fc10fb171669c0868621367a8140ada6a84086da35789eb69a0e3a870cb22a8b97c463c97c8d15320693cd5541f0d638e63940540bbe608c346b1c096c0b611829e4a08225ccd7a6bd0b12e50ddd7afc7c4d9e267180dc53dc3bcc714d79c47681e4c3aa6000f232635ce84ac02c11f80a28f6a97d2eac7a36b629d20ccbcfb0562af56716d867e619007a2c3cc11b838cfbd2aedaadbcfce25b14c419de2adb5597922cf509bdbb7f7c34067a040fd81389269f03962b17dc2df5bb6d58ce808c5cff959e8d24b1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3e32740dccdd0beeaf9d448ff81900fa60c711f732c27285a36a2fb7fcd0579942a323280103e86bf4a9a07249cf2c66bd7a83a0896f1a57b87d7ee8b390155c9074b8e4235c3766d866236d02bfa76fd8e0f0bd0e698c393253d16cce25712f35fa490387e394a5f46e551a6e1d5ae30c0a06cfb58631d9f9cd5d10d9b880abd108ae40caf752c29f2318c5028f8e8f91f60bcf32d642548f31320f26843a3998d2ae3d30a24c7d0bb36ec432d57ebd3fc2a31d686ff82c337db172657816c4741c7dc9838e344c8d709b59fa26a8cc27be71a71dac408055296eeefe7c2154bb65e033ce8fc0926c711bdb2d1f44270a24dbf35f7366b00751a2b1c68cbb79ef3757ae8fe00a1fd5e8fc5216c053b453e662c4c774fafebb773ad87593150f611370e6ca6daccf9dd011431f69fc5a152b94b3a6a627d65b8f7a912cc218469df5a16946418043864fb640cf3286f432b456af1b3ae7fa7565b59b34d2cd7969346ad396900cb81f108511cef1ea385aef312ce16bb0f1aa8da79b50f61cead50fc4ec481aa7253b912abe0cf944ae56a7367c5905ad600fc0c9445cec5490dba161dc8339565bb516b50a38a90e40448cecdf122e11a2beda1b4955f771794366100605437891cf7cb5dec85514c2f36c3e21f7dd4f721b87270b21084fa357d4a4e684275cc6ebf7bd8899454ca9ae2aa2963b0cb8a5c7b0e30f0ff8140b70c47cc1c2836bf9b0aa1dfe1e481ed75fbb433a8940296a92e8fd21121daa851bd0b415af086457b107c607f70e5e0466743a4dc3830f6c6cf5ea68c88b8a350b8eac6625ebbd7ce895d36cecffca71f9f77231e0a7c1b8a08cae9bee23ad8e83bdf1d18c2edec30e5a3991593f7432077265a2eb755b3110d7975c44170718f96c8752a75c99e66a1cc9c248a1ad88121039f57ee362446ef30df883d5aaa19de198aa945d4551b1bbecc19b611d033157a027eeb61dc2df6b6b2e35bce73b2d6303339d834ac70f6cfc1ce83c3d073e6c1cdb6b3c99a45a9a7ec97fcd31149d1af0b9922d4709bc503803fcaae8e27f0e124e30a4ca4bde606ff68316aa669a0962038bf9e2db313dec337ee7f3eb049c1bc906a46eb5966e5468b95474f3099640537b203ddac4480b20d0e1fd2e4977ec30d1f531ef442e4dd1377ac6aa1bbf247d04d7c3a1e454ab26c231fb83971ba9a0c194e496c2904e73477e13b1a4e18db8d813c10d0d138b5552abe8bf57852e82df1c1ae7ef696593ebe76b9df0a037df42661a6fbeba99f81d3ded2e2da6c0833d27079b3657f9bcaf0a0947e17832e776bc9a6d5e1d1570a42daae56520488fc97b62df78ffa3dc0931e01897cb596ab8d77bc74aa53ae7efc63508a994d36a928f93a74fe8cf744185c347e1fca4fb3bf3672d309b9345316a6e88af693ace9f9bc912fa0c61b9efde24974c0d10057a778cc775771be36031b0227953a370e887467d2e4272d24a0be6d6a0f5c98a6bf74956d1c1eef2d5a28008e6a8fc13d7b98d4bd314b709f7d5006b258e202a9dfb1c6bf9237c1885758ff1ca21e2e17069030c71ab5a7344fb1c2cd45f7cc1e145448ef7b0c0bfec56eb6c334c65cc990756fac60ffa73873243b03e83ebc1c0b7caed760f36f61c73111fc8d65e62f750308bd697ecb5a84c1a31584e3ccd17e8fad233a45ee95dc32eede9df3c7849e5dc00dafd9fc22b0f39cc429622e0bc875f4f499a85693fb94d88aad0a769bf6467f1e0249203b309ecf01ecd38f1c7eeba7f832b57843107de1d8656844f217b04778ed9bf69fa142aacf9931c4dbe00e876902be5383380927f5495920d51a830a50425bd411f39a7c92a9d4d17995411578c0488891ddf9b8a54b0602ae12a6055dbe0e9d6d9a392f93055aafd22ad5538be98eee7a78d12c7047813f96b2805f55d1a2c247601ee05befb9b10fab86ee2afe17305e0211c226d45b5467c2fb9dad3c3ee9b7401f04cca0d286312f945b1f35ce327575ce4f02d70bd36dc3ec10732a9b020475b28b490dc23c038446f18bbc59d028c504ffc6e7b3ac6830957be8c0fdf345831952f6cde7d0593dc9160e4bb27bd39989832e857c99473a146b553bae5d05b914374258f24766564a8a7009c61882586c4ce8ab8d0129dfeb2cbd314ce5276244096da90efe2a0c4a4eb572cdbb45ff065a2b823dfcf839085f8d12c2657b6f02ceb35704e1b3013770c00e5933a7373868d92ab99529aadbec1f759d687c6d0c29b2b47a06d5dacef1342a053205af0028e854db9abfd4e6a9efb897c14763657c9324d5deda479ac6034f4b4fef458cc3ef0ade447573d978ce9fe3a9e59604d68a84384dc6ced2d5bb96ca3e1eb17018c86580d2406eb71ef8b049a2c500cdb37d6db54f93cbd677947dbede260e900801456835e389f9cc87fe477ed46c1af882ea2a61773da2e45d21a28d02be48db5ab51fa05e08918e8e90f5c82dfadf03fdeb97207c3e9adae92332b81794b166cceb4b5570ee19b8d821a9b85e820536973f9bb8b5900e3b53ed2bba03a9845ac0df7adf4ff3875c84d4da541014af2f30d8b5e3387ef74a7096b1d6a5a21e21b84c0f68c48663e83e76fcebbb5b24fc18a3c8122b973e8b53e0201e48dd04b39efd001dbe53c78b96e87e9fea03db544b674a207c036b8f926ffa131f634c28ea6952e2557a93eeef70bcaf9a573e01610c17d1f5966eeb9a2abadf76d3320eab4f449dd0a1b2036fbbe1b93b33ba37f882e5e8ead40093727852e1d079b6f64176cd144d48b8ddf12363a4cb250dc6f30b6f6aa9cc724a9331ab6f017a9fcbc1f239b4e79b367f99766ba696c6c6881a51fe56799f2e7e0e5e67471d67276da382b167c40d4ff24a8c52deaa6df0febfe1daa90fedac8002118002b6529bc6c0ee9cc0a8144feaf0d3a0232713a0cb7a2b7f7b1618a1f5f93abcf89b2cdcfe76cf58510fac32b307ed41ed9af604c54de01ec3f838de97abc28ba9a6336e62aefd14d552b399e6b45ff2f7d9b5a31138526382b653c0b7cc7188943859f903fb68c0f6aeced0f9686a10495df5e2e566c985c24c1bb76e840ab20ea1934338181a5e2d82393116a16928ab2db62ea51ed1fa67e0545352e5dc6c2e860eb33657b5dcfbae8e4563b2247b85574b9df561b7c31ec725693beb63f3b44cff9031a304f9db9392e74dbfa11de03da8de9fffdc93272b5189207bb759e563dcd66e687a8e3d29bbc9a6f38b1fcdad24e8c79f42cdab3014aaaf6980f5343903681c0da619fd20056aa3c6498b3c31b5abc07a75e68cbcdbf24242f3875c43e79eded332b0d3078e12ba525cde99a2c4a6f400fb589328df7c01cc93686a5dcd9ac5f8053d3021dcad3234064c0252f8efbeff505f7c662319d3f8f194372edfaff0d83060ddf881db7d24996a4f1f5924b4138fcf87179020dce936585d57fa1375d97877bc86b3bbd07662798e0770ccad7ea347d3049525333dfa6c16db930c595eba486417a2a7fe2c01453011be8a6a81ab23058e4b92fc8945de13c776888dd770c7c5aa66303476703f467d2845def979cddadfd7dfd6c03c4960ea69c1ef359fb6c4541d09bff8478f0f24f925476dc2c6364b4f3195d2837d58284eb4a6fab0fcc1f691eb806cf0eaadbaa9a4cf8b15ace56d02f48e116786322dd742b868f1ca63ad76e0dba2d86f38473f933b5b6c34c87a3c87fd1e546de1fe75e0f898a864d1ec527be8a6442b2374cefe3fa6eea9bf0023ac30690f307b4c45a8362b59dc11ab1b2fa8edc5b0591c685cfe457195e4a32d5d1930017f8bd7af0ae895e3eb2f50d52f6a2f7e5624890f00a1ae7d9272b7e9087dd367594bda9b83d711929a550171c978d41f978a15c5fe0456078237e041019f90b4c6f691c3973a2b68997d9b2743055541729c020c972de30abe71db8b2f7229db4fb97337bbb325fbd36095abf558480ceb2534b288b3dc58f606cccddf7c1c7cd5e05322b086b391ea33967d37e6b9755c852f0e2d8af689bc1aa11cfe18b49da43413b7fb031d634819ac9b30e6208dc936f4e7afdfeed47b75477a20d43c3327ceeded88180f172b76dde5f7e7a66840975a48694212f801fc60c69d3badb30ab5761252080f5e078683182b639998cce7b7f28133ca4a3be775bf71e00b1fd45877c2506f7f730790814bb27f0aa9a0c1f3084fc4080895f92e737b917a0083937bd95d4572c75d011f32890011b891769fcf34f9219416f36b7617a60f3793cc17c51156b91f074e6ae8cab94e72473aaf93e684e874eb54975a07e0f29a0a69b72de4d420ce40ac4bcb307bb3a45c3187c7b5caf14ee89b4a8195caf517d07ac362785a372f256a730b620a16287def3f9557564af8f26992c580463e8ae826d104c975093e5ff2c76f0115b12d2b563ac4c0dae7afc6fd20d4755f07823fdf156f64ff1a19c6e11315ffddcfb55bc6876d2553374a71cd4445b820ea96f014f1ec6600b058228d548b7d3b48c05a8b932598eb66c672aa7e1cc0574e3c72a9facb499a4412325e338d426042577071553320ae33a3f9353498f68cb76311ade52b3e3c5f1f04720e730ef51be3cb8bd32e3583b3f52a6689961af0af9bbcf03586b67ae4228dfadc83620473369f3bea145765a9855b5a77003143bf88e1d34d14b066a35e497308f501687d170db8a8a7ad0b0897ba4461c071b721de0f5f7fa3e1b6aa205503528a6ad3ce0bba2fbde3fd4f333ec9c1d3d136c9e237494706308bec63a5bcb3c83efcf0225b8d01c36bcf5d4777ecdb33d31a7ec753656ab8036991a74ceb5b42b66da20d1c11d09ea89ec77dbb6ec90e15e8d8df5193d4938bd61691144a91a90c1bb37cbe4b90b0f0518f90541e47830e904d8fcf564f09291cfbe3f7f87710a41b3f61a7f3adc2e95ac39502819a81534ed111d4b4501813bcaf2a56f5ded8dffb6cb49779fa6301cdd47672d4ebf71a25ef51d194f630497169dc2290b2bd023405107e66d3b84eeedc3787320f5432a2fb5050e541210962ca162bbdd78bef77f15ee879c701a765eb02c5757b2157750c417ed1c51c2ce67463508fa3d53771a56e4c3c0174d1a96669683a6e1797d1b4951d67aa3c7170fd1a4ba2965e39c02ea880304b0f4711f0002981ac7f43ddd98f858eb692a053a4f7d5d78503f14798c245f7e1491ee5efd133d24d6ff7d53cc5f69742b238cc8e55a399c9058c0377922a55e162ce0536f836666470defcdbdc4a8a9e277fe525de53db2c8decdfec1f680ff4f39af085f248ef12bdaf9b1ea19a909a8cd4cf37775482004c2be3e0e5871555cd62d18521b2bacd69bda4c9d50e83ea98699d4f7a95dabbb4d13b02a533306629556978b0ef92460223c6e09393f8cafd8de41d87494ebfc2fac2a6042072eb4490136d9c9ba708e35dd2b5402ab946db5318d3af74ca22cb3d387b295f6a9e077107f20c2c6074aaf531a2e49de04dc47de450d792d160b150bcccfcae66933419fc73d57d1047e5e4bc6b29eca5236c93973aae64224ab7ccd09b17179999d90d80c2d1acbd74781534609b058d6078e9fc0a0a268934e1e01083f3e434815b8526cb108ca8e30b6e17abddff0d32c06c96c3a7aa0868e7abefe3413644e10107ed7c0ba81f7e121799a2baf79053a5c8d0790813a1d3b36d14607b4d22580d066c7ec7445cb7692bb26d10daa35173a0f7336ffa9dba865852784e7ace65edffffcc3d2dc78e4a98646259dd8674e6c9c8af24ab2b6021867cef618d90baca8030de4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h94c877faf08ce90628b8ae87cf32fe0589bf156fee687d54bc97eca5d021351c50d990823b30372fa86462648e316101d9a7dff60d3e62669ec8e51453bd874a940ca8b2e12858ec12867b1eeed98f34eaacab40fa5760cb355ee5aadadaba91da97ad2fcd38cfd9604ba99dac68587c6836a45d9a660a0db4252bc877133cb3c59804f0b98c6da2636fa07453281fbf8b819fa97f790a9eeee777b6f6202bdffcbe91fb1c63042abc573e98ec088e461defab1c297c21be2d127e6713f55cab8eb516352149588da3329edb9d4ade04347610817512328ae0e5f11cbcca6469c6da7c0507d9a2a5ddf4d8fabbd9b3142756dd7fedbed64e9638fbc998951afd14e0d9cb09effbef5c5abce3a9d96294882451f11a10323274bdbd0e9e045c7362bda9230e2a39a5abf7350a18ce1ded73769d72dd087e3083a4c59017f503b86a88e2de415f4fd53c4b08b76b9b4e561ed60b1b4bdf7fe81894492602592e4de06888fb3334166682a19815c50c7ef768597a7963b6dfc635f3fa9117344b44682e6a8b39d8d468bef7d5b2cd9b0ac533b5ba96d0cde172a4aec02287c52a5facda89e814c919eed2aa877eda0330cb0fb54c5a426a8ac6fe91bce7093ad5eafad65f23181c078a7c472bfd851ab1ab071290062d0926f22cae711bfb011b839b0db5529dd77c789db09b607e956164a62c02b583796c90f1333d66f01ce8c7a4d8d714ad761cca3e31a0ee4e458a66580b3625bb286de0ad56d79cb1463b635561d7eb54a299cb8319c06f5317c52d94322be3e8d39beecd09384c4b89128ea947fae0de75e918c20dae1b2ab791cdee1a24af24084568908651cc51c83f803681a458f3dd342252eeb0587472034460fe61280894dbd55aa98006e9ee8fa3a5e17f1a8652793eba05f82e22b958e279dabac5c590a25ba4a09a559681af6695f97709306d3138c9d0f7adeaf9271a6c18aba2da79c69d74a5889a9e0838169d91ffd38a48a11155233146f0af50e77bf29fec66fa08b9afca783a9dcce7e010eb76cc12593f85d981e8cbaa8c7e7abca1a602d399cd96376f9d293cad3740cd5243df8e7ec151c1cd14ea629f5d6b2364b3fbbbd0ea5e163ff95278a1828bc0455fd31c1ac123c90b3b971f3875ecd58d3bbae580ab35cfc715383400c9c856761c68be74d97d4188eab8a006641ac1e962e99b48b53ec9ca1a58ff7db50af9365d76ea9633caa606d71646e9b0dadc7db2b709c07b44eca5975cb6f42ad9b875df95929253a61d659b39f753751b73e0c052cf5b5dece7f123652f8ff886f1fe31a7ffcaaa5e61685858eaf9ed7371e961d95f286f2a4a2beedc065881b4388ee7c6320e2d4a29fc26d3662a220395d9253cf9d3187265797fdd40a97af59638df5c3d6e9a67b705677142a4e643c142387e650bb9c4cbe5573ff46b1fb96d252cafc5cf4692ed041e335953f4328f006ede64d72afb6d23d2bbc226879f84918186c6aa6cf5f3b835a7a4358505a1a9cfb24e0404134ea158048ebd66571e1813550c901c7f95fd6ad0c4562c830b1b4e031aaf9303a9083389f027db1afe76f2b42b4c290567459c8d0d925bf1f08cea53f1a62b2e074c71b9b35c8d9db1efc63e49a459238a122b8f952eae26f1f46568df1140b454df98438f5541cfe989859d5565ed93fe3f465ff7ba2a3c1b3017f7cea8c09b90122c8dc1171dcf954e5f5abfcca8834ce0905025ba09d88d6824f59bdd5722f7181165735a8fbcca37efe7c9a73d001088df26ec00166d3f2b9b825992025e982f3f5231844c207ffdee432d9c2313a7906e43ec014ebbdbccb4bb9fdd309a05cd68890faa253f213c26743f721d1de3d4abdac480cef584398ad1181d8f90db5b519723cef1d0bdb76ef7ddffb30030329f51828c13a28f554079f7ea84f716a1c97c66bbf830b37720414377ad08bcede940cb90c24b2a6ee0d70f84a13f5054cfdcf1965c152eaf87b395ba474975494ff644550fee8cc022033116d97a054b746857549d5d5bf7ea5c96bed2485145d4e81180160a17f1cc568fcae39ed9c9b806fcad936d7e0b7285a9e01bce2810dfeb347f57287df30b1bf33f95d86b54b67eac2fc23135375914e63adbac2014371441e920c098c0485c09729ed488973b3c24282c39a17c45169ec84ede99778875e527247d701af35d079699081a86a317c00b1bf2a6f69d4e1398efdc1ea1ebb9eb3eedfc72eb5b4c390f364e755194385b981ec1665f89d43dc459a9d9e20d953026ac735245523164197d6bd2bd7dd4818449b0e3ce0a6d0a4c60d876df8d348fce946f97c5d71bbc52355860ad6afd9e1c57ba5d1d5adcf7883551317b6b25a483f5c8c8729898ff1adbdd3f980a87411271ff1ead5db527169c6302f01b6cd2cd2b45f0468b0f0c3c0003cb83fed3460bc067b972dae9184bee05732bbb807cadce7510919931f8ac6e401c840d6bfdb162422ce8846ace882cd0c74e98432590a743525e5cdf3990766da159a82e422877e1d36154f726051dd739339b93fea7d79958404d305539bc7e526bca484e36aa5dbda332ce59901add7e94ffa077235b6987b9dc96a50405caba5dc20d97c898d6663677a9a06c4c26d94fe096f8df8cbe73eec413be6a234cc9007601ffadc40cdc8f23a1850cb4c56e1cd811c321229161ae3c56d61d439a9b2e0dad3a45c555edfaec5404288c72f440be54114313f1c47ebce9476be5e46089e659b4af0246259452247f041e462d4deac597748af46a3026c8ae4abe66d98d830223fd1c489e5bfea971d6500fe40e3d519dee7d06368f9eb3e284c8305f820a9b7e13de721ab38351f4ef4a68cfbf1d06a0a1d66a21c8fb67f2cc029f9e8d37c31a6b2e0e17bc4002bf2f9ee696d07f053b51f0c7072a9c815eafc59ecfe696c2f21e3168071055fba8040a20235b5c2934d0feaa9d3eeba47a9b2b727604244148b706703381aa4000502fd535110ecac481846f3ae723cd347a87f8f10741a98a754beea1665a8dc8cbb7e6379f2bb8f3dc07003680a6f6c9b13ac3e32411eb0e519849b24379d4d632dc42b32ba8f78bd17b2dee6bd09f2e631cf5881bb5d22f24c2d7665ee6f4da53a55e17bcade97a6092a5f7263610a9637ec4d047010b920106c82eab44065c45268b30d16a7f097de69792f73a4f8b150a09283ed949b90fc5f7870693d7b57e669d9aab826e356772398f15366dc1ade21aa1ddd67d86691c2b7ccb36b0c980afccbd34dfe5b7ff3862f32c32f29656e3bdc71abb12ec2654b38d12f3975be2434aed773e6b032579ae368e1d8c1f3a4509faf896c76e973b7c80eae0d3054962c8a9b69a29f8f66a3e69239e35c886b07d19856960a3a33dd429a1ea461bdce9a030d845f6dc960b816350e797b4edafaf84c52b1a09032f7e5219e15d21afd6ee7b3f718b2e451be98835b47956d7ba18e5c69ae4dffb16482f8e386f84e63c77b5bd4bc92d388a409a1809e8f96d5b261ec4c4483103d8dca7f152f1cbb2d7d948348fbe0eb56a679e3ea32239a28ab14080808dac8c74d11611ae175ad30d1c956860ff94e5acd18d2dfa521c332a53a92bddd970922bc6828e097be5d1d0156d265dd9cf2bf523bf108dcf84949b26fdcec24e3da5d63b20babb4ff8fbf63f38f9e06d003d4a68da73116bd1b4f62dd9fabf74ca836dc14ec2550ee3f1cf3e3c150809f13790612ea782ec677d086c9e9d6088f00ae1ba32584c51069bf50a3acc78f1ab4be2ec7ffe539b678fd600b4d87bc4134f3ddc49195361d7732a30e879e224164dfb8d996b809493f1821a77d9027907716a0290fb0eea8462738b18035510722017c919110b1ecb06f2493bb836c9d43163235920355931e4d760bf5b367bfee0fe7ca2bff73d5c89aee7e0837df626651f250e0445a98a9939abc4dda70b01d09aac6f22863e3adb20b7db04f609e91b01d261f20126791882a64d03137503ba9c75dbd6c40c8038ca5b1f59b7e9443ec104b01e3153b0661504896985939f732e1288705cb3a9a0ef49ca460acd4c33c169576af7f7c523890dee3042bf86c6c9fe779d91926522454adf1464d4058953675057f99247dca67181798b59a9d3d7dd8f4e354cea840c58f07faf7fcb81e75cc732548e14281cdb50ae15d85a89cd88ba6727d2dc27d9c3a3e5d608ade3b417b474ed8cd52eda6e7e0c3e808a3afe93d6efe7962049249aa7082698e4a7a19bb748e01bed0575e83c42fc18b651574b7b156ad3da7969d1729db830baa8b58a67c939739ae145214da43451fc7430dd2b69cae134fec0ce7ff5b7fbf523aa44a45f5ed37b8e7a7c396c2a4c50cd6b15f20bdcf7fae35aa754993c7279640d4fd925a1a9cc21cbcd16b9a9be39e89632cb39623d7f1043573462ca790279a7a0fc25216a7797a072064510e43725d04f02e487213b451ecd9111d978523c3d953f5bc8ee309b270f4759f04650040514f67cbd1fd8aa38efcd7c82adc835e90574cd34f421e66b3eedd2439bf64dad110c733e3df6093e976526a9e810e687fe03a5ea1bc321da067eb8d8b01f89664d0254615070f88eafab4fe7e03715b6030506dbd5bbad2def9fd28fae5661b92b1358ea2c06bc28593c35f2eb3587be9b27f133180b152d64ded3da171da2e2825b903b24cc4374acc424748ce379a288de6a9170781e19f791271a79f6281bf03bbfec841e4b5231b1c6abfb3bb2efc732022dced080c08ec74c6be392fec1abe9dc93c06204a8d483e65d1d795ff63432d276710c8c390210a9b110dcc6874437dc72cf4f617c8b99666099668115c09f6145e22287bba0fafa9b10cc26d2142628e4020cb6bbe822b8c66017aedb33d58605b12aa553cfa86c1d0a6645c74a963fa315171b624d1e20ff8826cdd3a5e931d9cf7c884f786f1d28df9aa628ef428a577b75e57684a2426bccbd6eacd5dd9150cbe183d2798d8be1ca99ec111c0e78d98087e8a201277547ce05a776ed32da55018d9a408e8d1b9b0659b078208380f728181fb8393f68268ee4116dcabee5fcaef8897adf1b830da88d70e929d45fa72ff8b67b9c98982c4041b7fea880dbc23136730b7c2d49882aae1c555c9ddd4bb1b0456d1e72b7905b8a8d3b1c4bc93f71b375a020b2a6228454ce4646dabcbb311c038caa4cb81f65dd812d3049e5b828035c985e885a6c320b086a8fe971e3eca04b4d9140784c97a13e97d087277540947abc0239f7cdd2cd4236e8bc01cb119b4587be5e7fccf5d898810f9012b46922fd846879c2ddeece703db655aced970a99f0092057f8ed22f9b97442c804c2c1b85bfa033c4c83c47596a275cea47c251dcda693bb6ac9933c01d00a534b36995ef9a32111d6da090461fd82b7175a99f6d04a1d67518962b300898a6a7d12ef183e763e706f80e84e51b122e1e61c4bf90e53fbdd8dd1d4ab49405e8eddcbe93d7b485df948a64f70a6b44d343e67d53c5804e9aea049a69678bc4406d3bcb180eeea70b2fce06324ccdb3640eec95ed9bd34b81d8f7b78b3d7a028590d0718b178d021b48c58197f27383c800fabfe7b0e42bec776271c2d169119ca45f7fc4dc06640752b627789a747ffe0140b8b0c5dba7d26c72f5cbebf54feb787fd3ce01621181f01b72b63bdee5ad37480b83939b75c4b13efc171182d9c93c11437376c559467795b72ec8b723e76dbcdea1ad0e4489db919836432239ba29d53ef2222821a4986151e8f4b77b10bc95118d96416f15d87fee5cea0f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h517f8b122bbf1251a3e5c1e09dbae4c37bde2a9b2956d021e32b28b52e0b2d43ef85ba155a634d7a195484a81e06b947ff6b78833d6a2aef5ce45ee67d5e0a1d3e7b96cfc1030d7b7702312bb3b4ad651824d56c658c203c5bbad9525b67f33bb8ccb13229e87a27b0d90b4566032ea1c78910d650b9529523302268b7aef2ce6c4cd3eaafb43ab3aa274ebac92554d95a91a50b130fb6f1efa038201a864bb21a746be21bbfa4ac41b8875160a9533f8bb9e0d238c0d6d148170d8e84f33b11890f9dce11d941774e1df887049d5ab3a890cb3df180f244a660a9ca526bfcb602a7d1fea1ea6b9937d7f86b96f75e50fdc8d3a2aa42e346630a5f2ba5e7e35310048aa65bdea6ad8d0d01a9bcdadc1e98ed4c16fae5b74a0739016500d2b9e360bb0ac49299ce8302cd14c641ee5096d5e6125e25a0c7d0d0ef6f73e144a00dd165133a17186eea975283d14b93900c6df78468125c8738fd4b9089e01b3cfa9ca42281ccca6da6a64910e485593e88838cf6ba3cfec9b32b26b9e8eaa49ea715837b8597a806b00b64303242663346fa3023f8af74e2563b29ee96960ba69b79fd5cf7434432b79c72f05a0cf069ca32a39c1feddc1dfbda24296e390ebb908a46c06600a303e780b4d9bcf15e410aa9cefafbb7ee92e81997de4b5e9ff155598a4e0147c764382625ea07ce9bd4c4812462a2f2137939dcf2e237797311036dacf0137b6c62caf3488f9707b085274dcb6ea3a65ba74bfb7b0666e4401ccb57e39541e4b452f263012741934af79e6df66b8f853ad98737e6513c46f1545fcc81beedf1f5f1930860c749af6846493d72bbc3b079b51ddf5fe90e3d87e28ac0bffc55b1f8af496d801b3d64231457a5314dee4df32bda7a5e9a45cf35e0b2162cb448b76bdcb780f3e8fbc15ef1bc14d90d030b80f260f617f286002026d9739158fb99dff769463f6fb2ac633f1efbcf342646de65428b18adf0f6404a4ab0fd63fb6990699c6279d9177c8f635d48e53f877299ac16d277fc73e6708e64096bb9bc4a6fc841a78446dc536f93102ba03114fd21d056df0d6409d884acb4beaef688c59deaa592b5778266557efcca08e4973dc93fc4a20ac26ab7447b2afad13a52ba04f0c5cc738bf3be087ab553e30b31fbdb1d584220855a613db1ddef97430791defcaab8820aaf0d07039217e2312253f50191f4c2984a3c7d6267d0a7c0142d044e61cc428b43a9d9b66fc2830024f60756306a2f18b91a1c8d17b1b2df668294464e866245e572017dd9e60965ceb82d0c928d5e8e89146ff4fb34288e793ff9bb8a52139efbc4b7376a71f5c8c6b7b7583734c7649ec8fb677e2bac074cd24cf9bafa7fe4d6afc98ca72608c07f9ef9d7c621c3f74b1776821e729a0df8d93b3563e4fbe696ffb7bb89b84f87549412ce0aa925e527615c6c8823337492663a3c3977d9022b02efef16ba056307029dc18645279a8049c8288de374a8c75b4168c1f61298b9ab52fc7ec58bdd7d4dbbb5318cfb344d6b55905176ad99d87445adde5838c61459f7be958986363b2176436bdcb579a2fc95a77f7cc87f9c46f5e0bb9982a6d5fb0117a32e4caeb8a882cad860bf514797624829f92218eb2bbb95fbc31cbc5c47ad792ce170a293db0ea2937be23a91f91dec31f5331ef95ea9eaa82c7f37b6974ac7bbd8370bd48620ad3731da63c0c3ac3c55310e288c3b71908079ad401c10f6deb34af98baae3803e617a80d0c0cb75720a42cdce3eedb8aa52ba803af303960e7a4f84b6a384b3ba6aabed20780809996423d0f2f2249de3b6c36e5388a8ab26a2140cb9ca94a38d526f8e0c331dfdae95522e881256366b38519dfc7b2042c056f3f337965ac64701bdc34d12aa8781f5e7c8ba7a57cd5a5be58ea056b999753f13633f1741183142cb519abc2de5c23bf6d285b9726ac326b6d5b293764c34667324b7067dbf3813f4ec27474698e3dfe759c215ae49aaef06a341f8cd284dc8c25103244fc037431754f90dd1f0fcbd517136f8b5f7ee2a34c03695b5dd45616d6e13fc9d828519ea39e5182437045daefc9e27b800760f7c53d98ba88df6e1e61dfe82ec0bd2f1814ec0c869b9f3876f015b2bff7375a7e2f6bb24ea0c52d6f4527da515b5849a7357c8745135f28a71b1b341c9a58e6b7ef6e313d9023614d91948714c0699405fa996fbf2deed355b4ab5374b834dd86cf94bc153af5231f1cc5df1daff443cc12844d70336a39ec7689414b1f157f218e45878e89d3afac53f9646d8d43f6396ada2d62373a0780b5fc747af614a7ba2e024f8cfd1b26d02764ed8a7f9793ab545c0116bf0776cedd0b711ff2b1fc1e5f8855568df67130ca1289792f353abada7f1ebd48b27433e0a57a536e339cee949e835113a20a80fcb209c31be435e66a61cb94a8cc11fee5c4b311e64a0f5062f8a0427e763bee7f3be04e068023f114ee0cc287b6c4b11f8f4d987c54bd04f1edada8b20ba80c1447a7b6a605216813d4ab5bd68b75eaf9e99dd2b703c5aa0f7ead72b758599dca2b64a0f2dd4e4a00373998fb76881c0246ac8155f10dd57b07d8aded0dc49bc955afd1f8eb9562cad423bbe60ac1450a4239611d9c70b4bde13126632d27dc4021ba012d731eac34b8a080c75d5a579c748ce8ccbe963b6f0bf6c1894671fbbf227be11940a7c0a4d3f5981f2a6629a1122588f779fbfb6354607b645757517b31e3f7a4b31022514edec6c9149f98b69b4b90f3d8017ffaf2b1a5ca2044edf008744cfae8057a091da69241bc0c6b295935d8fb5443c8b5c67979ca188ed0546442a6ca554b53c23608a0f882cc1d380d64dcdbf99bba0d68645cb9fd076daddcef56addf95e528f798fd053ec9314ea343f3649aa0347109245f5d0bf96135bf9b1de0f50f7637133bed004fbb21de88a63e7864f91aa4213d9fcee40e41968b94e6f648a1685e6dacfd8045d619b15a498641aba553c15e1dc68cd93ca0e855d7d007394780e2770f50d1762983ece8f958c36f5855e3a5b18f5130d0b8416c2448479c71ed82578bd461d054472b302a276831d0e00c82d5366de5d6fd54921c0f1058df94ff88df4ab941ed7d34d6b72806df532cf1955bc965cf08212dd00036f156fb9ea11b7befa3731d99acc9c3eb0c5cc20f434caf2656875f741857c9763468aa5a80976712036005a9725d49ca4cacc4acd91948cfab9c41c4fbbab884e32abcb5276948423c07afa1b0f7d74cf6fec17fde668c7728c66641fae42585803606e7981f4ba1119457a01d112fbfdd41592657200547437194f38772bd00581827c1e01db1b9a6fd37be0158f7172b86bfc7df86689c545d7383931cb208791a87c8cd2859c400b843f4bcd9c6b17195e4224a1cff9ffa4635ba2e292f4684524697c3d952b3509aedddf870d1590d5e44b59fdfa5dbfb7090a268a7f9420dc32f900bdbd8d008bb3b61cea977eb0d7a4b748eb3b27298606dc6c8d2eb7feefd60b9a7e3d7bd78da8f9d387c511f55de24438aee2c7c794c3c6e6c232932ca58327f793948610f90275c11ac7c143d0af8ca6a02f7c5e1b9a8b4ebe2aa905fe789de909ec5b785b132885e371d16c7172316378ac9d1f04469052537db1cc8572154e73a71ece982d74213c13471cc5dee89b405e47ed0df08916fb986f4053562c247281d6787c79989e943f36840dc202db3045439df665d742d6b4ff6447b2b71800b64540bc0ea0885e97992e658147bac97677d30eec8d1a6ad69ee39b575a8d813e28e097befa08b0b084c88e7376b42cae07a274ab29712ab076ff6645607f12dee7e31b8188da8ff330f1b98f85681237174c40406cd69662605e859e55a75954bc960770659d9aaa5a1a9a62ef193068cd37d3947bc690141219bb6c1e284509d95e23b68b23c166234950e3dad25b4b0da657aeb41a0d5b4c8b75b8f4c4f51d7c4abff85781ecbc0a54116d2775abcc7e2c8fb4a1e14ee212087d6eed5be66e911603e3efc52e2fcd45e89c330762f3620b6f20a95b95afeb35954e093adfd0148302553485ba3f7cf64b90aabed6c7b7ed62bb568cc8a03cb9d0bbaa75147a7fe5b664fc5724cfdf6fb2df261be287df0cd22dd42d5e706adbd0967e27dbc9108f23c1b4cebbfa8bc1ade86069758031ce9cc02ebe74b1bf2f76dcea17275f49fa7234900eca37ab1f9cfe004ba8f0d118860e2993f7a00e42693154839c87cbffa3e4021190333ae98d14b366fc08a82e0b488cdd036688adf1fcb8345430c260d2e16dd6aab275ea92c07b815250d82d58693cd3bd8769590ad7d045599e934d5b715f7d3f629c3e797ec43d451d43d7b3ff04ba5b3d5ddacbcec8f4c259ccf4475d4c87e29fd0168ca6e7e70a723d5c69f3d9d034e22c7a70772fca45352770d5a70144e45787a86ae7081e77874dd7eefe8f96f76b62f74225acf0a6c94ad4b830a3e79c39f96362f9a2d219edbe680bf02dc575da12a60ac1dd358b865e1985005e83b0311e7add9f1e360f7392ca6528bf4cdba0548d65f9c2edb0452a2a24f747e7c8f9f1652f2f822bdddff8e58435a5ef8c8d07acfb3d84ba65eada18a54e21b2220d5034d7446dbc3905fa862a9960e27240980117a574daa29ebd5ce4a60a90834746515163e8aa0e13e02abda24e6f493dd4c951560bbc1d0201d930423d74047a69ab49c6ab33a33d4c02c21c9349ac20c3203a7f8d1c9316c80e2e6b641c8c1131c1c801db6b5926299e18be998bcb68d4e463514ec083abe678b5579522dabe973897b88528f90e8af559bb041b1466661b07e66cbe01adbf8f4d0bf9190c543ec5c8e1d8c7410e4ebc708854ac448fd21bc9fa7999d8d617c90257ca2a584d85d1648355f3b8f6d042b2ae27f1c908d947452a2fe570f24e277e410ade8f3a4ffd45551b256d2b21440b2686b782ea545ee7f1b2e5d19fc0ac316352b80943ff4252812f14cc6a15d72b5b6600a92ead4c70d33961f7b54a3eb1087228373e03ec8aef040912dab295d8c7f9a1844209d23835c60aab2c14268fd7ecb9ebf51e39f539626e8ebd7e5f0d680db65c9793a22c01194390a58a89f4af317b5c444b75863af7b61ced15fd942c3b273f5a27487f06d001f7d5bba793905f8099adebb0fda2de4f5d34926b84081f4f8661655583e95306aa1eeddba7d7046bf93fe80e6d486887edbb762fcb9e843fc73231731cd431902539e18190b32f301ff421c1cf4d7a144266f1e220302fc30f6cb4ee87aa67c9d162eb9d30b2dde3011d108fccee7912426cc602b0e3a6c846389560855d56fff1e2cd259b2cde74a2e12419013aa2735380fefda72fb703153f6ec16e85b1080ec53dd75cd7e56e9dafaae00c19e0baca9c44e6d730ee1832e06ba7625521f4bd5550346d735547dc8f4eeb9eac64e2479ec87c64e837d802ff8403758aface31fff20d49070e036c5f7dcf9b240e27ed4b084b35107d5fe96e7a429d12e14b4ea07092d81f98cb7f8a69eb599f914f2a52472212a5907c7d7245a01ccd46e6b423021558d1b239ba627f17133d836f4f83e0c84bc084a8698014d7cee47ae53af814f1ac1ab9010bda80778c03e041e1758c41020e3014db5ac471a87a4c7f6740876f48fb67dc3c165296cbfe75e24e0c7b29e69d05616b2e582f8d324ba23fd55211f1aedee27b9cff2d77ef8cbb9ce50f59b95c1385915d7ccc4f891b2099983ea7ead6601ff3f2b83e17cc3c99c1a40f0701a0f418df38c470117a3ebad501d8c219bf4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7a61903c110080b8f2da39322b740db64de52e7710b49a5fbe5f1e7dd9867d091ba5a51dce530ba4719b3e02fcf68142bcc9467759667b8f6539a26de925834d332ebe89638b8cf07e7b5704ad37b696ab15d315547eab7a5656986183e0bf964f3cdcc671098196a9540b7b2fb8bfeddcf564fddebb45b28351d9e2f33b817e1f1b87d1cc61e074c459771d3b21a7bb9d39b4657084d0328db78b1681797097a637116f71ac0c513bfec11a0bfbaad3d015a796ab70c7cd2a81a1bd7b06c1b648d71f7b5584452b8c313ee19afede0ec9d7078c0993938c5323ba8200bed9f615ab601b1c455f2630cb0ff3a92afd6dd0e4fa7061d07b305a4abf306e4fb467a7489ef3ed1007dca09bab725b33152520b89ae61c70bfa99a2ea0095432a0733678c93ce3836946bf46cf8858457c1093a7983ab3a96b50c64a21e271e8fca67065ce5ea5560a073958fca72b8d2aa72caa828d36aee4702974274b1be94b69be4e38e86dddb3b8a7b7e0a0247488f97e96b03bd0733a8821d4eca6c05f26e8fc71277127d25a6485f5dc6970ae12cefff6dcabc550befdd2e52ff17f1d9fae4c8694283825bc07ec054a5bcdbc0e2acb5a1f2807e98bb9a7a9cbb1d108575758e0dd78d1b9264d8d90943dfa806b353ce0d5ec5800af907af20972410cf8303648e58456c266fa356a69101ca1478a2fc8595518bd0d2b2f7a34a8705957e32f13e150f5829f752cd40684c5c47b1e3d300dcad8fa08c3799e8a387bb2f27c4f5f3e07b92c5fd8b837a225b11ef1c36703aa3efb334d3c7945eb980fc1c7ca2b8ec576a3440f35866d35b56ceeaaaec054bc87ad7c81832917d1705a2c30d5d59fdd87569a3ba6a51f1cdf893b976878e7a6f419c6dd5cf35c4f07d2d1d26ae5cfbd957dd2832b07bd2a6d0f807ae37b242571037f8fe4a607f97f75905f722d353f34b881ac3d0732d90dda3e416a93256a1196e80cb9bacc98c16c0f9c43fb7874937d1bf31f80174c1aec53a2d50f6caa37a2b15db249dfa55a629fd282a09bacc54a36c9c86f02b60fd637899482a6dc89191d99644f07d0d05b35ecf24ea607b398533be5af0b9894aab24a6c1c6603fb8cedc6c35afdcd19e3ea5b5916e3455061521fb8ef26ef22cd57c9df5f00c0d2a2d697d5d3402528d6ceb15cf8f1742e8743f496c088d66d24078bc8b9fe1730987b2b0ea719c1a7d10eb5bcb1b0577a332e2d4e73667550f82360b1dc65aa1d02dd35bf0a6116c7ced1e5fe804a72cdefc7b2d0d79a4921cabe3888650ec615bdf82410bf569123fa9a8c51051c644746bbeba7b8a78a0b29a91ad419a970dc9a753e20588093c8619a947deff8e970bcf64894c00e832b5445a2c238589049544d105eda3d894e07261690234ab2fa9cbb678609a8dbfeed953eaa856a5b43a882410deda9cdce627f86cd3e89ade55e7801371cf85b84705fa18a3a82f9d4093ce0c38a047c43042cc43d0c9b0940ed2f74172dc28b13f15859b63c0f18e9411ae1e6c03ef76694dc0080555b6a4789902d50966bf34da19703cb1df3b1b81d9848bfbb349007155f5805577f493ecc241dade25dca14bd4964a90bf08aaa4643861245328ead057d2300b7f6a60ae8ff16e41c2cf1ea2df320f769a50b7fdfa6af8146b68422532d290df54bfaaf64b2d5bcdd728aa4cb1a5bdf64c1a65af2b2ab354cbbd580210ad0227de6c87b2b97a001cfebcfd733541b4e1d72ff4208981d5b24ba1b3df512d0c02a9476c541df8d1afa63833b96648a128bbfeacc353da59cceaecd5be7a21715647522c6ed93ff943a92aaf825e06e492eee46cb5682c09342212ebd326fdfdf4adcc2c5241aba0fbdec5296b637903a516c97df3211720b9a7bc4ef7931fad474a8a15a3b57d0fd7424cc0ed518480bec91bdaa71457de6b0ad119080e8286aee3435b1269b74a1cda48e54e0a8c8e65f168bfc749ce627f612321670d64e5386ab58886d99d816c9f1952924a9c86007ec9179e8919268d5c7082ce50ec66d775184ea1820cf9f8c924ea4b3a80870f4ea5ce916b72af13c51a67bb983c26d136aa9364c5f7fb8ce0ccaf79e1d97b689fb7835c677feff5dd3511d5638852af679c88ced35a37b09af97792f1c55e92f807e553507a4e2d036bc9290ff14f8559276957706ab78af7d702f8c9643c9c26946d4b22c1e80a455649abb627aed5edc58d8d4b5c486a906b3c14411d591249794ea675491e30e6b3cfee35e9f909a50f421f1fd635e3c4f7a2f4bce8c3846b6a2ea9e4e81113e1a505e233d8573430d0de77124c69535ac31b0114cf30e57e12057fcd1080260696c06b757a6d71adfebab9b354efdf3081ee30633f018661dad24ebc16975eb18fa81cd0e7c4fb2df22e691ad71721e5b7b0aea1dd451baec46c64df2baaec83517ca69883a742d6b2befd54f8708f56bfe5babbb462afcece94cf6c9e5e77b39a591687e319c9a37d3000fef0152618ffd419f590797bff0415603140340389fd4c43bd1ac1f6db2919c3b43245b92f0af8fe19723b09e755ec238c1e7ef9750be538f945498e4720b3b786b42f4b2e45dc859d6c01b55a5e98bba688983018b583c427249df02f9c254092ed7193945474866cd25252606a5bbb3cad360939954b75f254099cb2f14a984dad4924145d4b578f3da9de3a117a1d1d903b2b3d05e554c211049ef4b9207f7332daa3cf7baf1f0f3a15eb9ff80f5d8873e345304d6d7e6a3fa549b1e973fe5b7d5cf4ca8b3539767dd719988e343dc94a293f58ca2cc31be9233c02a5e24ae3d5cc2c2a07b07a4605759f5d69a9f0978f314e8b21b76b0268677c322770f1857c638d0e89e008552c73818f8f3d7d515ab090923f89842280d631a880bc6e6cc545fa627ab4d264f2558cd8856c8d480a6edb12619cb4ad656a53952809770830a1ad74440452dc9cbd51da5b94863b877b3b40c5f7d67190c5c9474a664aaed1b5da24be25107c7f3b987b806f336ff235046a744fcc7c0a5d83e10992ef311755ad3b72df7f3ef75303f7421e8f50942dc72a59a2c0afbbd01ed45a992c02d17719a6067625ef4db5826832d8d77c40b7f99e2e4311d3a3ebd0631c5bcc0abec6ef8a1a6598d52915007e4f02e2d23ef9b1dbacb4baf98fa737958cce22b76c667ac4f497e1d73287b7c0c72d4e5f25244a027ff2fb67efc98a4ffd5a2b2915d3f87c25dfe0fd8c68fdaa21acf82f9c8229d82701602762d92d32d934019f19277a21241996de1974949ea48c2397a1da9782716c404f10529598eff3bd98497e199b68a6373952f9416c6ac5df24c90405e78aab526473335ff51699686b074a2358fe41d63bbb81462d6925188ad5e33b8c528a0a246ad868226b856c676a61a88107dbfcc26d8ef3aa5b20ba09f7a65fa1de204461b4424559a9910ce4745b42123b68c5cda5d98ecaefd7a9edac0e71bdc08d2dc032a4411b4e79088d34f6f48e22b39b0c6e7b181b5eefb18ea65f4272ea9366dce72e7b3e5523773e9883d3e4e06ba6fd01e9436738978584be2d4ccdec4b0f38073e6c0454c0e6d2037fa590e72ec987ad53075e258dbe9950971fdfd603467f560ccf89d80ae75bad541c7dd0c517f8fcbf188e0e3a2bc748eb67dca68860b4155dd6bc8ff7b4a9966b32ea0ad673253053113ab7f5c9e0e80aedde9ff6e0d1591c3ec1908a4147d4f1157ffcb1c6f154dec95ab5801a2c7457ea9de4230b67ff609f002e321273cb4c43e19f21d385021cecf071740053c838f913df41c3803c0d35c9550b832a5fbd222f91c5b3e4996d7550106d378b696e2eba8365eb409990572fb5dfdb497c6a337625e54ad45e17d87bfc38980e3d3ca93a16450498ae22569a7a866cd663d218d0d6d0e4d11475847e9c479543a93ab17a574f4ff883c06484a6499ef9c1467a80758de41fcea986964e03a8a3ca435c935193dc7dc01ddc0b2ad2605a95272407bc4a3fad655f3090871a683a9bb9dd38287120cd2e1c7260f43484edd291941d0fe5cd7fbd4389f51e5d8dc9bb7f2439e35b28efde695ea2ce7cac4bba173127eb5be21a7195e0465863da4e8dbab58600e03835cef2a02ece9af9c1b0a3e946cc86048d5e2f934d3b1416a0a91e5558c00d5e909df58489912fd87f166203e74f540a0b66e3610b6a066bd3eb35ca25ac80a52399ca85a1f3be0925033925262ba7998fc66bda11eee8abb46b74f3f75769dd20ab9bf713e6ae005d4509c30d7b34262154b547f16705091645748ce112125f90705c62ddc6bf7ddc6628aa464ab4e2896c6c367bbbd57ddd004ab91e014e496527a5def2388859e9eba2c154312299fce2d9fcc40468ce1315ed8b49c602d8fcae7fcc6a4b742d70cd5270bb2409ed7d84c706822d0a3627d7b4d602348d5d299f633b2300a3c7c5946968092c1bd8834f4969a57f63d25d49adf682f3f27a42520d1698d94d4755ecfb9892ab2c94efeb813ce03766df2d13d939aadba5396dc6da8e5109d7811d8eb5fefbc4dcedb314dfee256d260f61297e75cfa63501fc05a0d71c52ba5129c2bc7a68a5bbb5963b98efe6a6065c422a55948c2db9e7f115ed877ff1d5ba8c0db048800039ced9e46bbdad9c865112b2234a70fcfaef89758d815c8cbd13fa72f88564d62887f65f1d18e182e3f201a0f538940470d47a28e44b88e9941d8a8501e45a99355711cf1df94d2ae1d393670cec84dc13b89f7244158262357c66f8e110ed4329374d2096b8de7a4893e30a2a5676d39bbe3f4a0e978ace74545af235bed9db82712cbffe44db8a8fc2b47d660ff08595c220c67cd8b512711e1f7e6189ce3356ab8a56351407c14a25c520c601fe98ffeb313e8f438238a2ea425696ec8585c80a6c253bd55cd9bbff44e48589d5bb9ad002d970ad237e95cbf20c0fa0847e55f2daaa1da642807687e031085f27ef1a36850c5df95bdf6a814248757581ce290412af15a1454d3fd6c471f50d445579cc0871fbd8883cf5bd6284fa1da17099adf86f59ed53b8052ef8018bb863786ae6976487c19b38dd0978e73d9714af9baa107c8a712dd6d98da30a8c316f0e07fb7e751e35192086c497a8041136bcd0d002b10746dd5cc3891e62a70e7ec005fa2bc3d4583d920863f30ed94ca95e425d6f09d31f0323adb490c47bbacc0e99498e9119ded8eef80cd15b78e2feedeb4ebc19f91913f8e9c7872db1e160003c656cf76b55970173c85dc25e0290f26cc92e5ad47c86411a4baca902993315771201c48d0c48c6c80fe5902ec655b22d874a06a1024906d854b592b439e627a17e59e8e89be2ad4236f68cfec7a6d2c6bf0f9b52b7ba4bfef455247a5dd0c1029a8d9ff4802a25f14b1c1248d298f1854892817e95239f77962f00e2a2c9e14de01d296489cae5847f8e492542091b773a0a1ed299e985460046cb9da9dd9f6d98159775dc162f2982b7e809d1388928521a35885510fc5466aec579a543698fb2fc4114537abf6fb31d6a422989fb6a81a4a5f2ecd99c2dc27f80a576387fdb2ea27a517f09564c018c83487c72133aa77c8589deaf2d201802739cbd729af3f67f411509df920e8064b63cb9f72898f6c63fda0b99ddb8f6105519d513c72e32dbac68667e3a3c37092a116ab7865169384f74ece9e298c60895fd708c8fe27752e94f5c73c381ff24c07c2806cb4089bfafa6b3ed43d4a3d7c9e76ebd3b38fff483e1f760fb96bf0a782344bf1d13f42592320dafc40dd560002d5bd5b198af195c2cf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h35ce176a93a1402236149c97a4f038f38bec07d950219f6b95597d8e7230943ff5d330f343ab72484b4df4ba3f8d689d540ab9b8157afbe3041fd1176e02ebad1109ece408e463f40f13b098cdea0019f76e7fd155872e78126500a528160e27c6be7fb2def4406676e7802a3b5448321880a434e60af49abb8d9c92e7f9bb3f2db3c3b8eec774ba53f8c602316e662009e444b3cfc484b02765bafdecfcb6dd4cad283590e6d9b2fce37156e0995f4bdad10f83f7f2811350c5189aa69bddc9c28790133b95b07c1626b115dd691498d16caa9b7e14323d609dca08c544871ac0be929726bd614d2bb12df9dae7b940677379889fbaa42e0b2f8365e48383fa860c156a6e95666dfda94b21624629202d4df93c5526b1803eed44ddb467cb3926da271f42e15369569db835869177a98a4a4c42bdec0e99829d5b7caa706b72b835718f5799fb2b5ec035a61545006f4968b1af7b2a7143b50cb1180f1b99a3a04eb327d84af263280b33eaba18e465f865b5c0b4d84771663c6bd37119416ce4b3aeec388e926e1a334cb4381aff16693e4133a90cc5e8061f673d3ed17786cfab4f14935934c50d56b9fd5206e4e925c5f44baf8e8e77627b02673f6009cfff89b7d47df47baaae91e19cdfce306a7cbe5f088d2abe8f209f5b8733d99e6ab9e845ea7a9a385c4d952f67a55a9041d797dc58a947f0388af2f8a6ef08d689e3680fd0b9cf4dabd64f542e8af2d67b8eaa1e692bc1aa291d8157714d8bed61201bbb7f0b53fda53aa8538b0a515f99fde63f7fd70b83bf45975971cd2ffe29998f06c1a512b706b700939a0ca3a92cef5e41923f52642e1d63d8cadac055b3a966715c9aa15103fa8405e094fc9b70c5ea0e10e01d51a8e5a2ed16b1f968bbd5692cba6513283fe4e5eb03733b9f221196eee78051d88d57d1ade521b0c094e9f5dd72c99e99945c7dc69a989f85793026eabf2c9d8d069b62929caeb815adb103ec2897cff9a1cf7360953f2efd49a32d4205722001da73d734896b471cfb21da334fc0df09939fc7855784ca8b3a53305b046acf8bc7f4cfee4409e97dc9579706d18661468d09d908b82014d4a3fc292e23ac548f525d9b50b933a2e082666a24a1575ae1cd68fceaeb3e8b4a75452c7875e06dfb5940562622b664a873145921b3c5501a3f61c762e81fb981e739d8f07b1ef48dd498e96f58adf6c086ff97dc01abc136a63b7297baf579b8a73257974ca43cd828d690e71d768c5ddb754b6be499f23a20860a7ef796be690d7b077684daea09beff3f53ed549ad16e9a53b6e94142f445982e8f9805aff7ecd67b551a3e5ca548b8a52d7003d3e582684e84a5c780c0c2e452664258490b16b2d61c586b5c04b4acc918dc54a46f6d804ab56741216f9738a48281a010d5db514c70981e8b81de2e8d7f426d88cd7c4c081458f3cc8d1f1d9905fe647fe0fa22e0652ac6f12d70e4fc6d2d551179e5fc53412c40d1340eb958ff2491dfdcaf506c7bc7b4948ed84909a6625c363963600e34c9b48fa3298c3dc00602430189d4d8edbaddaa6ef4ed202192bc983690c8edae2c4ae1da777489deba5f7bd314967695bd650b1869083d22b9966a2e55e96e70ff55b1c4b87dc177fa81c4da5239098d22cf09294fc2f8f5451133312dc1cf5e745552f9256c5bf1dd9c4a1cc947b45d428b7b015c15eb7d371ff89b24f67810f31ef53fbfb739dd0b64ced476e4a4ee1c4dfd0b4a8109d43ebd8c8bc7a71e8accd87ea410570f8d27a8fd46251e4a383a730c56a1f87961197d4e969b47781570f4fcdead63a5ac430d37a937d3baea3cf40ec3749969fd1e61da1e6cfa7230043ff0045c9a97a5040b0898af4c298129aeecbda9a45f173b0793b266cc72a1ef56e546463fb96f2052ff580af57deacac55543f9d706c92493df120c67315feb258936e3c2f304beb7fe34da28c32bc76cdbfcc6925f552ac772bd7adc503b41e359f6ee317c4ac0236b23f53829e0e233ed61cb2154d12b6d7609d0741f93947ffec6545dbb6201178d703b775c0302c42b4030a08babba98ccc9cd6ce24b2d5cf26e50a46db7dcc37d442225f52dbd9b272ab202dfd4416394d28c400f21cd28c27244d24fcc86c7b0c3652556cf2f9c00a6ad025aa7868c33541fc1756316c68e46a4015839bde0acd56ee0d3f581565ca61b3964a7bb1c0b2d3bd5725ef017a51e5b4e4a196029c86a30c63fcd5a836f6090905befc72189c11d290d8505fa0c7a260be1dd4f8c7bb9127d57977790b9e2389cbcd8a95f2cb758912ee36ff642d310fd389c4835301d286780a189454d32ad4ed08b52f366869dd199267cdab9aa10a58707d560091040d068ca678ae8a958d2b193cc754b159466b47198c774b2396d3d162f06843c32711da3fe08090c0680bb2407a332999928c71a370af299b1446920916f90463d0199e5565644b79efd21603893ffe565e8f0ff9c6c7beea1d50a7ed365b93d2a9c29ffe19020087a1748968facd2f080e6c24d6380da34549c2605daf95630631ff842bbb8917b43911fab65905fc8d1a969ff9c697f10cea0ec307823fb946bed8368dcac0103888d851bdd99cce5e5d764131ef6d87272d51c2d1a0e88bc874a7fa36389cc12988419080eda67cb6f6ea490d8817f4c37e696cd06ee7967b6b3b41d87d5a7eddf161c386f54128d64c838a2b7c71cd9bf90e922f4ed643abd4f493bac060fc36be8cde76ca96716984d8a124f22f75692a972f167468c3c198a2861d28e4c79b75b754de4674644a1ea59b69ff6474793e0ad95a43e3549b52a666c45da3b33d0d67759af3e71abd31046d17f11732189ed2c27a8beea6d39399d31a52fa1bea15c7cf42d9da64cf7ced6fda8190eceedf00bad2855435ce147efb3299e20cfd676635551eb99a534ea5eff66a5a19a0054e9cb046896d8d8b9cea800bfce38427a1ce44a4506df9375efbece8a6d99087ab6b2ccc0652fc33abb084d0bd4db0b985a53de030f801eecf0aef473fbc0b60bc8270585c41ef9de8c9d2c020ef7c263b59eebfe0accb19c6be1d2ef964d8ecc89fcd0cdb95cddba2d323674e72320e3a4b257a7baec3b6be1e9aa0a1359df9dfb2f17cdee211c3601c1bdb5f874c7baa871f2412bc7c8787c093b91ac3d0722a8736722d1a92be052881288babc270ea77322ed2532cfc36b39940ce83f41dc9aea723e28d7b672cd899c55f6abbaaf9d4d412d2cb541c63d7a88537395cd30b3215c9f76553622bc1324f239b5ab4eb7637f2c64ed91eb787da71111b125be42f9327e0b6327ab6ac2c7b540e439d3cad3dafc68ea21f3c434d804200895832a4c95da34737826ecaaf02789fd65ee28c2e036df33a08294c7ebf16e03488d8ce5c089e99df562e98aadf0f8ad257066c32fa36118d6f6c33705687543ea5a711bff82442422e514e10787547cff8155fec718be9de25bdb707f422ffb449df77b0baa786292af1513c6f9cb053d217921f8eb0fafba1db7af568d8fd66fc3742b147f8af53e2ea72d8a9bf85f77bf2f34aa91f3d27c07b09c8f2684e0cdfb369684dc7cac84275af8e94916283292b27b7f41601305bc73dc6854be7750678090fca5ddd1ed9cb01beb956632903ddaaf4fe4e827958e48ec9b6c4075f8d1c661426b547ac5b44af18b1c4a503c7e8c871ee4845262778540d2580303434d0b879c7f85e336663a024f9e15e086428c398384545fb3291af6f8815cda464e120c2eebf0356921ad791d3607d1ee03290616d32edf9ad0d368103821e5332cd3210095c31b9ea022d26cba27026b485221a4e893f7f2875e10541d2d4a1516bb1b207cf5d00f4a85e87e3861a7d4b1fe21fe856a8deeec90ee7388ff06947a49c729658c6e44076ea5660605e68d98e5e6d67778b60ca78d0f1ff8fb432df2bda83cb455f0396993f259b35c7367eff231aa02059438e9dd7998c611e5c08fdec17d8bf2c57dcee26abd43a6d4588d9a9758d876c177a082879b9dbd3945fc144def2359d4eb1bdf021981024bd1398124448dab601b87d345ee4c7dfb9a99e6e2dc68d4b9d1e0a533609b9decc36c380d12a7c8fcc9d58cc9186a94f3c77288790ce47e254baaed1d54d7069eefd209181e805b182f9862b1a8743dc50ba9b2ac81544b28b7b29ffb658843924ea2ec44a59385399174b55b3cbf78a8351594c5138ec2b999e042ec696334d893a62e26363a1927f892debfef6ecfcaaa6de9f01d9dc200d6618175da422c82d56509ef88ad8906202abc61fd324284b708776f3efac6687c23b7e4292ae0185005678e076febe350e2444d9dc75d84a07d2c63928df36b265ea82ae5ffe41036336c93dfcb25a9dc6361636595928192a40b03bc3ed2a743507d89c9d87708e03b58e5acbe2f6ed42e0e7a1ba1a8aa3feac5979d54d4ec4ef81f914b224ea7c785c75441fe08482d4051ef668ee200329205f58249e074d2eb08801ebe495f682a6b40d27f9b0b29102de5c1d59b4fc4536e86c0154189e2ba39aa65e3c6cd0822eadbd4a697e715393c4dc9336d6f47f5d238b9fe582dbbd7c85b2ac9242dc014e99601c3197627dc7b6dc48b3039ae61c2e7e8a91e00a6cce793c0e3c0b1a3c5080a61317a6503de6440df992f0be4ddf8bdb9ee56eb587f648075041c1a547a09ef6fe5870ab563d3dc4926c1e8966c5219fd97bb3bf2a5f68fdbbb913e62769d7d6a43ba37b23b4e0e9a89e9504061849522a51830ad0815f9e0eb289e414fc487860df37a6e4215babd0f04f6d241b4ae4bc07379142fb8e74bb42d90633596c45889cbaa8e22107ee7af6540d1c045e55f4f5134ce42472196a47ca032fbf364be8442723a2a03aa1850d9fb5d2fa223e18154d353f2bf468fc590ff514fb85f1d41605ae0e9cc9f06d14b0c787774adb50d121a0192d0f80a0da1aa47750c6ce53933fb311afe5cba337085141cbd47615632d6183a6eac7dff06ea93944f9226e33d9fcbd5d593a3112cc2e7a980b48c1bf04ba62a095c4887c42498b1e03a86dde063a998211e8541448cfa4904601bbfa9a759af0d7b0ae9ee447ad254171ba48fc40156fc3bba7edde213d4d2b3f29c46207418d8a049d865363c5c288ad5fd60d055b4f98326ca4aa33194dd99d76c84da5e20c806d73b0f0ac91bc03162fc13d6e6e5035469ce0e396811a11e50247884ddb542dd3990857b93d333a5a5e7d5ac9c3b71db066b8dc1a58796a9c875812b8c508a8ef663b4c1a5e8f351b8390c8e6dd11b347696dce3d0b0e7513ca57711422e66bacb3db43da3d7d5f8a61a85c89e34ffe24cf22111f601d0f8d6c27cbfb189b0d8285bf806d04b5287168498a8cf871dc7c15aab43bb5e6fe5e1a191fa0fe44b436d56952a1e1e3a170ae4514eed88b32ceda6fe250d9ba297a00185956f0f96142c3566ad442515cf3c87473ccf9250a8f3a2f0c4167c3cd9277c0ae9cca15ff8949b895e8b297da8c5fce83259d051d654765e03c65e29215bb0c3edc244614d8a00bc793c8109801a9c407373caf690e088cceb04356090a57cf5d9cdeaab29b62958964f681ccc73084d41cfb216f0dfedf71ec9c528727c47e2856a7136cb1ca48fd6ffc4cdd98e3cb0a29dc43a8ddd7160064f4e7d89c0ab72c701f6b6cabd05f614a2d4e071df24b8e7f51e4f282de9debbeb5f3a2066aef1b75d1d0865580e8296dcbe8c7a00ecf7dc731d8a3005dbda14a6978c162479cc652394d105dd036ead7440223c470ab028b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hffb3d50dc95163164c987078c713ca61866c44e42e03cb722ba465344008d09e6970dea1b35181dce5f0a6d8cc9359b02ada202bd12060ae06046aa16d174a22f8f8ba65a63b3001a6a35241ba6c8713294cfa2dc2f7f13f0c6e43f1fc4c9cafeb7bc404b17082a42b522bc2676b2e05686ab9f83e70d638a3490e5388aa6e0f94ee766cef46af7f1b44cf0550b10e6536bab431984063fcfebacd9f03378051a6fb71eb57fd308810b0b98e6b96b372052d239a033eed979c687abb71f3728d1302e646ad9f028104ced68e30f30f497cf5ca8e4f43323ac2603f8d317d5805e3d784dffd11afcc0b60db51dfd555eff53277a9c1a38ee74a1de36a6435b7ef6523c63402d58147f680afabf5311dcbe02e1c6473961e10db923c521c555e74b787d86b3d40fb7f0023b3d27c962a05d3fab2ec656377c237441db9e15a11ec4066082f95b42779f788d5167f326e2ddce4fbf15838c54a5788f13e9581699315a73cc09183e7fb60f722fa4315bb85ec89185a3acfe77fefc0beb12341a1838a7e20af1b914140c029f970fba482182e8628ccf9c1cacdbe261df5afd6b6478a08b83fc9897ce3c1e998da9fcb1ea7816cab1add4d02b55f9d39e1db9a33fd4c7a04063f3b917dd3388500248c3aec6dd227310bf44f425871bdd0cec46227df20681296649b8efab7e2fcbe66df869ebdb3d4b5b77f755f80ee563fb7198f2505404e0f55be988a19bbcfc16476af554b488de12036656e311d7f8ed9972e2e766fd7dc74799d84f6358851a584b3996d331a77380bfe0226de8e7bf3321e3773a65112051d8a9531598ef831088db9b609b02edd11984827f62cc9fb28292f73ea94877984e80968edcbeb077e786cd4087f9f16ef82e02798b43afbf84f1e64b9d7b0190c213cf3a614c647df853e1c949f34bf622631468d31dd33cb85b5dd8954e4380d1e0da62811495322049de236fc2d44cc69ccc5ce30f5032628ae4eca9a22525611966723552492b156b9fe00f5419ecaa29cb69d0521f606eb19d32550b2f6e9b71a5bf6ad1682a237572cd5ca791aa5c14de8fa844b9dbebc45aab61e3d713c1387d1daa2d23c1138979aa55d3e7dc6afd5ac27b697f427133b7ba142632c730051a035a2fcbdc2de2ece94b47aaf2bf31b76420051cee05df0386a257e1cf9152c738d76b43b8a78de0c4f16e9cfd30d8d06b604101250c3f8a894d9be051e2ee397ebdb4757df9f1fc7960dbcae4602dc81d3eb4bef0d9486d5b1c56994ee1fe494c288d92bbff44e6030191ee23a2a40cfee7b340f991a11fc00f943b39794128b4728f2337d3fcdbe55d2ad43f664835126bd0bc88fe484ec0234db14a94078217c0a28c1d8ade14c73c74b0529b4e4abbad2f213a4b7dce70c610d0e774dff8ffcd77eafa9eb531edbd890cbfe7d0234497430c0d2af1befea8d205379596314880e51205643a7c6cd9017bed62b6b9dcd45d99351dbf330bf210a7f35a089049f2c419f7e570586775e972d030f94e7fa691d2425da178c5f3a76747830852ff0b889752ebefb775e058f06e2ddf9d0d7790cfaec5d152a5ee7090b79a446471bf1615e9acd71e9dd3e9e81600cb0367f74c76bf7b6f96899401d342f5c7aabccacee9fe62a033fd7b369652ff8994dc429aebc1cdd7e8d513042a1cf7601df51adad289d6e8d5889decbd5907bd36560823a4f8577cb9aef462e440df2ad577580757c999ba5073a7376b057c8052f999c34485f64fd75d4b4b93733ca8417bfaa000d6b7243f7795b500306702cfcaf0c11f53f675c1783e2004976d7088f6ca5fe3851eedbbc9424ad0bb814e8510db56f5ce87560b1f78e73def498af1e3acfd8bfe0f615d1ed3efc8a5d4666d59221dceaedfd81fb4e0c36d997e6164f174cf1372ecb4a7b4ae98877e95ac2fba2c13bc901ceca1e07de4d301e0698e2d6a5794ea5a19a4eb36504e556d03f30cde5e19e44502c734ff7c3cbd572b16542398461b5a676a5b327bfec008f25e468e3653e88adf295f589b72a5a42e39d8e3def6dc9b304035dd384ae6af1192ee6eea05962fb68ec7b6c265f50a7650ff481f040717a97e1c51f7cdee3c741b530518386c9647da2124da94b52bf8540e0cdba9356fd92a76bb28f6d469c480ac73a0077cefe68460a07174119392ee5ed4c903e7891bea69a9e7ce4a9f4c350ffddce561bdfa9f1ebbed6747f67fc5861efac967a57b69b396cef03571b1e31466438058506683cbeb45d1ce3d677f993301105345f02a63c2a4005e08dad098d5524ee8517dc38c541536518d003e933780d516f27c4eba1617b6bc8b84f206e5018cf71b83e2eaa8b4dc23ee31d3a9c093a5e1ef68181903b689c8a698e9d3a4103335970b59ba936740567797d5075211ac412c0063596c290738b7e6cb06525f9f0b7f3c7ee68385b47408b51b5c1ead7cb05c4f7b73f659bab27da8172b6ed0d8e13a25ed579df9963e8160048630b3acb60b27cf65c3907c5700b2c9068919ab341457a60427767bb6486452a292010465deec2a6087ff26417f6508439a10682363e51f2aef5317f0050a3f973274d6a09b1ebef1f907778a50c9465e1c09f8b2d7691d5c0bcf39e9c4bc0c9f3b309fb1811f40ab80a6f91833d4169f30e684fc2e9646b508d0f38adee570f711cc299e34017f765949eeccbe4699beedb296adfa34c2a48c101d66e5bf0719a9d62e7798ed0e56d7379fcd8fdbe45b2dbd814bdb53df29677f522b83a12ce666eaae043389e9d1a2759805949b2e8d4ca8df16c11865348ffcaa43a596b1b4d0d803e7d026983442df27af1df5cdc1caf6372857fbd8507d068f4633be4170bd6d9e826fc3fcd2ae5bc0aed37d6ae8d892b2e52bef177726a6f23deb9cdd2919006ede4a84b61de4fb45fe1662925a7e61dee24ad9bc1d7e5ac34a501e387a291c13d05446b774e6957218cf5cbe639061a14d264945efd0587203204242ce23cfa2eeef4e954a2dd889ed630762f2eee9730fb1bd49c3d0673ed34abcd6f1ad2439b2d3d74532c595b14ed0b248534e9621bd6dca355c8fed0dfc4a11f05b3480d2bfad2cc0837b7e71bfc57e613318faeb58a36ffeea0252c5c7e61898054bb42f9b7eb04a136e14be83b9ce782940cb8eed5bf71dbd6b12187096f2a7ee5db8c5760b15888f76354e4f7356230eec264ecefb4070b3b0c6dccf9a4050c94a4e72081d25423032e7d9c96785037a3b7c78a42981f2249aef47a540ec34c2630157b7115217dfd85ecfe0e2c47be2c5c62e05f5d1b61e1fb23135873386db72b2f0cf6bdb0f3df13ece850fe545bfb6ce2465cd5973260cb561bde8ea27e4eaffcd56dfd6787287b91d1c7c4bf27fa779133017621c3eb69a05bef55b68da881702a190d815c7e2dc9414617bbcb729f28fa5a8b8a14d261a94fda32e41dbfbfbc5ffa2ad5f1a03f2c79cfa1de14e92664fb7bdf04e127005d5c8f219f583c9bf30a96f8efd1ab588cc73e6b21b81d218e8e3e9c1ed0a132f24b2a982bc70b387cf59ff1d2abccc3d338a716ad053f6d946a06957c1fb96d78816892b9cbed1a6b383dcb9f70a18faa6281c1feccb8797a347101f070032a374014e8bc4968e17da56561eba876ccd8b4bf646e5d3115e2e6330c43c9d32f2a8f2590506fa944cdfc300437afd75c7cdb1bbd067752c03f9075dda809e38f2fb42f4cd564a69c43478c10b665209b4536f2c3213561bc103c89449d1daa45b7ce1a2c66a3d4b412f7252ab3c142f2e644410850df68b257bc4b362879c1f085f34eac178cca8199c9e04048d746298c30b96b7b89fb85dad198c74bac7973fee0c16007d3e321eb8c49e26ea15a91fba81601ed18220f115f1327f28e1b3ed3a1d1bc7e35e3f6e75fe5fe9630df40097fc08f3cda25c15140390cdd41ca0d03ec72d2bd0816b4312ce526cf6a0cbdcb8a95754c5775d83533c6a85383773e68b6ac1ef619dd6b80a4c446797646862d3641e83721f170f3af224844e29fd060ad19d7b1a3a21cebfa68bbb81a7f50ae842fbad309ea68481ff9b464465b5d46588d4fa45c0c25108c8daeed7e96e0ec947f91649bbad38e8db8f9314b0ac43d6039426cdd3fb5ecb979314b8b565845af2b46ce19bf1d1c80969d02322e962d72f74e2138983d553de9ae76f60ef068e5d5354944b8d5e2b5d8fd36f43bfe984eea70b5391831fb2ba6d304b93c5a24d003d98a96d020525d9e74e2725c9b9403f07a41cf55b80b332337c8585e0768980351ffca797692d64963466ce63d7f6a4a044b1f6aab8287546be2b956f280c2fecc39a9ac2a0681afef7b02660bf59d0f82ed802f1a5aceb11010a420bc3ad1ff24459e0fe0ff019ce2cb414f0b4649d6bf593c575e469f83f59271453ed6b91d063c2c2f03547263af226b32ba31aa52214fd2c8cef1506be3b1673acfa97b276ac1b7448c639440d56f2880ff4b6bdd0e74e8464a73aa497e2b12cec24c15f3b75654ff4b2cb259116e9addaa3406c213c6b2ec66f103db8ddac58e37c6f49fec77fd1445ce351db113091cf28ac8b700cecb0cacedbdde7bbf5972cb40cd7168b0365ab483fabc46510661fb57f6dbcdee01f1b0d53667d1373f949de4a2c9627e41b634f82443c0bfe03562ee08ed40efa0a70bf8249b19748fbc87b01769990b5a68840cb93586312dde7fcc4c04b4fac77d2c8374a0f46cc6668b504429075379c2f024a6905dbf58e10120d58d3cdf751723dc4d4a39721dd6184b00611458c9ba2b81f9b860323d3d56fcf35c391592148a481ea139ffbbaa599a646285e5b966eee3538e9c1d1bd0e15c8bb913e1403b97e7352b0de990301f643b1505ba63c3a5015e12974ee02f233a8fa094691b53c7a20964df2b596e80305e8f2692e6567275c3760c4f24d8868c6c96cd02139fec0ffad432f824de122e2217263dfb86d03432b59d0229b097e7ef3ffb0f1f7c45d3a7d958df06e95fe26e4dba300b075477ba43a6845a0f689dcee0697b0c1150206b4b2ca3269c97e574558ffb568c654587ad5b6cce8cf31efc8cdbc3c8c504e8e13bceea4ca3da77d7b66220cf0353dcfd69fb1f984a8715ec27c2197ba8bcce0fb0607c72172a23232cd85ead3529b2d6212642dd5b3a6489b55eb6a18cff473e3188834d19bbee33f2f296e61eaea9eb2659721403c3847fd3d15cd05491f4c74bf040cd1e998cfbdc03be74bd3b68e25a07315c3992ad56df43b54363934f0c8a9b007f26075c377503e2b0b4d3686ce7eddbe2a56c7db2342ff33fcb2f0f46d73a3103337761d290bfbad0418149c2330f2b55fda71c9bc289d85b725241f525ceee35c98e86d8f79983c6b091c1f5b101944e5b4c7a2567462d8a4c89ae20c6953cb61e78e34cd4f4da793d0ad82ebf26a9024d6297f5975be9773bcd3ce0c95aaa45c002815269044d057d76b9bbf769858d1c291b29145cdfea67ebd71613ce2750314b5869f96803736667a88788f3d2224e3cc5f4749bc4f48934ea9260e0296e2ae67ae5b671d663d5aea9b3735a07d248280e06c0ae4fdd5ac0f49f3c1a8f57047c95c65b2b2f4168f8b2cc508d646901dcc81d3f716fcffa5b8d7df16481451590acc07d5c6ee0e1f614b5547a7cc8419deacee89528c472d886b0b471326504dfa5d5d955871a6a70e0b919784ac8c8740aa16fae5e7ec9774aad6f86cfcb6318496524b4ffbeda60503d58ecc959d4fa4d1bd492fe940e5edbfa54140e2b4eb109152c92e28be73e4b34a923;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h98035af0b3a7b905def62afacbff09f7fa8a89f0dc3033fabe0ce5f8123793d50fb496cc00fb2e08c469e9633041c7d3cefc65f5d580d50871108e291c6143dafa7403cc84db731be241caa132791241e2d1b0b7cd895b85beb496719b5347db248336838dcae71cb9ceeb4f95bd914bcd7302e0033e40a094e9031df35de8c1ecbdd386d6d533c6cc5ffcd0eda52e5512699782b80e400c5d7e51c139d7b028ad6bba6f99846f2f9ea84be6c49c9481036b64067d3e83684e298acd187d792f5f98f31c74ebc13ecf8f3ae7ef6df6ecd7b2311a390d49b39ec06cf40ce44fa19bf4ce961068e599c70b3a027aafa952c2ad8d96fa11f47e0d0bf878d6646dac7046ac10bef70ec5db3d1be4ab2f53236fda652047a453d7f2869565720731f9c0fbb80b5061de32530fa434704ea5575e3740b90cc86c368112cf6e21b3379e86a4b3eb29e597406d8bc8b7881af79d3e69d1168329e8089f0e439946736e4451aeef84833adf05f5c2d5f3116181e9f792730d8229196ae5fc80a348a36723f1495f5e614e59132eaff27e320461eb60610933296a45424d56fa3f326894bd0890f33473d293393f53f17c868de31277526ca052314fc16b7b2f8d744cad076cb75aabc468d6db83f37b83b771beb1fbd9959c4fd4ab79116d0d5bd403341a989d130d7c3c774578f3c473bec25947ccd5ea6aeac2fbd7f8340a4fa5649c9ecad62552eae49f93ca000ca846043d22caf762864d3df823e421308692d871954347a307545e1bb21e597e4801d16632677f2d8208723f94579df6c619957efedb07464a793a3f465342e757dd6c358cd98b0b0c3bde981a2e74754d2a9164888adbb6facbc668090036239b89bca13a62560340ac9d7d0a92ae3190aa85a8820e5c1b43ce245904bbd1b6b495f28e4b1edc5292bb3d7937a37ed15e6cc0de34f5779af4e8f9ecfd5d0a849cccce349af80138436206a84eb950b7238267a4b8a3e9ea36c09021e56b831cd5d437ff3d5ecb595fd4061089c83cc602776e405f8e963c9711b683365bcb60d4cdafba56320dab054e0f42efaa887e99961ad0a8d7e63094033d652aebe2c8b8a5933727e0f0f39ec24623046c36b685d3535effd6b350cfd30dfc8789609fea9c8e5941e0dc6945251410e7a0b6233b508ac907eca52b10b2193bb3c66c3fc20847249032e66e87bdd0b6119bad944b0fb203d3d8da4fada496c2d6d7e9e0b1f6dea9546797436c585d26d3ff95260ee767589eb5138580c9949c91091627b8f3ed210cf69a1941465019e7fc225d39e2e3c8f4194574f6d6db3bf704301ffd23fb675da7f02f12a6c782b2ccda4c6ab98c5439a61b440bb1131dede8f602260a890f09482c50d1145f1d208eaccec8d2c13797464003b9f9af3f0f05a9c31b9b181f0a118bf9d38aad7251d8b2ac41ef8928db71cacecf78f2f8b2a09e74304bc8dbf6b7a12004c6495f823a22d61a1ce4179969044f2c67080bc32d5edb775b4fdc4852aa1c74d00cca1bbefc138e46ef369a4629eb2ecf6fa7fae4b71d918d0a8b2585c7b263bc44e21e8109f391a8259c1fc59b2e6af52cc122d1c53c13a5dd86bd0367917e2c3b631c782cf92f0cdda3190b98c7ed06adc74a0718fabbcad745955c99bef3770cbf5eb4b89f800aff23972c38fe72b5341199c8a20d00935325f98d9609512b0fee69483cb965e2aa28de4db83b39bb3aa94f0f418bad5dbc3017c5b078c0677642f4d2d3d7cf13f1bf96e9e08e6f35d324b9ed74ed46743ca8ff3d7a8b350aff0a9e2c4bdb7221d36416d89d04a91f8cb3dbbaf228d7f08284f8f960993e86c9ef472c5baf80c27b76446d5d0a14d5277a0a9bef1f86150e008e3afaf59285233dd59ba578318d5c37d48fc4479b47da584709f145bfbf00913642f0d5e064a8ad260cc3976c32199fe8a977d899a7ac93032b30507fa14b33a7b9b3b7b618ffa68d6a0cab26fa45d4cd80232f98027d746711b9ef57c67e7804aca0df8254773991641288412a178870c3351dbd51589ab532797f9121f3b1ede317c7de8fab078d298f37ef96f6440ce51097e7e19615061e08437c112074d26ad63da42d1b52abf815fed44ff9c23940488886b7079f412ee167b5d79faaea3bbc74bfe4b5dd495caf367df9ce25a8e3d9e0b556378c1339cb7c16da0f417a109af591e37ac5524101b098978ab4c1a78fa56f170cb78d35b77be4c95946a6d0751b03cc755ee22c695742f1cb8de67738b5a89f226a5df1d1c0baa6724dffd186a52511cbea04fed07c2003058f6c6b368e428ceca2d497e80bd08845fddb5c335d8f68225bd4fe5d3f4a02b18d86e2f78c45b14c15833b28b2c26803dc0faacc2593a3162116e2e81ffccc52e3644928a794c9d1e9bc2754502e79a4c7000818488b02f0e280e8518509e7da5be77090191428c6f2e3d2f424c62b7888c6487dc9b4d22416796ecb102382db6273d0376a4ed58f6a137e3971884b38fad2ae967106987f3eb893d913fa51617fcdfffc46fed305936d983d2837a3739e7a815ce94e707761009440cb0ebf17fe3b3100e579b45f8c317efa00ea459bbd2a096b591d5322cd01e2ff846f8f7c709756aebedbae3f35bc1e3c82a2d69566110ec79e818a6558e8ef4c55a3cee631497b16fc3ee193a186ab6f2c0c3699ea3b0a12b913eb8e00a6d48e4dd8800d8db384ed89f544c3088803af4d7625f9c57896e057e7e2250b328a9c5b902087c87f9862c90a4e6599467c3e8c71785fc76c270566eec815158947eadb0572675e6d966d9110130aa2d720c2542bc678d9ede0cd22ac2b7f25e4593037a451fe20b3d46c6c3afc47358a508a3f3d5787884427cef660d5aa52cb3a25d6152d1db418ef457be110c35d2bb5fe4232ad76beb69ee571576ed71c754be86976ecae30e3bf668422a8acda73da7b54d77572fcad1e21fb03d2362467337637db123850ccd895eeb2ef50b6a280ec568e1eed09205bbdeda5f69bd938ecb4eb33613ff8465e66fc6e85ac833a00b2188d16459c0ccb4a0ad7f55aa34108e9c27a7d53a43d6fb35896f7ac62a8e15887a63fb8a07f3d506a81ccf8809375ecaef83884684790a891748030c4446809905d35b04bac15ae38eae854c5dd4ebc724879b1cb95a22396d671232709a2da42e2645137fabff41760eebf76b51740deccc9da7521298aa515ccd91f2105d483ab84acc68ccd1cf93e529cb700e7be96aad5464e7b329e5618f77d76eba5094e544f100082e35ed044f321a35dcbed6930bd0a17978fe42c85c1ddcbd6fc7d309837e589196f4854d5d4a25d84538cd49dede9f122babef0a6cc063057aeb4194a2489328146dd286f3c3ab356edc69abdb4cba620a2adc1be25f915c5f6025c93aaf89a8c8f2733437eb9f2f054dc797579cf2a42b490675e614fb9b8eb76e05ba015c1c0d10e06ff497596893e8c4b4a2a2136fa26a84d01d1dd68dec6113fedf06bcac0a4a89003c6a9abf94c275e6d909906baf6d5d42287ff58843676066e302ffb247f0e2261f7a58f1c27c33323a01a3c11a92aa3fa522288fdc99d4059e063132b4ab368e7ebd0deee5071d73c3d949410056c5334650fcfce8ed77c4ce6310fc4c30b6ccc5becbc989c9b1bda37fceaa02c8b400e1e81eeadf9f6ab6ec7b31674924cb024715cd716cab0c03cc956580f6bc175dd99cf36ddedb26923f857816535761999e1268a776c5d5dfe1de17937f2ab4c188b4956fbc1a473d58733bc25f8d8f030a39a50ab25d836ef831bc36e695e96fa27ba69eb269cd4ee805fa55603872a8ba3968cacf0ff2c5975d6b3b6333ecc063de5794f9e3dbc2643d1da40ce865dc2a4e6090e8c224e8b36504144e6e662f01e65aa74b5da9a681040416d4a1f3e82b571177c62ed0f8901ea69599d769ef3887f30b6434d7d9cf6899031c3366d6bd9fecca84eb81422870b71b66dc8c04b76b7f4d444b69ced90160d48e23690277ddbf44b5cfd07b90ebe049188a0756830be0cf9c080ca038ecb0e36b636515112b4ffe4df75d28ff47039a7156beb97c44f1c40d7043dabdc178af4d0533030dbacb0aa5d210f7d0d72d0740803e950b4a63bd1c46e83dad31def3a43fbae22af835337e58d854c36bce0dd2d6b34f28ab66cd93df0b09f27171ade6a0ac6939618c945e35dc51772561a2bf42f4e2b72a49053a43c96b8b625ab1df1a2b11434dc36c21be04104a758ed2ed08817226b09fc993d1b968a1038088134befa8503dc843e4a2a7653aefafc3094fd7cc23f8bee83a3a255fd184a45ca815bad81e201e604fe39c557d929c47b63008df2f88d0076c0a1b6240a1df2d5b743abb01da3cf494a97d4f4f258eb9582c8c9632b0177a56232bc183ec9663c3764181684507accfb7f1d51c7a925a384d44e52d2d954bc278f162e37eb87f68fd2860f453acd51ade426702e917416c112f9edfbec00aafacef8510a233ea790e03c6a1d042f96fc35c641213a0d03ac1a481f39631dde1638d5d535cdcf728f34a1d0d8863f64b46260c5e6bb40df7a535d24b54fdbb489e5d1b90b54ff0c9bc57dd914d5d671df368781d3c9d036d6e5c22022ac8f9ef316cfcfae46ce35d967b1cfde1df8959f6e90fa6c1569111bb74afe403a25120f9619897359fa8250f9dc0968665e032740aa7ff22bb9499f83245d0c2873586d6c51fac4940bd3556eda85f896569684be445d1617250a8c7111bcfdd22fbfc4067e4d71d0664c68c2c8ba2687b62f334e292d3b21331f3b78a885a7c278b1d810db44eea3489ac538dac9f48e4b9fb7bc884da267feceaed1e02a069ad444f57c0baa8ce949e40050f3f2a3340113308701cf3bb4cb1ed70175f2cd8fbea4e724a57f26daa3e289af1f72eb6db14b9d08dc2312c75f585fd91191e52ff923d019667bf73b7fdf0006a3fbb3637af3a848375a1c1b62e26ea1638b481e65de571bc621c7fc7b88960525041502685b8a1c9c28a6e123151230d451b3af6bb3be5a4fdfe1c4862508108422611a6f9c7474d1e8b2605a361a0fa1ff9812320a0f5c78da62598d2a69ac7ba56881e0b02830da0da8f506ee442d8f6d889fdd332486b50c12cca1438729301ca125ef37b636335813cc45b2cb5f99c9c227f072c991e02f0f64bd719f713482df6a40364dc874b028bb492738a5551656a9eb3dba5392502c8de65db38ced18c8a066916a38960cc1c2b569f943ef54deb5ee78d137b88168af6861091fb9fba257e353a429251d1597b762ac2ec09bb840b689866919681464791d231645f2f7fee32bdb0503e51491a41a5192bdad95338cc0e112f5738789a3e2986cfacc10985f9a52c6ef29a54c85d4dbd772626c44c4e99c0ec55701856f594fe3157edba4e45a6eaab504168d73b8cec79a7be4107537935d6610ddcbb8e5ef3d95ab7f9ba470129a974783878a34e580c9424139f266fa78846c34db385701d81e7f0713e5e61d7434dae097b01b3cdddce1bf086e9a28667eb9ec683b7656e1c1ca02fe3577238360042f36ab7f9cd627eedb34228bfea7c4e548add83fd015aad93768aaefeb71ade218d04fa6541c077199177588c678a221fcdde431c3a6ca8b82c3f264a860f8a33212ffc8fbd813f1e163e97f5e293a9549850cb0a8860f8f594d2e29e50a01ebd0aad5a78a015645b74970b27a2668a9da048f995617c44afbba549e1d7d73cb365dc8288ccad6fc27e0695ff28cdf8b48ce8bb6f5595d07127d8ecad76ec106f5e64aeb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcf727c6b17447829cba7df024341e88fd7ac5c4c23cf0bead00acdc857a61701e6266073db32cc36e7aaec592b23baeca27977f03e62fab3c71c128c81916f1bf58f0e21242dc749c9a2fc483e42586aaa21ac67b67deb01427d679274187b44af15726cb8356991798f6c5a54f9ef276c708a93ecfede96a92972246e978ae0b7c3ca0d067f9b64ec440e96ae0fe83dbaa023e018354877b161015f6da000014847ff5b0ec7f044051d7b49f1e771322b17f154202488212e66673070555c81f564ee2673b46d2d17b6c3380a764b802e603a4781b63c0d056945993101b2f2f5343dc39db08a86b1fd4af299e75cdbbf9f328f4860d5de54e660f1fd67924d2ebebfeb4939dca1fd1123bf0ac357b76f5f7844c9bb412b47c5c6861371ffdcc5faabf9db5058f93460527a8a8dce6b0c5a68ddecc594778ce2a471b8caa628ac6552077aac2987cf3f59f18ee931bf6d54fcf2ed2aace1908ed732b749ac7fa90c1b07b15bcf3cc46d02a1adc0f0513b43652ec5881797c18b545d009c1d9e1d4e61880139cf400e85586b3a3aae9645da5939c6471f362c6eb59d0105cdece62279f6bb9500d1de9af8e5600f6929b7ea86865a232cd92d2be2772b450ed4279ff36ce541762219e9c3f03201b442c5ffa0bbd5b4d243a390cdd0a1a5c173e657ea6a70712c27bf48a7bb3a0e9689119fe7a33fbf84110f25eb51d37c6136c25bbc885b5bf8259613edd3540747017e452afb105ae01ebb59af3f30520c55c66ba410c1cbf409c09a1a9c84c31a90c80218ff078cff985b7b00e2ed8446323264934345f6d627e7bf8e6929fb8fe15ce0c0ae6e2e32ee16407b9bcb68a81499cc00cc259691eeb31060010b82e9ceba703235d5a20789c1fa0133410d2750decdc7876bd1109583276a0cb55e553b69a74780595909fe4f9d3d6171ebeff960b595f921a274bfdce8b50f698092a807d5900bf04590dc5a095c359a56939fa65f4f356bea896b361d63c7f38c1666c7810dfb95c8f7d820a8e6edab7446c9fd0fdd46ef1371a556e46be86ff131713784db6f3e20f58f8432eddbfe139d2bfd3f04b58a803550da27b6c4b931cc8044aab0588360719e5e5834db037706a3f5443db455c769565f476994992eb5ae619eafb60a3732585d987643366dc0a3e2de76b3a570a0b4158cec3ee5d4f8177167999c2c503bda610d1b32cedab02b9f4760ba6a8579339b6599624715282a0e078c6d96f33a5c5fbdf07dabbb2dd1dfd66c9fb0d27e47df6abdbf7612d5f3dfdba4cb8397affd6d3d584b0aee31bdf6a88f7a7e38351a6fb812ead62ec9f9e67b09fb04c1fe34e1d6287cf3e8c018db487243c4c56eb4075e9129da54e2b7ac96743188c270c46e0b465b4f94b54faf46b202806467b00c030607079315326bf9a3e92e32fb8bb42f239989f11dcb0e8401bd5e01be248881c93ac552ec86a463e990c6dbe8eccb73715fb5ce5630111f7bcf048a339756c640e3feabcfb4c60372fc98c275c4c604183fab8759f2a6c399d64d24caa3b4803d925a4cf8791e2a8b899cf0fa7d2fbc5d72ee0cac1dab4e03fbd373c353bb114471bb02af586fba3f667221f8cf6ff60c182e1627b9809a7296f3db71530835196f026b48b7e06ef16d0e843444ce853c958a8612edfcac6bae8a38f587c0ee4a085993a4b95ccbdb8e82de82269429e28cb6e267fca116b7b98febf10251ca9d4982bbcb54bc48ce140de558f19268995d305f41120447abf414e9c541e69616d3a2650e0cb8d6a6ade347441c85b8aeec02f698aa1111423f418f0e175bdb40df13d7a68b7002dd2eb18c4c935a52476de11991cd3de01efd0308090b026814cd7d2de8623274ef149622a0c63938a12c37896fcc0595c2229ad5d143f86dbb36549b8e217c2e29800845c327418492922706ed9145023ffe6079465195354df1142616781dab000dd9ea08e6d6898b6457d634937e78ac0bab8143d7ccc8467c6110971b068acd5dd3165b8d38b1cca0efe8204255b3ed4376427ea6107e69ce2d85b12ed0156b7c1321be24cc3de86b889c0df01d62acdf9c88934a4e7931b143e585a3f121bc69f5264e132979f87c8a33a991daef3ed69b6377236560badb32d52b0483f9d08af74c0f335925b939fdb5184aa499ceae660be30d44ec55c1d4996ab3e671e22198bc3c705826f02d3977c56954fb149c69ba17134503bee58348549bd741cea5b0d2d8053eb3544a19bfbf25e1bab4a4fe7d7091af1ed1b9073dc8e2cbe6cefe9e6073c4ef574cb36e9ec67db8a198a738e0be3fba5ac9afc662c70bbeeccf6840596b731fecd5f10f6393430d7201c482d9c4de99969f32376d4d93602085594bd3b1c16bf8fbf3e7ebfddb290807fa72afdb86f8aa1163f87ce701bb389d7bcecf073b54f0821ae5684f59720ed9a376d33d7f354c84626240eca73252bec80dea2c9a9883e4a9cc70e05cb8560f100c2e89f7b60e24042620bbe548ff377f399e0a873b19a0f61983db7a4af443922c6d987fb51ab47894ff949af3680c230fd62aa5918c4dc72913f24088d281500b3839283e393a5224e5647b936571fdd0cd30b38c93d28013237b2117a8d5b4a4d37c96dba9533f972d392a85179339ce958c8f9501b25f761fe9b55f727fd716b9e396fb29bda5c3c2ecad240cf10cc47f966f86f383f2fd2087ab0c0cc7601cb5610e44e2365a2738372d8937edd99c35060395c135910ae54f6f8be7a21fc13d9b57f0be414bd94bed2f6ff244b380fb8d9f63413d0663dcb1621651cc29dae9ba02509e17d2b2c6c48be386ece6427443e93f976a18d3e02d4d15c7e0efec8899c4527808b0f27ceb00c2d64033b7ba42cdbbc0d04041e0853b5af9f5f31790a92c864dac49047882fbaf0d299f569ed0062903b82f9bf1d3b0f6b3365ca2957067556349c0654a459ba4106ec4a60e854721c5cb5ed9e2af8d0e46e963c7dcb1edb843b32555399502ac7c3afc4763916433a17945c73686e634b549654335e8cc7f29d0825a581fc145d5f26c354b35aa67ce27fef3fff8aa5e510ec26a4698d1ce0047fcf307f450ea9d7ba0ea49ea28cb96f9b4f6b936c28d12ac88bc13d2ccf4b56586ecda0a3a85df7a03a3c09fcdb0aa77071d953d77ee45edf77ceb1a4181edcb500a42c26040c89bcdc5edcd7ff10228409db1d69be96e1ea18593081efbe04e363969f7e11b6d29c15046a2c9dc099e9d22d53e6c0cceee8b75d7dd7d71ab2ac613db2fec075324e3af44287d09299348ae2577bce590350673bb29c9119002259052bd55604a08717834382877b19daa6551f92d3ff94c684d42c4d02f2b7a8a7eb54d0c98d3be46a3a3454c0e9415cec9b09d4a393c3711976896b0c9855380b46b384cc3f10267f09fc125a95eba1effe0bcc27ce373574f9bb9aa690c678af843003be8c622a354dcf714c28b809a2eeac5cad5bb31962d6676eabc72f2ab99a6154191f130fa12af049cfede56839022881a323cf3169b75f3280fb0cdc88c04b7c295230fda6d2be777b287b06a2829c99b545d9b29ca24546670f096f4e04ff70bbbcc94155b7f4650b65b93947c83b1e0096572747485f4084c10a4c30cca82b8e5492d5ad5b597b731d60bff3a710c71bc94baa101653e255617f712663b7dfe6c41e5fb1f2f2e5f1d82285fb97b9213b5ea6a9cfe70dcb40c75bae6c3913460c976a3b9bf67c12f97a1610c778c774bafc220705180bd94e63281e7e684c93731a026f43533a4ca3d0fee9dc24339a9e88b82a4642bddb0b777f1cec43dbc0c65c83b633c09211bcfe71876b93f3ee243476015c8009e8728237014b0721eb402043b7e1d969e3e793463338ae45078df8142c1cfe31c5659b9721b5b9b894b051a8ec69db45d9141bda18814bc0f9ba6301ebd769b95c19636391176de55a9436fa8bc37c69793ba808d63034aa6889093a270de3185725d258acd7435eac8e8f00a2136b0017829550ce305b11cddd1df728083824d0e41769a9a6420f448c1eb18f4d9a6097ef59e3a47bee787f3c5620d184a6c5e6e507196de80f723b56fdf24a08b778743de957e51caa98f041c1ba57c77fc00e50967f6c9ac6288af84b8a211fc66490e064d2bc3887469842122823bed008a383c0da9f314711d274b2d116a532d99bc0894c0fb844a491d4bdc244f770662383ec1e9ba449136607387e4246ed733eb308a6eed0fe1a7e890de68aeccb1e6930d71aac5eb3cb5ea5ff3ef203a89901c887c693ff59f40feba1879913dc21e4e75dd1c7e85836023e1c46b0826c71d98f645987a04a5f7bb8f64562f466b40221b0bb32a199bd7e2c0fe7aae5f85db93aaac9131d47c3d824420bb77724c415883f39153ddf4ca6133582c9683f175f91889eb62b6fa306ecbaa2a41efcf6355445e06151b79726426a95c2c680745e47461e4c6fc47d5aaafd18631eae7b5233ccee0fd50a4f541c71cf2c96e874a416e339677c58806eea9d904c84bc67ec92f30d30a7dcf9d701bc10ca9ce332d9e6ad1a56f2a6bd224498df507026e3af3f289ce2d9c4a3a3879fc975283cf299e94a189cbe1311e3bf9810aa385237cab86f5042c8c8359140bda418b568bbde3bd08cead2d08a0263fe902dea59cf5fd3e9d26b346ef409ee387a28ab68844ff678a1871d83892fad083905b3eb2d8c55c307b5bc7ea9df09f924ff37fcb05e8f2505132c45eba8987a27e4c931989f1cfd3474a5afd2240ba639b943c86144ce8d787b618ad983446fd3db8cd2ea7324a68612f097c6dac1f55443e9ecf5764a5439d76f67a7328abce651235fe96f6572cdce62cb81c36885f4531a6808977ae01aa6f2b7da92c254dab2076a2920051762ba61b317280989e28d94fd505b6c42958939ca545263540b38eddece386781e88246445896b701814cedf84d702a5512aed60c21a4f0848fef3a329ace267e1301f76e03e176074136595c48c5443c1dc2c160d3de8396d4c3d3cc98dd46b6a1ad862b4c76ccabbcf3c3ffd47f3a4502ad8bb06c679d36b2592a84d0c0da592cfd8e2d3a1d8a02761a4fbc32d8738a9a94a07d3cf1b6424fd0853f7ee4317acd33acdac786f521d73808ad69e7d38d5af78dbe226c0b374caae09269f5dcbf38478c7a3108f89dacbdd232655a454ae1c833b90567cc49d59b5fe17e1ea2d6979add96d365b76550d4040b2079544874ec3335a833709e11fcf8380306f3d0483fc823425562ea4f429ccac7a267231d197f8baa8d88f5a07935b17d04b544abca33b6dbd52f7218e6cbe1d9591f2470fc60dc09736a9a2670f60f3069bdccb2dfeab75fc59fbb2bb060967eb3b1d9ea6342a6f219ab2c5d3d8608857e538cc35a9cb4d9a64ed75d69fcc5bfe2426199a8c119b531b4d9262760d4b3b922f52f5c94677e7e4a9c84a782bc35463ee20eba709432d5aa0c81b9837b3d1a54a86eeef0965b8b73c09894a9d7173d3b8e0cbac6fd921e8ffe0a7f89a2e29ce255d8ffe2db6836be262d4cc8f08840662df39d789bc8a327ef028163e630b634e638d18504a0980649f91d3610d8219d7f89b51d78de52e269c4b93742e899c5194c014bd73914134249980753ed7df6f11363c2c928ad393548294bacdf1234ed8e7d4c0bbffa10f94b5fb012432b0ff3c60130480f2f47a674322827e57bf222a9d42a0ee4aa1007f7dc377b45ad01edc293046d4fea1c4af1a4f4e6fde3ea1438838d4b71bf04567cd9b285b85301064804481f099ef;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h24904979da3f1ee851fe867e0df153373368b7cf5161f179400e2bc4123a694cd001f57e097cccbf85aafd400d010e3047ea148aee9b5b061151974ec252d48a42376253fa8372da83d4132312ebbcc4b5b8dc6448798b12e7b6f0c7a683647fd6fbdfbc31385db3ab8fd5d3a4137f45d93bc7831b8a03eaf868978b5cf9a8a139173673169377f4376a83d47637b3a3477ab4a8e7514ffa797443e5b0d6e2787e5873753c3b4293493e17e408ac07b38588a1f6cd4cae2da2f545dafad9fea0781a71677ef02dd56b2c68b91c37884274f7472a3c9bd12224c84259816817ed5847bb47ff595f478c61a4db093f65f783f131511e1d6c0199a968485576af186fe191b6103d5520a5a586b100b72c86205f882bffa43b74a8255fad6fa4b5e54973937b35bf38d25cac76a6bdee2099202f7d35b0481d83c84d52eb3fa4bea800c8bd9b9f80e6d7babdcb09618f0f6847d27f62217d32955551d37e8c3d5fe170bf522c42164cfbeccbf9092c1c6bada56293c973ff9987470f582465b11eaba3027a569a3f94e9427f8d2d335e7404dde893ca2bbcbcc99f5b948f075697d85c4f65db37f968e8d6ca3d3643cd01befa550a387be3951098853c40a4834c437c4d27b485c1752a4dbbb88b7ca87b5aec3c7505c65304da1261ddc987592e01f845b5fec24dfb42ece6390cd3f84be4ad2310116a752d24861e79f7843679be74fb2e8447b4e9f1c57350457704689c484c3ffbaf6b598e5fc11cf00030f2c5572342fea12b668880d67378dbfab3ab5b4c457b1ac907509f883cdc9791c503a3de2367bf6f3a51b3635f08738173a6cee6e5eb818efcff551e58ba74213c7ae13d65fafdada6731ac74bb5b01af1914f89775c04f0af1657f339f11babadf73998b69adee43f0e8035306d0a372bc36311473d5acc8a05b69eb1f691adfb52f5ac6542918462398036710e06b97b50450e38c70f1e92ce6a78fbad8b4fbd6031165f9044f81c98274906a7c024bec49cfc0cbddcae8b31bc09ed539dfd3c416845bcfe31db3fbaf2fd073b15f1b881d4f6dddc6a15af96ec8fda01cd0ecf1fa1062f78176a2ecbfdb3751d65a14a6d958c5ebe0ce2f3987d986b953c7f4ccb08704b02e01984dec9d31df6d8a4e2ce7b66769b1e8e4b6a3000c3ad755d2a47ff87aec0e53d2c9933333a07e790775e5c72a8bbe273fbc31239ed0a54899e2b6c954bc31b3fcf59013c10c4882a8095e4c47135e691a5e0191d409ff77ce113f35ebfdd8a2156193ae2008f717e975035fe585680fff6f6fc54f239d0f5a586ddce3f96f7a285f5a62b0bdcbe8019db1f59faee22a76167075e5f38431e6f463c2ee065c60681b76384edaa34e49888e35066b7b4503975b3fe56aa18707fbb06fd8d2709f2aa18eaf32f535b0a67d0665c9326d3925e8d0a40ad58976b5a0da754201d7e3d7371640eefb0185403c4e1e32cf49c2a2570dcfbad2031a2945235bef5875c7c672987dce5e518bbddf351cced1b7856db21a5afc1c26ad1764d897d7f7c0cf94e597976bb2eb6113757d788e269cec2a08506aa91d9a9bbb075cc5897235e4a291a873534f30f1d0416f5cd99ef899f31b743d75d076d3febec9b8c46b3338f2eea65c64daa0dbbd341286f1bcad0769d05764c29bebdf73fbd017ad5fb8d6cae9a819aa1b3f78dede157a5395e155d70d02f790a848e0fc6cf599d5023d4c7a27cc5d86b610122e98a231d652b0bb505fe9919276e38560e6df6175b46a01fbd370df6e507079af328cbc2cda08b1e23348b44a90e75daef436f207b21f5454a4434910a3c58ec712d6c2426c1b2dd1b2fde64566bf60de3bb1f36b387bfa3dff8d49decf7fbb25788224932ffe4cd402b7ca127875c2b2d985c73998a5fde4625e7c7391af18a2460ca8c4fadaa83f7a0304a3ae9f711ace2d8af7bc1d783855e260918d552b5a0b248326b65afff26cb59aa3636596e606b5fd0d6e241f9c61a2d8f1be3495af8ad306e7bd0ba106092c0e00ec07aecfae76839a3a3a4a11b0a79213a5ec72b47d406b5fe60ad3fbd5727c400041843f1d8885d2416cbba44c63c453b8a22c1cdf17ee34fb562b2a982e589b5916716243c1af391c44656f7203ba638937fc1318bdafe9e39892ab80928a2758653d7b91b1fa6fd302afe0278ec8fee1b79a295a110ba02e5476e6e036333b05ccffffff682235005fea6475921fed2455cc038799779869fc535f787cee7deec306e635f4927ff253bb27ee8f927b229ff91391a508197a769de3a92280cc0dd1ad022c9385e8852073cb53001a17fd041dd2358d54310ab6394b4be41537806dc57d5247d332d0c21188f6fe0ff565abbe95339f0adb6e0a6fb6aa021e385435c3e2d6ce3c921bf8dc25ab8ba9b8ba63e064c620ce49064113e7eaf483bee2860875805619ac585e2a4137e17cbfd6003ce37990ee56db3f8dd745b77a7d916c2bdbbd2969e291f1c7876dfd198c45e7f4a543df349a52b7ed2f02ac7d90f8d292ce3587685f489292deaf8459ea5bc5784b66a72045f5ffb14fc131a532cd60fb6ccba42224ea64ec36a6f0c2fa48f23943d0e2edfe15a0f855859b19911e83ed5d1b968debb9676502737abdba301b27f26aad728d5e3c01e4416ef7b5feb1c383a0f0a53c45681fa92296ba860327d94d21c36a536d31a508f39dff6c0a937b74f7dc7303430e68f00ebced3dbb26f04dcc91a1089fbdadc32e06fcd94a541820db3c8000f360ebedac02b09ddcadac4a94b58dec3318fa606aa3f012ee0c2f14cb47d05bb9ee9efe9c2b1ea33170307716541ad391de6a720b430df77b7606e6af970f6fc47a9f0c28617e5d585ba25cfc07a437bdf399a3659fa83d122fded134746e12bc063894b4c87dc167f847f602836dacffc1d0a45897b7343ef88127d8e50749382234d53b2b28527bb4f9128887a17886a8fd6fff540adbc9ef1d0a95cffccd97f0b4c0f4a6495d4ee0ca7bb747e91e2d48a0474ec2267980ccb0b115c5803640571fed2701ebae640c61f613eca26b250aa0cbcba1ec0436a2d0bd4453d8373e4fe92098dcd6b946e7e0a30593d2a283cfad8e594bcb33f806ecb1aa3fc17db894a7e44e8e58ed19b6605670492261ca843c11f0f3f60425aac24328bf660852efea716c8865f15a563b914101b111d4e0826a75c37868d4217ee3b0ec7374c6f2fa4a6549b818c7421350908a053aa7a51a6449f48aa7ee551ca85f4855df573465dd2a5beb8d1c9d530d8fb39e0070f7de576cfc66936d4cb7e849fab10a92386a52ff7b86a26abf71b7f8ab8c6c88cf4c260130dd0d78282eef57fcf3062eaeb35648e82a1305825a0abbe6457ed3f00ebb99f876ee0c68e37976487385f6d33ce7eb6366f4091da670d2e4e6813be9dd992c1ba102aa8eef946f0a5666bac2fa94c452124bdf9a2ad840f6f4a552c5ac7a8aeef7d7c46944a3eccd2029f3918f71e43b331bf582f3ebb838067789af7a0e6fca34c541d8278872961e8a86749fd30fc199ddf2807e39db7783b058688a09c0e2f76047424400588f136837c312f87832070b4221bffe10ec761e44483c24e29976cd6f0ad5d0e89c87a8f2cca492d6e8ee50c6e57fa4e3669ebc2417ba6967584a0a14826b32f0d1e329a86a754b9f5c9fcab7e930c41e4bbb8f76ee8d638f87255c55fd6202dc70cd8160ff22237f2eb5b0124f96f6fd0473eadd18d3af2d3239ac758d5ad6196660b0168e14fa2ecb5f3469f115b358cc3af6951f28f1fb0e81d72de64d723c3b38705252e7f0a902c956e4e1662ee93963660ef4c15f8d0a14664c28b1774cbd1065648d46b8ebdba095305da549d9acfd795cb17b6763a261b4e3bb274795f91aa5f17a0b2e5acb313fcdb4baaa8804be188881fd4752cfc635a380b9b623e51cd4ff523b82a7b4626b47847e4208f66a9c413ab4697a87d7cf8e0d05e774079c11cc668a1eec38c5dcf42b6c5797e52bb462e55c2a944fe879a08df5464ddbcc743eca8000602085125fe47202001365bd7b41915eab2219e52d90b5f8a450a8ad46ceccc26740e13f3d584513f1743bf1fa58b8b0e63224ecea81e51fb5e76ea58cd13c51c5b355ddf800526a637647a69e22283cf54e8171a06bc992c7f175d646cdc94bb6e0a5aac01a513bf1ced3f0995062ab9d53453d30709848d00e3c3e501e941c64109a2fee481525386dda1f136aedb279e35174db1a6c35ab34a235ea7188bb02fe5088f0809b642978829ccf8ebb26a2960e9ee050adb0b7492d3cdaa9aa01e113279b55f0b9c49b500be6c688d52ebf94356a3bf830c8f722e69e0874b1a0ea8a406bcf9fce8a0fef74d29892aad14ba8816041548215c8796d8dc8a73aa1277d9cdcb80384aaf20a13af2a81660868dbcec7271f22388f1b4e449c1eb393ead9517fcf9257abdad79821e84b0c5c4f208d7e8204c0bfe5042b4200db1cf4ae18d80442522944525fb96272fd8b0c4d07fe508cd413372096d67a69a5cfdbb0c336174ed8565263514b9c90222a72c675fde5c7a018288f3b841d26d32fe1b93309f8c79fc42fab0c32c8efff73319c908d8fcd6cd175fa2a1a1b1dcf91ec799b728c824726a25e6590ccf0b873e8038691a64fd6697164c524e4a99859ce922a0795b8f1b47578fe1d053b2a2c4f956866b3c1f12cee0b7019c2f5e267ad351cb58844fc143e07641ba8f32c343c1db7f9258865462aa0a8785092c2f7964f46aa3c3e17a84ac9c9640a7c9237ccc1aaa810a1ceb147ac7aee08e26239e93b79b00cec8c38f7e9e25ce18aef92e473f601ecff8c33923c1effa6e9faa223354b1e24a92e79f2c9cd22d4f55c4d3d23ee7bda7035c5906a05d654f746e9c2081c0a830317d45d8864e859566450b83c72699974b5742f712684645bf75b604fa8c180e9946a043788f578e6d2ecba6b2aba5544bf4a560286dbbdd6c25d50cbde1a12e6624bba3021ecb52b8c3ed240a39e7c18ffdc2e3d589c63b0270e26c08d399b89d299803b5aabfe16a26170cb66f066c6813f53de0f4eb078aa9c938aeca6e233d2bd2ca3589316cc1c2ffabbe1d6e7095cbf2c004dc67a005944d9d83aa684a2fdc018640f677a55f7a43193bb71d08107f54be1bc6593210e77b666ce13e596482c7049525e257f7857ab747e31db6e190c8d3b3d2e828e684aba893db519f28d4f23e11a75ae7d3c21b091372312d91f62a3b2a3c5062ef34450cf69edf650ad99dbb9010ed9f85b3fe72a2001c32b97bdd6b10475d3097bee16fac82d15c1dadc7db4d353b6732183cecf000f62b3f27f5c60bc4fb116a288988d7be847ad536762dae2f32de7698c048bbd432988c5c1eaa0b1a8b27c079331912e225f05632342053cb551b89d3b5be627ceca2fa573e1a8d88258daa3da9fe16162e76da990ada353cbc8f78a6df5dba0eb5a55b56aea77417d0b0d56239d9df4f6f727bb40f975cc1a2f15bb126e3078e7fe0b01bc31da12ce5269e95a6e505396487a1dfffbfe9ac32a2fddaa8f5672752da9c20f59effaea2fa85448131d8568bb8f34f5acec46805aefc6bf40791950ab021f51d27e9fb993863500734fcc4f10216279d20ae652aecc25e5e3b6932409e768ad3302ab6c9f11143843d68eff7dfc19f574445892c42345b0184507b1f17688bce7709efa00e1b8985343ca41c82b4df649c72f60d744188b7a9f1c3a3f540d54c96439fc7f785a355631bc88a96ad62b38053f70c836de194165ba11dcf51e82a7b4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h716e7abe68de33f397f6d0db6f0894654879f07460f7ea15e5caf4c3dec5862e630ea5272eefcb173ed7c3c9324be630d05e8c2c66e0abc42ec551dd1998e0eb1575276401fe7b348fed42a0948985e4035f950b18354e1ee7f3717f802c76d3002239e570126f58577fddcb5c1844124db9208c9148095a9cf70e890c5fd22671000e0dc2495f72f0fd535bf3a13fe22116ef28ce3d3511e4a6786d2b1fe9d69821eeea4e347794cdfb3ce3496ad18f064506a309bce9ce57e110a671daff2d9cb837b2b520418f4a6997cc011338a7682f7428116f6c1cbb1996132f03b67cc20f36799b1bf4ae2d1827dcc7fee9a4c94f33dca84e1532599c1d1d9655f9e950416aa64b4df7018be738a4592eee0baa4472fd0cf85d1e9bd5a66a48ae21bbd8e5c5294778da0edf223b2f2dc653dbcc1065179203776ae5944bf0582d9b8599adc12ebd04567ca6043ce47d1f5d39173bf16a172aaf6294ad127f3fa29482984860e0a08ec02ee352e9ae23c5cf152999344ee1d32ddef620ccbad2ff6413c16f73f33ea040cf4144b36bb18c7c30363ca7d084447f05d7caf864ca9abd897404fc13e93262d29a7cb54023af54bb24b274f5fa6e8a21756057a19a674b523bcc8c5fe5e463a157e8ccc5776c8d89190ef2578723aca70ef8ac9984b3f49fd06d1a942b5562c8f2f5588e773c7c12580d0c5fe8b9ddd8a6262062851664dcd18a6260e2285e02c596867a2963e2208fec4731a6dc2376c267ce1bd15762a2c1ad321cab0defb3fe7e80ec53430d09b98d3b80227918bdca3395c895c9dcea398db3fbc6bdad89cd2935a42024e65230d9a2545092fb3b7f9a3bbed407ff45581a8d99a92874d1bdaf21422af2b9363ee48378982e19d16484f175464cc5d6d73a780bfba6cbecb6d7fd368a3e2c0b2091b2ae4a049a594cd742a0a12ab8917ded36242f5bda53a590211abe4168337b53a55f3b22693e85d43a8b90142ad042638dc9bf1295027e377c2ae7aa34e1aa7e93dcd5ba53a426f345bf917eb3fc28617d9dfeddd3cb08c7efb531be6b88ef6728ee60485d5d09bf3b5d271b747ae3fea353fa5ea765b545c2ed29494f0cb5269eb6e879cae51c41929fd2d23ac73599ca57526f720d1d5bcd2db656e980e9e5c128d1572296c09629b8ba908feb76fa878af4a7b9babbd2667d20ef5230307abba8889308ea1753e564f0bf0e6873312d347ce561a3ad66f041788f24d7e7dceb84189388e33d8d6b5017b2f916236b9160f8b5d4bd1b98896e1d3a353b7c4c2a8b19886cf023c716e0dd9c00310fd22385eecc83fdc3a6fb35b11ff22cac51d0e7b17794562b7fc25caaa450897a6c32cb28ea7cca8b2ed01e3a60c86010c320668066f7e998f07fc36ba93eef7bd5f7674a8e8d236aa92476c1839f53c5e26301f262fb0f6fd9aabe2660d1cd4dda9b98067c880d85be73d744f6929a765baf7a3473ee39eda58389240b84273d4d06cb39c82fc74548f10559cec6e71a6d3b8bc08fc9a53c138a9ba369886fb0a168070b04d7f4b84a84b86e3c36f505ae73fb04da38c42e1dc76acaf7cede154de14dbf1e2824fd710635711a5bf4857cd1c153a4d017c4ca2ba36db8c34716839a052a71e0293e990a83d1c37ccd5c363d6f9719c2d0be130d9698c74f136987fdc07c63539a0d5ec198a31ca35e269280962fe3bd7c3a69cc3b98c7c2b4409b3ade2dd9eac6f9e3515fb57d1be85464ccb38321f581e60e3b366e8d8a575ab9feb04e387aad4cde218610075c6278d8320e141c6e07994293d018db1d8c37bfbb796380915bc42fd8f8c50c903f5641e620732ade837f14c8875ce68ac43380ae76b4fe99c5de948ade694f1df6ae10214ed06f07d6a7d62c1c06256d0250fac8fde1cf7ecab283023adde16de78b97113857746fc6f2dd810ec690853bbbd83edaf55266dec0c22c4698c1cfb1cd2180092321e907f74617fa27df21b59e077f6cf36b3bff3cafe78f753bc5e43f08d0f810a79c8f04752272a080b3b916b5bbc71a10a76d49d1f67f8b4132668696d6b5f6820f7456bad62c7ad1c8681fcee091bd21b8ce5b0936deed7a9ca776b5d37f8d276334b4c3f3396a19bac657773f4c2e4dda9deb6f7a15fbd5fca5720f463c0fa432e7504a08e783552209a1b7c6a27f96fb0c0f4867950f6f36c41e407d9369478f4e17d1b7a65cbdf41cd3463d4f0c6e7e56174c9e0616cb3cd733833a359fb9ac3b7714a0593684fd135cd11565447061b1528327ebe1b8a29a139ba1b8dd220292b605b8ffd4084a90b000aa5cc9f66044b6ec32af9957dc5d1d273c1744a339620243cd378a9a47de2aed0b5e9ddda4217d146be5c795ed8b1f61ff1c5a35576be9581ed4d4a82414afa7365ad585d9d87db288a1c3ee4b570f45ac55a49cb6848a85528525cdb5307c8bf02989cda470d600a2a32731e068983d41f639b65d33ecd496f00029c253bcfcf4a455f920df01fc060b13d5d0518651f24d3e6753b2ceb2397512419621bc4751ab6bfc889cfde63c6400ee1af6c95bbe6c9714244e71d5922cbe565b4afd14a6b4a64a085a7d5e777072a575c84c41b2efdd5712a01eb641761f143522d89e07f1152fadf04836c711f0d711952b92519b6f5f545defdbd7f598269e903a21ffbefec33f49bd4301c8ef0b000ea0840843531e8f43e33a041bfc9c1f63431a069b9ff68e2ba5ca7089c882819701c262c9d84e52e7772ad43da58ab694faadd953a927b0d5f169430890f308679066fced03d4e7c7deee3cc7c831e6db3f21eaf6904e8db57bf75d26f835a9050bb8e883bd05f340d2f518c14fc9cb920365dd91423130aa9e22957fdac920c0a2d8db5a0256c9eb2c952b32c4830ad91a055af49137c2727be84b335a40affe3fdad211544ab6003c9d6d81279972e5904b170ef0540b08f7a976c0c1b362be6162e2418c91994d5d8d987c362e0a704621d95f4e4ba495b1ed8c71095333eb42cac36e355e93304f43f330322d794d5f95ef9ac78b77448012651a1cfea3d6f894b3010dbf027ef844e1e37047b556e765f159aea7a094d8473a3c088077f038b25849e3f940cfe64f2d2e7d83f1d08da36bb6f840a210d62d4031ceeb6f684d74dfeaed21ba15a1b112d1f104abeaa929c2b672a5eceb4e3e90526ec70e3668409054c165dd8435e407dab94cb42dc99b67fd12a06fbb098160004bcac463c736820ea98e6e3eaf6168f383771cba0d71c3266dc9a8d53b267417b590d6039489180a9f6d28710fe781ff5b5aee00c5f71643401e90ded0193fb1cab9b3e263ed1fe70c5413d409850b77ab4839f888edfdbbe67a15e80485184a87c46f9e9a50df570b519f7b1fb0c9bbf0aab518afee91e72817e5fece6d943a6542f7e46f2a4ee25318cba16c8c38be9c908247de772f0eacf571c459823bc8870cd087433f6ac14996e3ac85378a38c7a50f4e6fc8aea7df738b63383bf69544e86fac953fd8a5bbd97ebf86b69ba90cec3a9a1d6c67e34ce99cd3e73acb30bc93bd5c81303eed2151fb384c74241aaedce7a9d492981b6e1163795698f0e41e7b18a823011c986791bbcfbb745eecf39fb46551b233d725ad4f3d4fe83b9bedb662cc4d9632f5267d2499dc9d84bd7bfe8a5083a7a0b0cafc2e3844bf8d975111f0ab52a4de761d356501324f02811ca3ce7d568ac428c389e960cf80cd2729b1f5efc9f62e713edbdc4778ec5ab7916b0524f7d9657647136673404fb594cdff7f713aa6b8276fa2332d17e0e79b962ebc47309ae388e2f48267498093eef5e159f8ec7a99bfb06960f7ae8610186991b3e770fcabd3f5feeea4cb377d5939ad1fa6300cae99e392d3e82ba202c858aef1bc49f33d1cc0f062387e79f93aff8f74edd3b8257e27a50852f01f05b9ca5eca048a7126ca17c6f1a575d1a2e3fd8dc8cebaa5ad1fef0bbc094d71ff0e20e359dcdb84075d4ff0d836340ba48775188767d983621f4fac5c844db078c90b4a2e7176ce474bf5b333194ad9f5eca9e2f35ca852377f9ffcdf6c50b8de8361e70d50e725136701d95202f5f5a25f0ec2cef49eff5c3a54048f5836cb5a0930c6914cb654d93d36155fa1957eafac7b7c6e7b17234fa820ad33b897ff11cfb4992ec11ba1367027096f8a2d7f581b1a55ef900f21facfcfadf3b12f63d9529613a198fc02b22a674689bbcde65614ceca4d0f1e97e29360c0cf2d1c8be458068cd7e0cf33f2a8af8a4d1193af21c5a72f046d70395ed962644dcecd21aeb08bff25ef404614d130c8576f5d9a1bc3c1770da2848b0ea09d568450438123e8d27ee15d18f730c627ca97d4955b74603271514ae3365a431789bd4eb3cfb36655a78ee491fd6f24b25792c8bacb8b4cb60ccbaaa21478bc381b4d6f2d8c0a7460843314e86c4504f78f4dc8691ed27960d492c693c7647dc6edd31845d20d68615202209b22db7bd4cd1965eae21654586239ebef50d31b605d7e23dd14d6f8ce721d57aebdef0db3551a3c5adfd75dd229e8a988a012964e1015f04800537dc2a522325ce39bfdd5741753c47c460d3d40284ffba77e2f1ce51370b7e5445388370c9a64ab8a55f16c597d49a96a40475a7647add5b9648a0d817d0b78e8307d077ffa35178d610cd670852a53d3f6115698f00b8539f06c0addacc358340ed8a64109721bb05215ed0247e2fa7eb05afbf5f297c875cafd6667683070d77acd46c2fa3e38f59a46c5acd71971ac940ddf23e097053cba3d87b340edb8c4b381c9d51da6012d4670cf83354a10214e67513b4914cb00f412e2220ab5b7011d7309fdf1d48a3740700b69d108a4e05acd8bb1cbdeb81e0774dce547e91d5c3ff4d1adc7811a70d99ceee596072f4c2e09e61375120fe81c5a93c5bb01580c6cb4a3d3942194f6b25ee0669abdc689aea64074ea3bbf677bb84085ad464bb84ff4abf18b4e640ddc836f67d167e8dddb892f016cbbc31d598b8f7d89d1c0400cf62d561e234a58c2cbacdd2150ba28ed8f4bb3dd27b3eb8f9912c7b7940389dcc6ab34e4b3f769df1c34c1daf1275f565548d3a1c3a2200e51e386ee604976a8a135a495cc903329a01a38babc4da24ac1ca262e27dd33e1f3260c0760a5e3e991db41f399301ae81d51f83a1942c9662a692aca3dbfadfae2a3fa2452473b920738fbba880e3726f11b0c191dc3ef6f2b463dd186856d95396247145139f543c6e5a7a545bd7e25045ba396a9ab55c4cbeb02223a4e66ff07dc1a50a1c208b786bfa852aaff61b1f9159a16d3532a775f4285bc8f83e4e0f42279f39c4978ae50cab3ade36f5de690efc53e5f845ef1c9c008f173911aca055db641596505d767b3a5e5afb812f5f7eb04a5039462546c0aa3d3a2ba4cdf180dc6553c1183a8576bc752107087742a5f4f98ede1c01343056087d6eaea3b3e066b470e5eb6fbc8bd86d48c353a9f09e17abc8a7fdd4a1f5c58097ca70e50cc53880cc0496e399951eb403b78f345cc18948827f41424a26becd0743e99ad60a5ed45737d160209d93da8d41f09ed5f713448ff3fcf1d5c97e5d0771cf4fd2d12473edf6f9bb5f65e859ea11635cf1d574fb2824d3a5d633a778f186313da466de3edcc3c5dcd8bef0bb12ec921fe4b37041e8d1fa9dd86e065138ced0a93f681daab362d40f1790b49c6ed32069170b7bdb0a9eb7cae54de3c7f03200add9dcc5328bb40b1809134c25db8210c4612670b204fdc9726f52d30b0ce070cda204a9df8259726ee3a5987c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcc0e9d14a2dfb42861e0614ea26b63ddfe739b68ab8c605d24c997371421093b97f12d88a763c2175160f65f9a68c95e432dedb4b245ff6b400cbb4777fa94fa847c7900cfb4851d88357f28345b8a910a12a12521cd4d1b2b2bddadf14f25ac422435b91750fe23c7339c428f270bded338651dd6977e2384a6b5cfed12c6af1476df967d8cd7a2fb4ca5baf39e68b20e8b27bda4bab54fbbc4bf43c18bba2a0ff2531bccbf106c112992cad5e70957cee7fb049e05ab849f4200a27151d24baec48dc1ffe40dd3a38c8eab0c36904aaa18f90938489baef02709ceb1673db56c609492bbed80e9890cacc2dedb3096f552ecf39f9ae5ef17dc01eb319fde83a2e0d22884813a18430d15c6b429c82ddf9692d43e5f53055e1aa9c0dcf31cab80b856c1b80dd953c78cfc5de4c1380fda82687ed0a45442a571c4cabd12d18dccc6a4d0dfc2765a001629b722586484bd67b7eb4874566bf03a8f02f05bb3356fa94d90dd007be0a584d609774cd273fea80822d842ba0e5ab5910a9e871ef858d48ec4babc2ed4657d8497c609e6af838daf2081e36ce199d7044610e55e110eb4c198910ec7bc14d0e70aaf92c053227988e6a521af528142412af0d5c9348b9edcbbb008c1aeb28251e54e53473e6d56c428d4f3299edc99973991434e7e57df94ce14c3a54e12898cad4ca27a391f57e497ee4f28a66dd2e2af52894af9ac6ada8a7eb2a3121f252971e215a68d4acf67181bffe8b702ac4ae4f125a3510e2a0f825fb7c11ff7dccef4299d3714a0ce84d0b1b190b888f141a96697eb9b8097730907dd7eb542b8ba0a7762760ff8124b3e07dd6dfde5d52d0ac2ba9826e2e2d56066cfde7c5e7e0617c145fba7dbe127867f6d3a76375d9995c06eafc37d2327a0aadee57247f8e2696c399db78c348aab14913fa1668ed45ab51edd038369aebf735783f8bba7098e607f883349e6d729e2b281564de0e7055118a05fe560ca5104c738e1dcfe677ace6169ae62c1b6e224a1a0109d2eb970c4d7342e4ded5e23befd402216ff3a67e16bd5857ef1077aad77dfc6f984e15c2aa48d89584b15a0aede3947d78e115421446077bbf672a4315f9ee60b0a04e5e5d66dffe01564b8541225ac32981dc75d6783bbb6263de5f939947388d34510d4cda4646296f060d49e802842acfcebaf09f1a0f9930d49cbce57fe6dff41caf34490c1633d7a68b11d4f159d3e6a5537fb9d9989387a9ee98489a653ec4ad931b3f382be07032efeaf12949b6748aefcb2249cfd6b561f491cc8cbada07ea13d24ccea3a97d68f673f4e455b71889745cceb555e59c8f29654d1b7c0f029cb9435940170c13ca4beb158aa2e415ef1d7e1f9864f2c03c193e6db31b93259d2a7e528da36d3baee4eb31d4b90859f183ac56df9474e62bd427355d6fb3b1cedc4a3d8a86eb0eba2b337608d089c5cdc9b871a4a3f38bf7c353a764b1bb4909f4bc6d2fd199d0c7eb661d8834a8d9f16ee6cf1d2790fd4cac68078cd75bdfc0e7a6f74cb8c30ea67aaf46728dea2ca460c0b94fa9c8dedc903b5497c68268914090233f4a873b0018b52c4d026b24579cfe9635fa87652244c23eff46ba1933f1dcc17e8db484976033e5c45feda59e6eaef42c7c51c648e1f4e8519ac19af0738edb259956e832afb524d09868ff44f5941d67785065c097d80dd8d52ad13c91c6a5cc31f39f02c0f78cbc26241f613bb82fcb4f8c6787fbd3c893f2afccc03d11288dffd706c8b779720c10eb32b71473f1364b857deedce12f5d92991995cabe711313d3b482b616ac96337211aaeb58787880a8a095064630539a7e5af6ec03b8335161d13aa156c2ac1564824f6346d3626911ffe05bbd90d375c770d101228792afc38b73bb02e29b668063b73b355414442e53e9e95b65693ed231bfa6cc78fd8d31ab117a763d23e3c61b126dc22ef798715fb6a932b2a25191e4ff3362af5f63525ff5186d19e9fc4abffb434ac807369b2825403caaa65a62e52dd44570b7bb2148bd4295f0fdca7acd43b07d4caed4e4f29a2df9d64bfaaad04624e4eeadf82ee9f89aa374f4a80a0d09aa0c2933f808c4d8c9735b5a3e577021036a8b61d802ef7865c791b13fe910e3369d50f50018f5271755a9e6c9ceb332f02303f4ca0acb88c58e285c9d5e85b903a21097c4d75fdb5f3f68fa6f7200fb4e428092dae1e3be5170e5265dfe1f6ef08a510a76d80ca91756fb646f2f3e7e6694445b1401d8952dc27c448d75d31204eeeff61ae6318759b61dc460337b1fa0c241ba00ec5424e4938b5c70a31df7be545a9cd60632ae4de2b886777eaf726571a9e902d4b1b73fc7df8ef8b20cf873d55107477702d418ad47dbf6174d528b87c8abe39796aebf7d60841bdb3cfcc60b122a2ddcf3ab8a4db46db300df371032971817a2e69bfc06383a23ba403949ef228ece4a12bd55e8fcf32c2c95ac4fa3c5f846ed0255e98d48668a98c405c2d70bd295e0f5d0e5154c4b7478dee127375ae3143e96d6b92fb1f91ef38445c1de195f374f029139e49713c9b67a4f2597f4b084fd2d6fcd413d48091fa6d67d3d21ca81bf1d9e99e8725f4688c4af3c98713a701636d8ac6dc544f6acbdd979b1ec4ca4038d8b9bff19a2469b7e2fd0d8192d9f77ea49627c787622be9a3ae6085b6958eb9533ef72d608c5dd810f36801e1e18c529d5fe726f35ee77b5aa411c9834341832d6a3f32f0d072a0ba4bfd1200332e7efe274791bc6ef75b76007bedcfd007bfff396aacfd580ce82b342570916edc2082e16ecdfc1f640681152c82a8590821535fcacbb1e902f498acbf7f3fb25bc98053d516accdec508512b9f01fc7d9e791049624a56cafcab2e0cf73b5312eac35bf478836211a78c3a81bad117c910d695783190d05be3bbdc544e2ce84607cff7916ecc8f898e0aecd125843891fd2a8bd32cda211e23cb5a5ae7c8302adfa3c88186d6ba5a0003f1a648dd23fa3ef3e4ff8a72f01a704d3814485fae763f492aaed8adecebb9e1970a177786f9ff8c19b3e8ef84770927181770886a61c0d11bb19703f56c19ac8cffdc4e707404694c77b3d2f980a155a501c92aa3f8576a39f41393222d9a5d7491c5a29376d71d2301afcb7325dcf6b59d27e77f9d653b3f5d1543aea48913c62bfb950c314776a034b5a712cf06ec0395ee1e0aafe5c823482a1165b1ba004b625a19d6cc48291f186acd11b52f2878ebfe6e3c97663aed9bd7e19a11116aa01c77c67f71bff85645ab72bab2c7b43dd10d13c8dacbbcf865254d22b4e1727c738e7da585f8d7fcf4031b477a23602ac9af2ecfc43a71cc895e4793da8f9af870d60c7ae15c435802acdd200fb5f2ce389e4373f5bf54aee578fc8417eeb158510f4e330a60e988fb028b53665e17d7bbc6d11dbf2d8452ed7e7768bf956008c5f9cf630276135eab4b87d9d1a2df3203fdf852f60d228147594aee2dd0226fc85901799624b0e45a1f9c9378a225fc3fc681447c0f4621b3e60917ee92beec4c2182da95b27a36084c4dabda6ad75da32fed908e339190ad8ecbbf04e702f684bb6798ab080c3ef4d2de94e66b3406672bfd56d605baf633cac4063c9d82857373aa9d9bba89b1c9d86777222f78fb0d0cac0c2a85641b54e46610ae2281ce25b72d6e88373df4d33967cba6d2d4d6b36c7e1707cca1c559a36edc7b1870baee67d623867e02e9a36a2edfa306319f1b8c4d27e861f38139a7c9356b7c83f7f611a570e0a60e244eade8c79eef14ecc9855ae16b3e31df9cf7cd67ee12e627e2dcb74850ff23dbec8ceb5a6fc955f44133e7282f5bd3a39f7b22016ed943698ffc6e69abd0d7d19d4961688c1efe913d503d89808098df3905d608919a58536b874cfbb42c18676e71bb971cff4579962cbbd22fd4b33e3358ec0c588e794904646981e02b326be9438e49b04a86b3f405caa7d8abbae751503d845f277c34037a58fa8fc6b52ca26133d55b44cfbfc450f8af25b60557b8d2b83b2ee1579a6032d3bd98e3d4e7921135c6b3001886de37d277dc0474d102cb1617f3461777f5d4496a1d51b53bcb4197cc68c91de2eea78a39d37de470c5c9defd9b9421437bf7c6f7cd4a882f5ed2eb144c9860a15400b7e19e3f2d77867b23f1b7e98ef964c221420fb41ff36438fbd83cae6e90b240190029d5c83746901f7012d886ba960e41445766976c0bfb5319fb6622e806be42b696d66d055ffa2ffa502faf3113b94906f3c5a042498151a9ee42e341a974ed8612ca0f23cb29ad403ddc9c994669a9979a04bae4cea8a64878bc5cc7baaae3afe3f8920aad3348b59f06407ac19bd92759305504e624a5af7a66ee3378534ca25fc494da8831bb7a28a3c9ddb7f3f9b218d1e204079f82218342fddee323c6ab7245d81df0eb729a7ad97036ec8b9002c7f5b4a0bb628a127035cb171a6537b425cf65285ba7c2f78a4fdae41171580a549f078222e963ddd7802f6cfe49a55011563cbb005910f53780d490161610e2f55cce4ee730edd264f2629028f15584dcfb868adf7298c21c773dfc980979705c7b4210b9e893c2b80b61f7259fa3cd9fd17f10d2658c7ecc197a94251291d3baecea429c40a4524a6060847ccfe4c59e9abc0bfd30922c9161321368c0b215f5da7247b689c4a89602e69cddcda8a8eacaef55d8ba21a4a61b1684419abe3355149a30e178c7b20760b3adc6a3a02b8db9a3ed9eecdf8432b6d24e477f7f185f68df38eed311b459c1b5f7fd54e0a088d09627130a0249ad7751d6affe9264cf77fe1c422dfa92db044e07664f98b53705316ab32b72e103754c9abdcdb68f3d56ff6bb5d0507cd29b32cac7ad4e1944a403f6003cdf8000b61e296233e5b3b4b73bdcde4e0213173ebbf957da2c6b4ddb2380346ccc45ceb75d9d55e510d0b4b140655db1b57ae8aafcd5f24185cf97aa1d5aec058734ac3b42f6e00915eae3eb648c461269738bb8280475b04f1b6c9870f69ccd7c6aa885c468aa4d7d4d169c2006b36cf2abb2d44cccaeca19e1f95bcdeeb9dc1888894d130745a27a0872a5ae76454a0118325f3a41865928fba62010061cb799abe4e32d0f1953f0866a8b4246f55d03a4f19a18432493871a97468a4a75d1493e2ca0b55ece9cabc8bb4ab2de0ddf8e7faf45b24aa0303a89d9f450e78ddba8bf2953236d7ec86a219d33f0578d3bc39d6d702efc7a452aae88a2737d98c909461193c4667bd089fc07a66e5d7008c56825f45094895ce43b98b5f55d411a3039bc520e554ffc2704939efce3065a17f8d997b411ddb699b7df5d2fdaad66babeb6dfea414a67e6e5e7abd40e8caf4635866554531af45305b34ba51501db56fbf32d2119a33247d139961cd1840408bf5e5d71f2b9c9cb285c6b7a47902f40d2cb6025e74e02e5872934d61e80f378d5cd0ee49467cf66d16b9002baf3f8018fc78624b9ec93c04f0970c970dddfa83ea523080fccdc74b90cacf984148556da41f25977ef3801f70ba8f6a4f3edd9c6732b878f62e86ddc16042e05e7543e6158bce3a92dccb26516c4b3f726d6ef741dc9abf4d4dcb47e9ed57c0ab353adc4cffc5d6878c8bd86277597c2ce4ecfcf6cbebd9eaf384dd608decbbeb937a3d9b25bdaa301e156f3270374b49eb291496b2f7d41d66408b7071b1006b3648a8a11fa738d6c5d7aa8741208e2c82003b6571ea444cfab668938f4a50307da96644260df41a7ded422315d94c81d03e07770a361d42285178e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbfb72aac702aeb4ccfe4b5af16c94c6892547e3157f2ed9fe12db1036633e9969f3fe25399bfeccf6df8c60a53c1963c2cf302c1890715508d08f50b813903f11b9c342e26ffb03e202383d0d32834e623d2cb751200d043afc37195e3c4cfc79356250cc77a8e3354675f7e60a08f32569502a59e6497abddd81b3f0dde09b14f071c8aae3d4258f1e27818ff9eb4c899baa72c7a4f88b333558699cfae79aa8d817c4775ac8455b7911efe9529333bffa4ea32ac0f5552cedd158af7854ff204796a9aef61dbe5116c058172eb23c5b688409e9fa62e5b6696ef4f113e00d6a03efc60d171ffd9bdd3c0322077f66e0cccc4aff48c0aec79bce22487449689702df467001159de6793abcf762fe7c57458dba616163dfab496d304cd9087df17d95d239e6bbfe43f004e5c519065d73879bcd4668e94140d16f4755d4c7a2237efdd32ad3a39bcd2007d0aa22c5f637372f8124f812b7a3206f082f8790d7aa687ce4118c5f0960f43f5c12b5434fafc4831f8f54c46483e73c4d419ceef4d92e3c2386ca1ff98a98a2c391589eeb1e00ccf3aed81a78f67398b09ba5dcdc44f30fa6a194b86151166c2fafb4578d201d4748d51da44ba915be572216d4e444a61a6a4651a1200b17f2882ea7c897e3160062c25fc03f120b585973687b19b5b8a0dc62b518cc8126f08807589bfeeca067a30272da5785c90342f6c9b08c17f3bb772af529d91d0b200b7631fee2dc1ccba97c5a6095fce8a31efb1a1be8251d2e9fae22358a6ff8b611bf9ecc9f8971353939402862622e13bdd2ff56489bed442f43069940098c7403b4e5ae244a30c8ca211c016f7aec93fd1842d4dcfce1f8ff9c86ffe3f5047cc0ef805ab75d53487c428c33500e962b5e16d60fb68a4b19b4f37a468c62e52179c9063633b7c5a98d6f81701b71ee03cdb3687ffe0ccad49f2a688344b56f7218138cd7b04c38ad13f3eed9f856a69b1b8310ea07977ff20e161b059050b48d217f16c80d5685a019af60c4dda6ce2492d4701afa91c46e2780fa3fa62e309f15feecaca953260cc8304eb0439ce005b90dd32921b96d01d77551a1ca8d72f61e3d0363db2ff28b1e41c6b7f51292bd5b08e05ebf1e8638f3ce2ae690c7ff591ffeb5ba91e741971adc19ab71496070fbc9810bf9555ef45930145f5de74963d55ad13e07f0aed29f6c7425b0767989a1d2405f23a997f28a4d5dee590d685e0467189b4badee74b4b59212ed75901122aeda15573785e1753c179427521491d816cd27cd39e58c77f51265cf916c785a0d60783934a4266e0300d39bea7459f195d067d5b24b60fbbc1ebe13e6cecc49fe3fe413f548fd509311cc440bae06ea12547ee1d876f123a7e7ffb97c2d4eb7db7ddd0f1d50391d2e3101ee4f26ed76c14d61433838266176be0ab1c8a630d133e5f87c78277158362d17d7e1c95af2db45c56beacf3d84796c32220af272a57641af2acf6d5556cdd9f93aa1fdb854dc2a9268d2a8772261ade0fa7d023f0b8a066017e483394b2312093c77286888bf06eb638aa89d26c5b23f0ffd72eaaddd745885a63c053f0eae942bbf24d39e3cbc9ad8fd12048f244aed82c407dcb68f836d57d11aac42789dc4e8d23cbe250994fe14004e0bf617311a57797b399ed216dea4a486f20d7a02a50453d8c4e7b8490a6921a1f1abadc3e5f3fc87bedeb22c8c8b036d33fc3edff3c84fffd36a81f972a01f9cf4e01f6df101c06c3570054428026ab82d246f3df472aa989aec0f12f9ee32214b1a35fa3681dd5cac978d85781202e6a19998714633a251d08f8b797119e72f462856354f057740629481803cee4ed32d9241f0e746fd68fc8fff2a80fb6a27a7b4d9335b66a98e9c37b72eb88cfae1bf256e8b37e6a124e682b3d25e75fe6dc441d3394f99bb8765efcf4e0d74b9aba68045ad3b485703f7775e27cc5a8f62835c2f565a4de69dddce0f9b5182dafc35421af8f81da1913949ac315a302bdbe513ac3322c9f622424c195066d988ef5bd3b5b6138793da0103929130a75dad2004b38fb0384c12ba5afa8fc8412c56aab9539b14356abef0318f9fd8c3d6079059e728ac4055d5be4432652e4262384f6564ca91f9416f172a9088f9fb8021ca2a510f6f2939f70e161be938201114c7cbec8bd2e785f8d9ba5c6b81415c33893657ecf50f3e4383a13df457ac544dffbc8c78d2100d0655c9bd77d890647c47d977f8f44167e89d48877dba27da808cea3ff41dc1309cd97ce0781edf52b981101c94700842312c4c3dbc2ca8a4298adb3b093fb84ceb3a4fd2b0cfe79d681092bdbdd612e75c99e4fd83415bdcdd29d88bf434e6cfd1f0c0f2953c267f7cb41718052939988e938b1eeb1b142a3d0c75295f2a0bd74f26195e54d2fe4fcd0f88bfc3ad6da075e533d40d0a246774a5085b6e6d57e68502d492f192c9eca77008725228225545235b425c8b5ac64ed0f4e15fb945a4318775ac27d5d1b3fce9f1df8fdca491a89a5d7960074f038b96fe27abb5187b74de67b7c20033467570dfec28ea89095de8cfebb15ec3c6d3b889843058fa420cff9499b6150ef66ab666402bbe091c5d33064fc78eb815939f0e151b3b43b96b47b90b133930a90bcc70982b84e7641492f2009eb53c7508e74283fb41c4531c13b26eb9b9f42001a900abf301edbfa962c2bd536b21c0587f75418d27a141c5c0ff41f31f3ffa28f758f217de35510ff9b29c16e6c8c2d660088c7f2f0f9a26e554b83f8649309276f19d06304242e98c36f945c7d3e06430bfe8e3fd615a612071c846a81579a744bc7df0bd0f24d74bcb649cd135086f976b5859e829491ff9fefb0a04bf47823e979611e82ecf291d9574bd73760d3262b62fda41823ac908b63e081b0df213de647d2f4e99333984608991d69e6140cd6f4f5eb9126eb957a10768d992119cc9c7e7bd405064971ef04d5094f0d7981987f480deb4e6d3d73c88d1ba02688f376dd8b694f678176e4444ae7cfae89ac7ead5c22d86ddce8f9df438bee1d200a5e7594c2dfb2e66c44767d0ff1a5a79a67dcbe74e00a2836267c9becab3cce4a67a742899e0c2a8c28df406e7630f308fcd8b8d8426e1a41a00e622877ba45ae5dc6bfd89bab70f70f7c58ba30e16bce3adc3616761f20fe342746c8fba48a28278c9a24633786d33d20bda46a3f055324e03b1070ead65fbdf785f8475467f18d96e432e68224ad1a6f439a49ad59f653c1a027f3e831a3fca86517a534ac05821f86c517b40b58d9e70446be13aea06a4d908d46d0ac99bc702c3d549b06ec67ead7c8860757681498bc7dd7a1bf434b31af00bf4e81defd17d641011b7da3bd64eb8c771660975ef1daa71abc1e20c464162a47aa117b4d610ddc1e34741b10ee97ed92e895f98f47d49c05586193596197224419da094b73a7163194b9503607edaa21e11494f4618b88df8f64259a47f5b66f8833b30a3a6d2a6545e60db4e2b9a65a795af0c7e3e21f3c596d2e1f94d89349690924b9cce6763163f440d5a49e024c7945ba4ecaea45e71cdc559d7955d55e87cf52e10469e64382c01c0662c1c525fe1580602c4ec4daa86dc60ca2fe2b53b8fb4e0a891a4f1b0f5de626dbc6a56bb13d9077e63e2916a6b4cfc586e5adcdec68901915ef8155c1bb986fadd837c599401efc88a49022617f66e1928de5370b84b305cf1d9b59a52d6aec3af1c703e160a573dd18b7f73e174c9c33e25725131272838cc91a102ddb97acba0d2ea13c63180ea7e48dd9ec14f52449b9778806ac90e1e57fbeee13953971b81a6570ce453a7b9cddacb34f50bea2c3b71ea0c460705295a77bfb15956b485e52b6675db9e30c9f1dd9c19b2945c6d6cf58bce6ace26ca6afde43b5902002efae634dc57778b68b5a054bc6e79891f22640f24997b13b604c0e3e93518fabe3512dbe5c6de392a684be11e76c8a5ea3265a6055ec0542a23cbb77cde15b802e434ea6fd7a20d0968dff82fcd876a81f4d66838239ad2b21d2267fa596d78c1750aa57d6fe07ef027327d2be4df7ae6d3df2e85c990503756b415f793dc0f1ff16912c722e99df2a2cc867d40784555bbde28770e27b3c9bc3d3f86ff0cf368a783015dbe8032fdcdd25c68fd143529b3592ae318e05a500e21418985ad8befeff366b5abf82a2f2345b5230b710027f360dbe3a55024676e89296472478aec9e43d196b097ada3f2905e42525898942c18bcae1ec350cc863ee4613ddd3ca146459cbdd1c8927546739d931c836ce2e5dd511615decb136c73698ab9c8b5ee36bfd5e5221f29652f0726209492b83ffe7336d9604c047be0bc9a1c6e4edd15bda1c5e3d957843fc07c0233a3a77b3030cd66f57f181b1606cb16ee67c71aa341516ab8a67bcb3821d4bf063a5ca47e83c36e19d4a1bc3682f7f4e770b49614853bac3ee58f003281ff58bfddfd1bcf95e488100d631d03776b4f3011987974c0ec0f372cf8320fd9dd46d706b5e25cb032fd46a1a50ee072c07366c6b61c8c111d05d0d97ef2c98d54645f7da765e8c4bad6ee22edf96905157f803b63a62638fca98aa9436f120a46738f914ed65f2094fec9824ae1f436a26d309e6ef7fe0a7db4512c0e063189718127202a53418c3a82dc77c19bfc37c5bfb2521865e38998d7997844ed71923d857961c46faa94372bc747e6dd3ade07a672b1d685c1e740863bcde5a4e4af7aa00951e5b6d165c0045a3527b4956f3e8e57f34550fa002513680b86f567d1c433672e0cf97a1849bdae6f143ca0ded0d0c70e8de8d6997806b89edc8dd23c2c4f73f66de7ed0f49d805bbb7391dbedf675fda8f94dfbc018bce0ea7c0c65d950a08c25179d14fea340b8f153b6283993f1cf9fc2cf6456c1e5708c69e73b74854e5e7c8a3869624a2e41b4dca227c89c70f971ada15b374be216c68503c7fe51144f7b69ee84f282b8a469ade8151013f3dd1c39bd1ef7d2c4d191e3720d83c9aa082fed81400c8365af8e6974c7bdc8c42e9d93380a814668840b6276a792a379dc6859ae3dcf74cfe912ebe4b8fe92c66d83d97a0f11237f9146be8699625ffa3c81362d3f12ca031707691d54456008067509181a841b607c4a2954768c0400e43366982e1706e2d97c777de7cc204bebed5aaf5f149b9f8f5566d382ce587698f4efbbbf1389b927e71b4509b11a92a28b85553e6c338d6f96bc16372e84991d7746a1e52c5228c0b888e74a2a12d2dc0f0a081822436abba471aea99b7d90ff6d27898fe5e2e538d9b42a754d227c49c83b7983cbc04ccaffc349f939be92f44f5197d22ffd84dd4ee0acb61011c4b0e26392bbcb3c13eda3ee8e8eb2da0d154b438e409b9956f7e102a1fa67a8eb538adbcf274f7575ea4f87aa3ba373eec2c676f39c9711165aa27c2088e89cb35e9b914df105e13474012b34fe78a4cfa8ab49fe775598ef9d43b25c9892016614850a41278eb26b40c4de7fa5d1b9132e6686bc6eb2e05d1d707f1ce0b2c41e8d0cd569cbf32fd9aec912e5c8e624ca3f524a75723af5f7749e74d67b0c3c3d9e629e1111b698c4f12aa8253001947ffe07f48e82aa47932f6be361d44bab03d3269af4b16fa4ab906f1c384f96c11258f0766c30279ce87945dadcb3fd2aa1e3fc9618e1927a6155d975c6748e7f397546797a85fb6039d013c3d60ece264c05b09fbe3bd5006e3198491004aeaff2cabce0f52fa767e1eef16c65d6a4ca40c3310898163f34e710d303554e7d471c6e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1a57e359c48220e96b3af3ecd2055125818885d49dcfaf6f519e84013b28b53893dfc2593cd358b661f9d6eaf128490bed33e5f6d82cd7cc5a03032d3791c80aa75ca262027fb78065afeb86c6adef51caa8480d4d735e0ae3c948d3df411266040b50714daf46dc0e054f38e1e8c2b5e354219ab29c3f1b12191a4078437dd7cb80870b2e8b9f43bcd5a44c05330b51c44049d7e9b717125f91491c42ecebdff876882a60311665ae1a40f47cf1b7fdbb98612accfed6407d0846e300026a478698a300ebffbaadebe370cc2566529014e0b711ad1b9105df3b3fc7b285ddd1eda29e2ec0d4f98d17e1b71f1ac900ea565e53dd21ebfebce9558023d7e356ec529c589ac76aed6a287840a29ff596863ec61384b5cdd9eb146e814dbd764989ae88514315af592f2ade9c97cac1a26ca8db400038b2e0af8e746c8e40cc7cbf60984b177523818e3f59566b640ab82d92b8320cd10c68da1e8835cbd67665b9a2804dd4e74262d2dbd4ca0d581a250b6b040dec81d85bec21ec8479e5656d4149be66ec5c3b2629952e1d8b7f84e1b8e65bdf34cc7301daf70123c8be1574b8ab4a0c2b3606e6165366c3d11fe6cde4f7b936bc8df9b1b97c2976ac16a7e6abd502940bb01937c6cd63bf83e4af3cbbe54846a11c68d76e63e2679bbe45984ddd3915308a640f962c8d619e817fd1ccc12600d806b7d029ae97ae5a02b6d263fc4813212e71cedb3b595b19b8fdd315ecb88d3a41e8dd326e4bb50d909d2c15c5c4a03550a3d8ad1c47ebcc8a4a22102849da72d25fb2105d7152198464c73b4db5e3bfae8582f7ef7e54f1cc1b6bb6a349c80c1a90feed87c2cd51b53bf188eb6d7a5ff459181a99d8eeae6e4632d29e529f6d062919a51473a5cc38cb491ad576039e728adade542f73b72642e7a1279d8d5ee1f4b321dbe8eceaeb23fafb06fd2f9c78010b89974616feadfd517fc45835f4c056fd8b82f93c6ba82cd5d6ef52bdd33a41343f2bb988e2791c66265c4f73e9431d752ad1c5cfaf8eb50d9cf98d97cce58c7f5787bb3fb8043be167fe5104dc4c8cac3fc7196496725e8fb8409d795f9cbd4cacade6c494a1ec25a0f972fe65dae410a69dbcece4433b5a365c23f756de1944f5b65dc6269aa7dde18cdae0a64486de33cc0c28842de398ead11264b0e0d83a8f2761543ee2867e12e09d10b6a23cc485d70eec0728175d7ba67ff4c80e3641d1af235f7d8e4c811ed7d4052974c6777214265f4c7f040cdc0c2c48e4187ef455a413d8ada18e699193d5cf525df772d6252a49470c10f53f9265b972deb6d9d0417a7bcd2ccd4cfdf1f64b192188338369c717116e01d55310a34ccd482f27b3ce865e0bb907dfb98f7a3203ca2a20f8da3f2c6e47d3b99c95ec1c75e1b590353cc8b667bae736eb39143e48ec18db28ee8aa296418d2ab80e8bee8cdd18834f67564e295ff59178e673953aa3ace49c99c2b82b8ac68785ddf0797e0416f22dfc4902e7b07a96c099f91d33ffd73fb211c74e64980daa11c54c04925e5b9d39eaf020ecf9035290270451f3c8af071a3c786b5c150ec0766e91c6e2a6ab9a8721c141b7ef9b51521c7409316c1ac7f64e5833648e15a5e8b10da7a3bab944d2750bcec33957e8456bd69b8f55c7a152a558bee7e6febd17df578eef721083cd2dfefaf72b7ddc33f5d4b26a027ef336f9197d68b10caf7eae34e80098981c7fd040c3521b517d5d835a3d3fa8e4bda041fa207c2343faa2bab03ef2a9bcc17d33f870884c6bac5281ec02e09b961a7a57d6d4047a4da83bd7e3ad58c1705b1cd8747684a3ebcf385f2fe4087e819e387486437da644b5fa980d5ac24b6fb6cda4e272ea12532fdeac50b61d8a5b99e136510c974cb422545ee10c02e1d0e249fed88692ba94a6b3761fba984eb1958d5451b5c0bfc08adf4d5ae530eede2c7f086b588d9032f6c7b88f6af602127eac4a7a1beda63f40ccb004eb59ca594e0667800036a803f009e63247bad5642a3765bd7b0428d50b497eff83773ef85d4e135efa1a1c383fbbcf3e0f7636e42e049c665f7d379690aca822858b531edc7ffc30faaa40b10bd03fc689b0ef9a317aab2b2598a97b7eb92d59adaa9d49f8a8830b1763097810141c576f4fe1243892a75452ae9845821add044d949e8cef6619b339e5340111c12c5f097428a0b488f6d7118969c5f8bde12a67ffac46c50932cdfb6b67eb8cf202de6631a1238f64a602461023e44cdeabbc97ab6bf7f6884d00ed4a9ffbf5d2aa331e1005d65fc6386915f7ef34f53b8da9f2b468ced5061414b1d04e1e59c16dcac8b77242c67eac5fbe47601512530dd9cb7b88107ab2a114c4b4a3e557f450058719aa1b3f2de5f6c1fb245764b91b1f97a600f4acffaa35f2434a66165c301a4d3ee5052fb749ebf89a84e4e205df1e357fa1436e50726a68a42a7c6a49cf3eca1005b33e56211838fd6193682e783c5e3434b65ed2b83f80c59432918d2dc1edc161e22ffdc16cb120c2b891c8f0f1c9db6a049243d3d6b2cd13519b18fd522077aaa27cfc4324747d8d7739ce29b13e874aa146a4da02e03b4e30d11c46feb42bf27879aa732a4eb46fed1ee211bc6513838d033f1e584f622a8d45be67d400243b06489b6e823f413b055323a8a172749f1c5bf3cd683398816eb07986a73f74fce3ed67e53bf2fcf399f4c0815a1539c7fe0a52ca8c2653d2d4a4a2c0b86e9800db106cb1230459f70e29050d4e98c9a9bed4076487b13bacff9a0ad27d60bdf36b947a6839684133b92ad3d04b8dfcf4deb2b190297c8fda76836c1bda7b00adf0c6273eb757f6ac5ae93c7406d4c33b57739f712187b66b7816d40550a6d333922f61ffb454672d4ddd4a18f4c472f02faed9217ea939bbe7264b0212928bd45233db42cbe5f87bf8e88fb6bcb5caf74e7d1ea0cbe49e8366bc19d2f0287b6263de2f34edefd3a13b3ce6c1319ef3a82b75da5abb9b50960c01a83e1e91a93926bff1d7c6d55b326d1ba17cbdddfaebb6059485494598c3b2076c8c0569b47500f7bd84a5a0e76fa4dbe4b8af65b5250afca2138eccf7a93d991ac4ac36e644e16a510d2299d9e66d8a8915c232703ecbef18e57b40afdb8f4ea58a109278c342b68fb1820bbd061055df42a9080c96ecf674fcd40cc4e3de24194b08eb0aa3d34d95901f457fe9d333d582de8f3e0c99de183145755803a1e536fc059323de6f6ad928748283ea00fbc471a16148008aa5a2a7e8fc440df6bbb5359ce8bdf6ac25739652e47180e7f46b2b05085ee24738219742f072a745e865670df64da7b9a77e2a0f77865b4a0c222b22ed61bdba978c2e394a18b6ae378b206b725d41e7c0479c0e62cee0ed80e43ede604ba5f4fda3a6e9c5336cb6cf070a9bfcc7452b0720825450115f4d790eedc2dc96607ed1186f7fc5d07915bdd007d0cc2f12c5d658c3bbd482a12949a43f36adfd34c4ad21b025d9629deecdd1f70443d39875e1ac22cad070dd89451e9c26dac6eeb448ac69a678baa1fc86658c2518f4c91d36e30cd221e5fef27e6fdc7894d2f317272f688928f2fe1f95c7399a1d31c00f823a79f86de5690a2759f63db20bd1e5ee4778186e232a29e49584f1f21e5c355eff7132251897bf753f2b1c7b32ec7a12a21f8dd8870e92d40d8a494d379a0a5b8e6280cb579e842b7dce52801a34a88936a91223db842c8afea5321637569cfd14f268c32ab0c05ce24b433b0ac82a55603e5d1abea135757060dc60587c4ed01c86a1311451a6d996a4409ac33edb132e0b3115c93fa4f9d1e55715cdc7a604b21f8c269ec8255fedd1e2484339f722406918fd9378153d4b9a5d9d49b870e79a5731656710cc9a7a82d532b3c932b761b170abc88eed0b8190c57ee79fd5e95991fe31d4e803eb1a9239593871a8de7896e3705cdbf60c790e8130af38e2aeac70a082a73aeee7cb2ccac1feaec8f468196d8d8088933b8474bec720b7a7641fca8d5b95427cff75f547b4f16947799fc3124eae0b8423f804ee9edde41fb5836bf6327e8bcca6e362de1e6c643333bc5402b7983935d1cc43cd6cee61e37644b3972528745356e04996655950d0374bd1d6dbdbaee4f4efe21ab06fab5d56e14a0be7dd3d37e7e497506479c8baddda473e7854c31d5dfeabe517ceb3d6d62207e710ee0ba7d2020bb80b5a4a5d492f4ddc61a4ba704f3896d9b31d98333f53cad6df17380abbe46f679cbadf0de0926cb287bdb7444893238948f1df7a4792377d9ba0135926b52847d269f8a4a37b5ddd6729f6916de5ff8a6d6b1ff006943688ca2b13c09bbf6670d4b24cfe6a5b97366809e43a8b6f58469a7bc51fefe203c335bfb2344390d3ad9f54982b358d2078946ede38fc6a52342b79540e54a8fca78c78c22b051cfb312df2caf4f99666e714225e142aee1dc2a43079247ed88476254a1364ba9c09506fcbb2eae42e4a4dca216b5fb94e2caa309ea69a0bf5477d22e39b2f460f6dd5d78146b2f0c145c65e6963db44ee6268a06e60fc1ae94a53c75cc62cfc4aae0971e1000c52e10697314583f658407df903ced2b3ae73f1597af9bc34f2662668803e15d9b3fad8dd058d31ef4651bbdd3a8a70cf78b245a864152286b905aeb88438f917074adac4bde1dc709ec5fa3b0fda6a48a29c543b7256e31919104eef87778f2f5de19914c2d41b258f6c724296e18058ecf276215e6126e808166a473aca3e25da7bdfc5e10e7d60e5be53dce82def30fed12bc6e2a84a7d19d9a2f11bef347c58776e85703e0525d321f46bbc08a675e38cee04fa00cad714503c1cf1d5c9452f8de26dc069673d67a77af4b20610bce1d680c2ec6d9a44d16112f9d67f85d7e507f0346c2c002423f6e958840a0915fd7d79fe86b90d79798776c1713bae68f70f43e9573a65f542aa28116107d65569a7daa8c17d41b1300d1e488a7e894c0f9e9dd9ea5e9bcb36b3e55cff8d2d0a78a5583f4540185e28eb2ebd4f3ae436a1359da0c4d8623331fe6d72229c6052e3210d78dae2142535e8d05c60b67fbb7af8928246370ce12f89e5b5b30abfe576faf863ab9db238a5841dac843f8873d70a06f75ad21f14653ddaa153446b8f5e22be9b89a396c7719405426124d0e9d427ca264ebc7fb67a7ae03741923ac2bbda073a91c6faefec5c8878cc90c190e59b054469d8911d20a83c6fc42455d9b599df1f0a52b347419d2a0cd27e9dd6500063bd8d28e25b1da2394d8f591552e02334bafbcc1b6e93e6c33633113e8c4a27c8facd32b514197a1d710b4db15cd575a4190f6d7ffb5a070100d0dbcafdd6cd0124296ef2f38f8c8dbfd6de640af5fdc2a2020e04656885f4f4fee95189a678c96438f6db6495efb9e25b481e376a15a8dca7a6f73a6366d5f76084cf834aeb738ec72cf4a3dad5f155a497e4fa28ea25faf0214c4deff1d92ec88c883b1f36804c45b9aadb30154c7a1d0eb00706e71257046fadc0445045220a4e0fe168f72119b48dc46c66c0e91670a70c0a9d3581d230db8f7ce1278b6641b794321cb6837a1bbe6c409e82956ede6084bb22228bc5c04f08ff4af850150afb04b6b29ccaea3fd8c22cd7b706bcab6f4ce32ca100bc7961f55b696806ed3a1f2f096047f92631d50fe20d77df822308b49e52ccd8a3a133dd73c55dbf155cea1c89bd63d3c9ec2934f7a0b5d5789c7e813f101708560e5ba494bb89a5db03e30f2be98ac6586083e0e4eb4c686faf4f295f41667607c37a278e75de;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h99bf3a887cea514aed8f99bf20ecdf10aea84c2ca988f924d8b3fe3499a594c4ae722cce2bccc8bfbb4072a690e3ab8b61cfc8f9b92d234e3a4ab1805e1e92e018a8d0587a66b0eb863f8742ff125944ae875f2b582fdda2af10d66ccdaf47a69b11772b18964d5598a1922ea483e87079c1e9562df85d62b53031f62df84865e0c1b838a1ebdae26ca7ff233e78ec2b620c52eaeed8c1ccfb33849eecd92e144b6c6f991e77490d6b0e9a3f7a1c7c7be9bf088114e326c0822b8575d2008d81b0c6c086bf9785c803fb6fe7d3cad2c14a89253c579c68a003c565a8c31409e7e204818ad824e5ca417a9aa5792fb9f00d4a0a5f82fa9dd28ac8fff10a7a408f90ba147b017702cf6e885f50bae9e598c22f8124b682c438b07fb98cc1fa8f11b5f60540126f65bc6f978ae822295e9a0d3eb2881e048f567a60d5b89bde3cf7a07227b438579a7fbc3e5d09b0b2666db3d160558095f392067027d5e51877fa665f9d6ef8af291e2ddbd79381db1f55f8d66658f11d1beec394351261b41ae4ec991e90cc25a1fa84c9af49ad108ca2cb1fd10f284c801dbe393111e3d2f5447775db070f33d04e320e2a7b23419666f40cb5ddb364c9ff3546f91e624792175cc8d9be253d9c9b7d8df25f54e10c189c175e09d248539e6ec81aeca2fd60544318c15cc07ac0a3e3164445e022192a3961570e1454273c96cda63645e71228ea13ee262f3d4a174a5ff130ba17c2bc9678f09961724a2c19baa3d0eb2d27be0783b4a68531bfd82794f415207270c413984d9530c5073da4b1dbae047b8742317afe300d2a5efaa685c0cd2fc93608d030e09ef742aa5afa21401b4a9c2a436e8b4ebe199e820952997e80bda5b346cefc5ef3513ef105754718ddc64f6faf1d9d14ed742f6e17eb56032c36d9c764a6cf1b0f5b0ad55e082c7c157b7c3a9a7d64b46ed69f32c45d810780dda02c165a9a89b1e3680b45f924e6b21ab7a99fc3ea7294ed9ab1a3cbdf82d77f2ea82189a851bec75f1c21414514bf1078e46e456450a65f9d97c9a42ed86f66ecf721af64026bce636f3d631d9f1e6316aa40be230e74b11d7a4796bbf90fdef873167c5c566eeff8ca470eb908facec2db7945b9a595dfae071ca55ab81d5e03209fe2ca60ef05fe0d460794c2034c06d483f7c9a59fc5c1de2b3d7c253c4de77aae41db0d3405f7c5b33a854a2e370918ff0976f41d31d6713a7d08a460adf0085c63750a7ed28acc6ce5048149c138a6adc28559e8e199868578a540cd3365c8db5d86c95cf322c42e83a0399c39805df73b6b79edf1fc61f8d06addfea94c020856192fcd848164b9a641919345107f2eb710c21a4de30bb090f678cfbaf8c1428fa0167bd2d917556a1cea8c5be231424a09128da479b0fcdd2eff87f4f9dc9e8c3c5c18dfa73b643a6bc17de20cdaf5669e16ece09ff95de4779aaaf0d7a7f717ea0a37a8b4848b326bff62adf35f0dcc4d921f8b7aacc404be15f27a4087d2084e67124fe605bf2d000db347749d498d43853a64fc198b256af55c7c87985ca6eb8df75132fc079297f645a0734e8c7096f5a0ee8d72082cf8e36aeef95c83d15fd7d68c76e3bc4b09ddece8e225dd5c13aea73faab17cb84eb6281ec963ae200b84ce1a9f519cb2dc36e4c2bc442ddc1cb3b32859dbf43a4445588c0a7894b4b8d430ae78f551c317d325b715b07c2194ad262cac419de24ac31f88cc7dbc24f017bde2065121fbab9af7c691fe4aac1a1069b0b78acc20d93e5b15b5ce3d38e4b5abc02dcf389137bd20fdc03abd319a26fe0f0fe06125dd996218cc3c31c61c6aafaa21f9bb7cbbc9cd798d51f40c25213c008aa84de52b2b4540a2c5742808bbe81b1c21ca33c717fca3a5cbfb952b57443e0e6f4a770dc5e41a905f1f9d4111f8d23a0a573799b7a0453332839d80c7f4386c39bc17b601afddf7b38a0a80b8f7efae67c19851b9c91601afb999401373bd969a7692dffd0837751e7e3b24531fcbab1d96baaebc0f66df9dc8c3e1658f86c43910bc810cc4b650634b0750fbfc45e78c578740870b1f7dcbce9ca29db62c9abcbfe030e538bd19e5caa13858783161e45a76952dfe44eff089ff9768a3fe8561b7290c7dce01b60e864a640b7293e2bd80a4121ef18fc84dac69430e350dd94f53d4fc30ea78d0c0e0419b18b51c0d8d9bc24aa1b8e123c8284d15de861baf1ad8888fed82b3fc330e31fa734289e29457c0c8ef07e394cca5f3a1d980ca11b07805797768ca8b3502602a2a8a0589b4459534072408bb10617f1c9f3e4826ef7741e77108be725d57cbb0354bb91946f8efb8a54b700a32b1703ead295136f38321383f337b34ddcf01fec0138f5f01c548211000e839fdeb244127059d4a9d7642b792ab64bfd0cf300436aaa26d57f09439223a0b84aae0eba87e273772bb972906702aac2f0e2c494dc84f505ea067b49b83adca7511e5b0038a370e89084b3ce8c450e94688cad5f003af9eb7547c1cdc1026fe8803da74f156dc46429b67537dfb687eb84a5cd252da2e328be3b5811b668c37b956eae5f83b64a38ef768078296e3dfcfe4a586bcb84e9e3c86aab18f96f780a8fe6d43047ef795d3529dc89a3741ebd36d56effa6d073fb5e40c087bfed85acd3312aca6421de743eb0259ed70255fd1eceea6a0aae801f72fd8cd1d28c7462e4fb272ad97bd29db1b30deb8fa04561728cac87a78d371ac11f6296e7b7df747e3655d1e3b04d5a3769e709ef184fd5bc9961ee3074952284372c06626342eff86123d57c566b3ca94e143c629a381c5338ebc0cbdd13e949fed68a899134d798f589a7257640cb48a2595ee3c4b755b863b96a72f9d226a4fd3eca02d9a8d58e91305aa18de92dadd2f478d172384815ff484aab4c451cd11029f898db14e09d9d55405799c2c342013068c55547f9e4d45540be47e70c5c67c62daf1aa1d087fbfd1333960ee46b80b6812fb0a6e5efda5d6d6f1dc122870094bb55b0ff0283c1d28f2b176a6e3ab6a822403dec69f8566f85b7e8e5a56fe8f49f0fdefe7f412db1f479e5995be5ea1bacd6731131c244c3261744e02432a91481fa5085a607a48b10265360f58f022e69e48904ecdbf0f0be3c7568f7a6fda7f4580b63816a5769503c2bed66e74f0ed15f5f95fe6e293898b940338880219751cd703dc349bff7772341a9323cd6a1005f93dabbc9d464773404f06903dc404f2e7723430718424c0f09f4e685a3eaae4b2868166f2ce667576b818d04651037d3a68b81bea700170529d13464944b8cf746f56fdd1e5855b47b2d3e96d5f5da83239cd20005a461a4f5322abfce11af2c01735c9ffec3d9c067439c04c9b36984e3c3416d63ea8ecbacca9270afe24147f87aa8cfba849f22264ab0db2dd7961827a86360cbd3cd8c5912a1abcfc040eb1fd30e510b48410fadcfeb1dd32f1904b357bc4b50043b940a5b7ace1d9003ab0c72d56f8f37056b5a83a7a9777c582e40d4bc2a1a83405e41a2d4485a4a5436eeedef4ce1eec94e155ce0503bfe0024713ee338f8d83ae30f6c3bb0ba21760da39b83cd0dc10959a12a5dedfd0830182ea93deddebd94d60918c9703f8b5970b73778a8b824fa845349ee8a52ef650a785843f8a107205f4ddbdf355eb18f14b418039393c4df91142faac2638fcd435fff332c158b110647c47cd4f394b1d984e0621062a5dcfb00df34d7f505c106ffaccca98a029824cc3923cd0e8c992717ac3fd360b7a478734a9e2c87c874228ded61b4b80babc526f8d957f40161c3fa04e5dd8191d03ecc4b7a6860de27c8b60815acda82263498e91b189cbc4bcf10539ffa8bcb5ef0c77e0c3cd89fd77a1884dd911764b5437fbd5053841475c21a7ca0872cbd504c798f6884440225b43da4656dd42b4c4c7504b2f2c5c1ebeffdd586c34663144c779482ce0b5f5c5f76ba4be2ae0b93633886b328f80314b886ba3b886631a230fb90064ca5abcc5ec016bbbcfaf2c7171d39469d3a586f327a150780fdfe87df26e52346ab55978c8f49bfea997320aa7a6e1d8cae6f0013c980278e0b2aedaa352a603b4e1998ec10e191bc0d84d0abf1370430de92c305869c83e2d975120710b65c7b27d1ab3e17c777780b3dc226ae36aefdc7167645e87817db5ca7f898853134773b1c51e81946856594e500d08c4705ef7c2cc4d356caf88452f8d9564628477bd22f93f61935c4918103e283d962273ca2abc2da822dca58e4b2747e7cc4f17f2fb37ec61d9f6ecb09a4d1d01adae2f532439f3317a972a2e1d2c0a9935f83b4caad78aeb324c43e3c717f5bfe2a221234730cb55e21c7d2ecd7eb756b48d0f00db2be87d2864f8ddd091c67d681a89ba9ff111b1712f2a1f6fa65560cb5957cf14100db943ca6691b7f221e38497e0c1a81e3a48ff43322e6764f4de024c4d1ddb82d717fc6e07b00d3c2424b78aca47be79fc3e7bb95948ebb9b293919ca810a50d2ad2d0d26f1695cf76e144f3ddd6eacff31b7b88c8fa043c3dde9047001172c618d11648ab2751072464494a8698876fe12314f048b391fc5de7112e133b38e0f2a8dfc6110ef9f2681bd08a6fec7cee417542eb93bfdce29c4c6d94d737549214ba9ab9b64f5b51bf3bc42d5bf797e7daf22166b1a114b65b2f6ddd34f517d45e44d684f711286eaeb2250f64cf6d5cf1c1848c3665f86da3c408eb0ec60f41057fef635da97220400728e5fddb991efcde5c935022e3de7e18d059856b0d154dc46960905ad316bd1f8fa1485b260016ae0793b7979ff33e52a5e770ac31344114b90f1ac996ed97d1a99ccb942281194e590caca020af5334188ac834757d5f23dfae1c40ed83516e2486d6bf80f7582123943f54f9d47cf3b117b57acd6bf91a2557a611d079a089ad72fc587e4bb9c6aebfed2435d19f2051b3e5b03abb50a96c5895113e79be5993073a148956e443e39c977cd7e1723f04f6583418c87eb0a89674420507f97728630b5c9b95d7d0ab8a5f5bcfb2b76547c916cc965813bf0925f973d520442d4f3c61fe97a7ad0270223dd00a831320a2eb0a651290e918e854017b427b7de173db3a92661e5cef895bc9e6e8c39e70de0b405c3f8db9d337d8b34b43708b5140e55d49c3ed5b6cc8f78eab5442a1a676e73c92d44ac0a35a74e4c006b1caf74e6e03b8090cdfec23dae356ffe445fd56729ca653a44f806e7ff30b0d716f5a64458f05fef7dd9b3edc51fb2bc8b77df9bbdd4b7a22348bec3da6d9a7f7d66b950d994c09be8b46b6c686c35b1d3ef13989a1c4af66672914269e8e006acd5cdaf70d59ebc688c12ae4d0aec4417086c58f60fa776be5a4aaabae5d6b9336bece0828351c1d4028263ae0220b104a9566f7e7882670ad8e643a9f60ee321309d422b4db076a2025e4100209a7b10a99fd197441141b1cabb392b03357f1eda300b93e7c8a37e6f18bd6ebe3049a696c907f4c29b3efb85d63fede23cca395ae89cca6b98ec497101e5d2f840b881ee0fca5e2450961f707bade52dfddd42d6b1322703d9f91dc7b6f1b58cd3029829504b2217a3ae14097245596856573908862246b6d25911124684046ac9900ea8051c738f897f85443666148be5a4e84c5bd8a428da544941e250b4e3065e50da66f17cf0d6cc5c92cb35110ed15a2ec1d529071218a3e963ebc583a11598eebc51c7984bc516959d117b522b082a72eabc45a4591120e466dba58928d7e62ca965b27586a56799183986a70680a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha7ab8b09012cf13c360fd13d4bb16fdca810b70655d4d2661f28101ce4f0631945903b5e81e32fe731801ce2b2a7cddd7f19cf8a98c1b08260566d72c517d8293932b6ab7bd7426e92198b9ccc5c458dd366ca33fc6bc8d01adee95ce5c1b2b8d8dbbb0c5ee6a1599b76264ac706bf954152cc9a6271eb09d8dbbb12acb1aa02f10ed763d5631fd84cc737dab9fdbcd1bf86694ef474734e628a388b99b868be577242776e7db391bab93e46c0a20ba601f10708d0475c6c627b541d28b8ab3c10f47d3900281e2925010d2407ed10cd606968b77d702ac2307fc0345bf27e720a491c4f5ac2bd080f196eafb763c1d33cbf8418ed82be4c6ae18a91e99d6af7bc59533e007ef35a0d4b7899d9716011af5e07033a2a5052b99285d8e5936c85cb898ee7491adea176cc6ed87197a8076eee0dfcd07ef96bf07b4ac42439eb8ccf6e4e03746f4c25a14893707f13d183aa3ab967b019953a2a64bfaf2e8aedf60dfc63e72e2633051b15338863b83eaafaeae7d5f05464e607502a7ce074c4669a1111df178a3c384baddd3fab569a539baecd6772845300779c8e99ecdfd407c5ecf90acb518c20d6cd28e303ae0c960abd2e7135b79495b775703ca899de133aabb8ef891ecb1fdc86e564e72297a7778ea20026e02a996574cf694fb6ef7e3211cdb60a603299ed882d34583e9354c16b93f45830fd2c6c9003d263f337770fc9a1eb5a4e40c09432996f31decb846b692beead049eb1ed92661ec5f7825351b4c31668a366ee4be16ea54d214761ba4990a826cb0d3f7ee7628efcb17ff0445f14420fbe826d2fb23288165a45658ef101653f80252657eb3e98a96a2088181bf29dd8f865b694e683f07ec923cc7de74b1fe45066bf164478b6a33b4c8f9580241675470d5e12151490825b8ff2cf0d60eb2c432b91b81453c0bc832c9102eb44827fc987d55665453048d4a23b897b9984cbf63eb6a733bbea7505fa11faeace3fda1a50fc26d7f776bf23cd9ba915ae367423c6cee5f914c042040fd9f84131b986304a2310e32d82f2f80bbcd1ef79d8545ab9462f0147918d80f6b922fa96517aae22aa28b754be5676be4f8102809d42b97b852ffa64a0997a1ffe332c0ffd06394ba0669c8990941ee7a86e02e3b764e7755a174bea43457ed4a6dc5d18d648ccd1a13d745b53c1475ddcfe125e105492309d749a81c347018102c06eaa1af1c2e9ed8c4c5f573276c828f2c777b50a6b3260f5eb6974501774af0630f842c0622a729b1080ec7f6eb458760836ed48399409bdb405efe3734ead69674a370f19ac1fc09158dfacf616d3a3a7125f0af3e59e154587f8f5a0abb34e46b2fa248d4883f0cf150484ab8cbc5802a8adf0b3d39564c064c2bba9f8f2a49a7d1266cfd8509f53dffc89ba23abeae8cc83c6954376c19f953200b52f7b2b0b1318e7fe2799b7de25bb1d65a0af996e45acba30a1f4d5126135a3de85e0422a1289d3ed1959eec46faa6d71ac513e0d0bfe91bb952d49da73a25d688242bf751814344e989675a8f869683c57d2616137a0528b6ddc199b72cd46935dd07ec52c34e4780e11c123352ffef774c3d3513385302d356d735109a69dfe2c806a90ddcca229d1d3236c43e30faf398d46ea4510efc45cd18f0db56bd319c765a8c37d401fc89a5993822edf9d6ab9d488e2cfb177976b9c9b8b85a4e7a4a658da42c4c4d1a6970234c615b704c18cde8b58872a13c6d22ca29712ad7c81f234172a747f41936311170a21f2af52668ff12bd2379873287a84c0e6f824871f0ecce75caf0f78837dbe9b4d6985ad18939870d9422ee4edd721c15d20a39ddd71e7304ef248d0855e5941850009f11e531e5b456ba1625966eba7234182ccbe785a7f2ae6728e0ab45e1cb870fd82cf678df28297840ad6ea6293ee946b6fe6646ce8a0247590dcfffe4763e2d28f8c74b64ccf808f26ff13b893e92451a4d4fd8e0a5d25c92fe12310546f3580afe8345cd80644a8597be7f500378250eaf9f57767518131be2206815d26dc65c77f55d204d5143979474e61626bfc5cbece13996b4d834fc589d14142bedfa7fedd6ce7cfcf009d764f3de39ece3081f22abac036bba74afa3b18ee5de4e9879d1fa2ff984ca4daf6b52f1f0ac2aadf45cc428ca25cce45897ec2788e5af2264b145b000622aaa869f4c468ee04f23a4c4aa0cbeeb0a6efdfb9626fdea6b335b9f3fe584582dedd386ae9d941d5fbf112ef195b8d536f863b5bd07e7ea6fa21f8ef68f0fa9123ee26fb0f6a71d2d6ad32ee47df8c9c09aa3dcc2b80ddeb4ba9c8b739b6eea6f1683667f9281e039787b1b87f1537bd21415b2002c13213e54a915eddfb60fd926b2e04704b6d9accf39893b8a379413a157db1e78807d4203438b2a992a9b4859e35f2cb851b02bb9a230b715a84389ed910bba91bdb032cb8478dcbf029ced0feb97d1ad5e740dada13da1f06603232d0c32c00f3c5e2dc9349086338e596bc9f98c6e628979f2ef3d103324b2bded5832de82e332cc28ac02a7e0f610e960177de72fca50421d8ed0c7fd262c674de3b9c28a52137f57a0913c7a76a32e6be8c8098e3ffd2bebeff18bba9d690b3e3217fb6c6e51d3e4ad39097822660ef2dd637d3535589ffc3351c70511aabbc87ea62f4f54b946490707931450277cd6d8f11a748b107e60e4d96d70aac73e165108e91b0552de0504daa93ccad640b5c6244d113bfb05c2b257d854f8100be361c29821fb06c99eacf968d9f1398cd923cf6433ecd9b1a2dd9a7f4d0d43c2f925e931f8d867a13256af934d42a5bb50ccc54de2e5aecf0ca667444221cf7add1c72ac7cb2a02b8008c216997df3803fe207a9dea725e6c3155f09098047bf7d36e0fc26490fab3ee7768b5aa8405be8e3e717d28e8f96cfa3399978c534e68c11f50f07c973ef1f768147b1782208bd7912953988b0692ce5b4304677d9aebc9fc23f2a3e6ec5b8410cc4fdcd0d7834341834008f22af7c17184ba0aa2f06d3420b575fe06d3d7b90c3985f148a531dc15a1a4bc2d02f1b0f48cb56cf067fbaffe1e163898b156db1c1c46064a424641c40cee31af1921718bdce91f2b584afc627db4f635d8c4f61093eda07733157b6a13389ad1168575da073ded041257752420553c1482978c332a9f3c2c63f5e7f552abb64f62b79aec8a0f7dbffe1237e6cbca5e14d823c751dd5436298553ff285bfa2f4ca4846900064475a659761337e7e863a47448d76b9170d4393eaf403e8d59d47b96655b3f8abd66fa857e254fa2d9738c18f2fba0be7dd9cd2b255508d0b12663351d8d8ffbe175276082f3ca0c249e11766926a45e7f87ce320b65c3e50faf5739e399be165e75ac3a2ce36271a08140bd0979a50c6c2c825df856b8f52fabb2fd776d331f8a9df08d60868726486672c007b7d6ecf6d32d182e1f8112435f489ab60e1de6cde2cc21bb8af42397556d6494f5a17284253e09885f68e696315852738a18ca74f27e45b3206ef0974fbafb5048f065197e88fff5c556ddee28101bd8282c3f97351830c5df2dd34434458fec4b9ff4b9523ae6380b93b76df108883a062011b0f54189e68fcc31f259f934401cb3fc8f9af93ae020551a4156a7442e11aefe2ad36690c1162851cd8fc082e7a3dcf3480cf71b2258e8fe3d293e7a1cc894906e8872c87d5c6f1d5f607555cbebd66a3978eea8f30ac00420967736635b9e8227ff6507b2267deb77ad2d09866480880f68aa7025f4b6299d86f04346a069682ae85a2c2ebcf02edcbe1814d43f79fb5d5e4117e460b398993c105ab64576ea957d94df15e581a203f7768916500128aac90cc3a42abf47eea34a59ee54c041959f8ad3066a75732c9988cea1ea00094d6d60cea3e21542fa7e10df0298a5df04722a3941418a57592340db7decdfc7d69c86fb1cedf66fa7f9908fd02b299abb1988190982c651f2f8e644791c3279eb7749eb8ae9993969c8f3f6bba7eeaa232ca39ff405f562e08f866a0991972898d82882856bf7588352eccbb6db9eee19fdfd56514e06ece8cf59090f6f4c9b56803a6107b570dc049e53afef380cd6921b561a0787e7748b01e13121746b13efeefdd216e44ff4769017ef136cae14e580081aa060950724085dac7cd598399b246168f0371602015fa074eace7b6bef82650baf6627f677f60f333f69a7f0d58897546ec8ab6127e4eb23fb8d3d09ba5d4bf83d3d3ee1469c4b79393deb6a9bbe614c2010edba4ec911e14e32b2bef683852eab7f1d7fc757713e5a55eb6f9545f934b06423f355d21fb66b583d612e552ba17619db88946b5ded5bb252e8df84db111c1c7962db517b271d10d4a419070d09eb44fddaae4157a5f544e1a1168211088d5931082a4cd0bd861cf9bb5f0331b2c9a55573c3cac06019519a0893350290fe8e90a38a8837a862923a6eb0d88de7b13b94b035309e1dc25f5e20c5860c64d3976c8ad0c169d5740ca5e215df125371db4616ac8ee448f4202f02f1b168c5b1fbb6c7a185bc40c44bf9e69a2f4d5db31c67f0fbe1c44dbda5905edf64bf355c27a840539b8b11bea5a8851d8cd877038b266ea1cbb9714bc56ae2063f600e561c054d549f29c8f7e2bc6a24aafdb10a6eb88655c38e69b3bf38fe0c31558ac95bb72df2205b3e561b2d08ebe644b63bbdf380ab159ce95e75269998397e72a03be9800158e8f5af71d96bebbb9116a67515bd7f66c7dc288b551a3e43b425b5c3d4f004f9e0cd0e64957862dbfe813f71121f35c1b54c1274fd721aa0d424ea4b6ab3a0bead7c1cc0fc867ea9f088f075a97fb42fd46decd28870653cd166171274f7364ed779c472ddc7d97868d8a68ee3dead36c1656e247744c2b486741a3404fb7d00a520e30055380c9004f68a9adcf06ef599653b4d71694964ac5493d35840b51d5f0a09cad20f7e7bea82a566422b5997107f1dfc5626ca544d6e3b47a9c08bab58d1a6eb4bc19302ec2a43b512682caad4834bac0db62df66996f4ca0b99cb0f15d369b3328a1ce47463b135dbe41e89abcdd5abd0c813bceb1c6c71f7caf1348cb04d56de51bc329ff9f99350964510ce99ff842e833f4bcb37861a98cecd0a698389bf9f88e1d2233e176363f180f7af7d3309a5b376ececa15c5fa59aebe7040336a417880ba769a487009a49d75ba6cb16a3139ea38858fea201c35fe71ef5ab4c7626e3414fd38de6ca8a333ac2e6f5f665708d6b1e144a91abad699cffa248c7a0845d8502ec2c1a8a66a491f3b50b69142d68f5bf38694dbab6bc61d39cf3511e2ff726c03923d42d667078750296adbad87eedf2afba4475dd721f3d9c4b2eacbbbaca8960f81d167d2c54455135d573229fe917015a85c8d0a144036fad83367001481ed6106f478e2cc020b714444f18f59dd47fa9abaa4ae8c183c586ac6f08852f9f43aba16127e4787e3a4721ac85338e823486b30d7161a0fe6a3861a051474dedb2c02b7eab14836b67935f272fd7be98f9df8e0fbf89765026c243d4d9fcaf23e9ff5b80a41438240f73c607b577127274ed22ccfa83afc16827b187abd29966a6a4462890243da8ae798d84d1d2da616a87af294b6326de7f29cb7866a1c5a3e5ed3834f3ee0ab9c166e8f60c8092822061057613bf1e61b42b7c226db7e8f0d4aed9d91ce5e13fcae443689516a636d2c8c08b6c58812d2378e772ff5c431e0f532257341c279f657e465065b55e737099ec0aea5abc269329541dd62e9fdc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6a5afb25ef464641509a43277f0905ee41a4a33da1cf1b509653915642e70dac1fa065152d44c578a907473987b33ad527d7d01d0e7f0f755e4a19d633fe14dd5e62d825cf79eaaf0f380cac18a3ec07d903a8ede16975c5d22599462cbfe637835baf6bb881e4788487e07f5185a6d5e6ad1afd76fc1788f2603e4147e61f5dfb54350e1469ceec6bba53d1e298a18a6461f5f548154673fd630d725fc6209eae9a3dacc3de4086c74ce8ed3445c59e64253c0f956550b740527859a957043a0e2d523c7e937894d4d6d3391f7f33599f10f60a20c6536af99a9f328b4e6cf83595be4e1cb8fe6e7c7dea1a869c4135ff01128a727ee533a9f3204264c4dadea928820e4f3a0dd03900a10b8fe3dc3deec8135c3eacee8555683ad9e2f6a1b8e9b3bccf2f9318e9997e717f5d894d9b4076ae780a9cd2d1a2cf1f15a7505493a67573dc49fcb991cd4e745b6a9e59058417a60e75a8e4d832030738fb09435ee63197966b9e5bc377f4fa5cd663283980eae6d5de0bfd216e1cda165d527d9d06ac100e7ddd2df48bbb9f22998395276e4b7cf653f7d7ab8cc2cea5ac10767698e6fe5a7ba38e01b7bea949924a8ec5b1d9778799ee5a68200919e4de56bfec5fae47d501ee29a9b6dc5aa4ee1f2640ad3ce774704ab3bc2d40dbe5510fce98a0ee86963e830d449c07b421c357ddd7e5d5ca56720db05b5062d65d11265f235235bd73a833fa96208dd75dd7e8f3ab4505bc06f061624c72f21fee10f8d91c84b7285e16883ee6c247a24afe006745bd90a2dd2048c562741115d4e43ad637f8f4a72cb0b3fcacec006604ef6c5de0a8edd795f63b642402e40468b0c45cc205ba92bfdcd1fa20a74a53ea644f1201a4b200f597ca9b6b1867c67b57f5891ba98d8107bb71b63b58aa95b932e8b43e63c65553008408bdcaa1f57bf7ce35423e877a257b33cfc1684a6a154e5433bc941dbecd890f11dbb48f62277cc559a24dc52de19b56e3f8f13df759b6ee767f5c6b8b7f756d64db23b17f14842e0a589c4585fc994d652e81ff46391f5bafb28ef73557b2ae02f2abd4b079dfc7e9139e6936d1ccbbeac76b6fe0491e522dc74a8574ec32df9a6c5a7ad58577591dce17004c0fa65b21223e9cf802fd7a03dafb8ef26e0276b5f1c9ba2ea852680d095ba92bccdae0ed0fae504526ce88701f445a22e776d8fa39ef4874bb7cf4fe51b33386615e741bd20386c41cf1f4f9f8bd2c4066104710e01fd92d5b51634696bc3846997d59950eb6fb08863fc5750461eabcbf6e94b20fb166cf60610d5a9e468b33d1a1d8f62b6a89498d035571e9d1b7f2e2b5bf0292cf58da007276e6bbc5f5d7f26089146ab7e44c86d8f317db2df70bc1eb69e4be05b9cd1b2c0981085737553b6b847f525bb51fc3b37f0149c010ee21205575796b15296682069d5689fc089a938ad5813c2b9675b4d8d7de9b9f6a5a6cda27e8d27a216ade54008cee81b907956f8bbb4ce3c7482127ce77af578a0deebc0c35e7f89fb28f1e52993af10cdd17210db78334dc349a11df4b8f72676a855cefe53b1f1d7517af45fa691d7721335f462479d5f83c0f8cb08ac50dc3b17135370c857f5e98d5d871b109c22790d6a36a02797251c92bc2574f1612134ffb0211ba76a9156922868d071c1d510a891fc7ea66604aad0b7d620359d22f04bc9bc33b31b343a552150558bf31b1a52ca211ff7a3def93cb4910116cbd96465e81935be4ad087d79140814c4c99bf5db937d5f4a28202af762290738bacb93c6db524e67152dd8b2a8136bcdc8b744fb884cefdc82fadc77c2b90d4333a5f52a2aef6c595a0834f109c7fe70ecf55bcb908b4221f256318cefe17a1ebccd3d02bc8b169fde7e2737a3babc560037e338d1d552d26ff75dbd8d163ae0fe096e649ed84b1c773d81193385b52ec8974e982f56d254247138dce09739104bf264f3df8233dcf75529a15304542e34381ed43e1e83535876a5f088dd9bc734e3db45e191a359b68c9520882cacdc1a02d406a3d66fae2c8755a76708c6278b595c02b68d1267116222b51c35f970ec54047056e838ae5fe1ada4a389140dffdb499e8920f1af3ba21e71559e96380c1c68bcd60e8eecfbd7f3ef6cb65b99006df3d07e7b4bbad8b26d4f785b3a81453872594dbc17129244cb585b07b15729a244c00f112a28debe957334b755265629d8413996e70f8a890c524b89e759bdccbaceb1c30f85b488fc94aa7c7822d1e3ca91db57a5a24a4c0e54e2637e76b2b87055fd81e27e5540d7ccbfba396a4a3cad1ca680eb2cdbcb7bf821b42f53c10c5e7fc02bc3d6bb0f1675d58f0ba2286136cdd3b8d8e3ca407149d921849cadedab96a8eb1cb42df552dbe94f23c4d14110ff1fcc4fc4df854deb1d4e125ccdf58467c45b04987e45e13ed0c4d432adc450248c7c9637f116307961236f5a2fd91f70d715a38a48165e2d7f53f86f2406640578f6a9e2e51f9240c0f21ab649034c11bdde3766b79a31d9df1428677ec7e0b8918cc5fd48b61f2eb47dabc2468a34ff048af797a8de2e6f70e8abb51cecc14ee423af67efb87c4f1f9d276df9457c911c67e01e2d1e333c3c8b86bab5dc6930a098ee2e6860408404ee113220d653e2286c05d9e00fa03b7c6cc06556a5e8dd4ea14f7dd94b574f2f1994548344c3dd57bb6b454cbcc4e56174982bc8fd2ad13e04bfb03cb0ac0fc8f6cf5a3e5407ae4c8ed0ef5afbd04874bd336d330142cf1dbad4e79fd29381f5e25185f12de24942a506d8ca0f4b6ea4b349757737e261608a93cbb9132d69c6acf0f1c1b8dee2da0e026375eab7afdb16b3b155a3b27d4968abe949c1708c63dbc7bd8cc484ddfa3e06c55605c5002725432580a2d59c98119122677c7913d366c59dce7c92d18d21318a1e4b3777980b099dcb89e659734c0a43c645696bdfaa17fdd611c247911ccbdb8f736c0b917aee47a07a00018f82eb09a74f0f856725c98a777c353594ca60ad90757f61810e1696e848d364e1feeb1fe126a44d61362ffc95d94b5a22816b182dd12bcea1b2a3a2e339f174048ba488fcf5808412b5e2015a1e1c2a2bcdb5aa937898085440646947ac9b0a4672d7e0f730fcc2e4aa7c803b80e55f7323305a77ec815f384a975f7963b0b8691a82bca38ae75dc2021a83e9f89a7f9e5ee5d521759473d3f24c2c62cfd04c1a8d52a5707826ad57b7c2b3c91a82dffc0bd3acfee38c9fd64fd4edf94118a58d69a6799d0b4b8114c345081776b17f20eb4f08281fc2b05f4d4d585da1a8399c4d5b491cdf93ca533608b7731fa9890363dadc50f2df5d4abbef3c5a32d72a3b825d833167cf074156c6ee322578e35af8e3b33e30d3064418b1d7f95218627732394daa1d05e8649c79e9a41b5873319c0e1233d80cd1bd13a7aa531db0242f34baaf4b07cfc79f7ba14fe71c2ace35f3bbb2d1b07dfc5417a834f9672063626aec20208b0bb9666098b3e12d795f14d6fefa19f01811da13e9cfd950dd6fb7cd3acd3f50e47248951272d86e16e15f957a5b86b0952c7a6d1db5a49e2533a088e201398e11613c955251424289fcca33ab5e3f5fa7a3eecdddd726ac40f006ff9fbbe95b5d73c2163f2674face540ffd7ae5c4a00e07508d102aeadbc1f6c377559414d7b97c6440081f7294f99a5c18f041f607d8680c2876f077f98b9c83ce708d6a81f9af6b6cb3d1bdc8cd0953f14160f54503803bb066ea78d3df97723b87279c97e0ed6ecbebc082d4bf8633b0fb2c953c888ab2694f0b17a4dae4ddb1584ae46cd185b159d2c0a986c21f29f305e9f26babdec716267328b9ae8632be1778b59215525ece8d4561e1c0ace41090b0774e681e7f9769bcd06f1f6685a842e954b54a1af5142dbdd5e2b2ba56f35ba19aef94807717e38199ee8f3067c3e2e8c743424108942183374461d52e9e2858e6b69c89ad32fde07476922bea9d8e67e16f824019683333f538859ab225aaefbdfe8435f05ae5882651a985c7f0c302c0eb4979fbc62288e5cd00fd45c0694955ed3fd4f5070cba979bd1f5cbc4354cf08b65627a9abc68a31f575d720cbb50fdcad33c10194038a0415f8529c7e60e3c8413a2f6b3652598c5077f0669d2944beafea8e41b76d7b207ea557f8220a56abcec02085d872e663f3dc5147a8e5c7d80cb12b3d266a4e7529cb98495a99af0498352db09714ce9e6acaab2d32df4f7b59d855f114bb9e5c072d2ebc962a624b95aea9760b69c9472a8d3778cf723841398c19c083eac38067b1eb659657a80fb676468d307c464939433c0ef98fadb9422e3f580b4132dc435196702e420f2df784dc804293feed979574e35860a82634e0d9f8dd681650e96d050364d02e7662b3778762569928e82a726df859bb0f5ed705f2a91b4589a4557c289169d6a1d16028ff6d7c1e353c91e2eff7f35b0b1c17169bc390f10cc7404b7a06553cdbf02ecc44512a6ff7a73d90e1c6c7b57b2d8f25c7fbadf688738f40a8995d960bdd57e89a5572c33ec6162e6a1de7bc5d24c89a6b97c8ccac7152b493caae18dc55abe41b6398f0fee1ad31e36871dafaaa9ad6b343b76a0d27ac45d1acd62c1f62570dcb39ec1e78606dc8f2697f28c55f5400070341428311fa032713edb52f2a1a4d32cfd7fe794c433794eaa01bcdfd1250098e37deff72ebadda3ec5b936a94586892b6829bf6e2234fe36ed6b57aa2e993cb79572d227b99e23a32efb94dcf6fa0f38d202d57976a3a2184ce8587a7b5dc03d4e925412127e123e4151bb624ce622e7d33cb97b9ac6c45d78ebbbf9b307825aaf02a842600d1ca37f4806ca9f304ba4cc09d3355c3c4da50ec21e0f08feb08d7b5d593d2d51bcdb5f6f8b6c025138c90139298d7ea32675efe3b28d89e5bf8d7eb8d61d1afd131d4ad00c95151735217fc2b9ae316c4d017cc4401785c617029a42046cd3da64f90ca3aad528f9294d14001ee32a2197248865f704d51d1fdf026b454c3a120cc040b9a5c7b24ea234a40f5e864bec6453e1675de35f3acd6b9cbb2195d03115d5ed80800c95f57f42083d2735ec9e152fd84888757fe824e40bc977d0d83eb4f98bdca3a93701d0bf6467be0769269a569193ba61335b6d3cf7a40dd06e3cbad6f1eb5872141a35333079de83be7248d62f9cfa40f4f7db784c5ddbd43550fd064621281a32e98f352f7b3430628ad51a928ae885d4e215ffba1d73898640d8f229a7d643c4b50dc78d4a1748d34eac22330a58820d5f2f98e4c1e7a3f4904f8d4da11ca7a2c7030f17a27a9f8e5e8a719d520fca749e4e358bab556b1e3670dcd0307ac4301f7a6ed99c6a8a82efb94e55f11083ef41798dd6a9ae1bd78b2eaef538cbd593ec36b26813d8ce1c6f1c03f85697cfecf8bb762d53231c1ba44880a691f8b5e97d3f3265d5bdf8ce754db56c205960649b0f9ba5ba3d1a943db5a5e89a9221d4f1a9f7bd1ec7c2c52e363880b473b1b4793a3c2afadce8822b5d5c40f026931d51c78cc87ab4c311445761870b0f78bbeac07b682c75954cf3ba9c7131b1d6e8bc23a64c01049ebcaa565427d25fa20bc35db4c3425813af8c4a12f9e5f7f561f3597e1b810de6e9cf911d6ba00fccbd38cb4e661fa93eb522e4795c5be93eef3777cb967cdfa0091266f8e4169c3bbf7c31b2924f351125424af297af80d71066d8c7c803e05e07ad862898d610afcf018699fe5a91f3aab5b8feec18d9fa632c5dc255addb926ea87e53ea031476ce1bb6400;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'had7b0b00e3f4b894ce8d2da83351fccc7da11ebffb9698ede6f03acfee7b00bb01ba4ff6a775021159199ebabb056d9dac3a917eb9acae96f569d2231800e23bca2705a09eedf0ef7d949470eb13bd26a97086f058608485d7341b83bbf3b3986f6fc8817d1d62881af2f576cc7071347d12990961350c0acd8778039413ab420af95d86a96dfc250881fd37edbdc344bd17a220e520247d497e5f9793b6b1cef2219fb8e9947c5b9d34e467d3ad2da9368cbd4f36d4f722f69ffc4d5c46bf0075b0e9a122d1237f7c0510b8e775f9a9ed864e1832bfe82e54153a940321e0a6f94848e39f86639e9efe4484f19efc2ac54c3a6ffccade729897fbf4a6184537536d4cbd9ce2201e87bd65748b017db7b2e0611cfbc7385eb0989dd70c2b4aaaaea4407e72355d7aed6e2d3adbb6660eb0298cb65a0cbe88a5553da42fb4b1f0c3662c847e2cc92043e1d8818389e09482500214abf77fb3f83a44d005ca64f85217ce69f4d20d95789bac3b1621a67ce6f438d4254f5086bb5065f725b69a24a41e6ee60fa4c4326e559056d796f28efdb0f70d16c5aeda7783a00865f0231150cc63539dd7020c05aa54c149f15495e8e5bc4f69945d4ef93ef64193725ae8e87af2b66b7d1e470df9bdd156f058ce12903049afa2477810c4004983d8c7e9b6eff467479677c257dacc5a3d66f3c110f10f9d863b050e76062a2229a36f7900ebd8eab4b7f293120b434ca3574932398c1ca833ddbb442c6a4fa2d7b59389ada7f044a89b2a14d5293df608e0aac1c4ce88084c5e852df1e75cb9bc18b9fa9b6fba2f12ff952081a175b592362f6a18645605829195b4d07018f1b0d1a1174ff0f3b0e60ab16d73e5bbbbf79058a1d84ee6ab1a3ce981bcc4b3b5640e526cd8201ceca9beee82fe7481dd694d72c039f68459065c73a892c53a72d60001d12e4d43aaf0299d923e784cf67c838e27ce8fe090d53f77b960329bf9b316e1f03ee692492edd5f31f06e3e2b9e6894b7cca5449c2050724b6a4f58edbc68ea8ff7261dd27722a777aaa90fc7d383341ed4cf2786f7559ecacb66c7f4bd7717270f1c992950f4ed7cfaaf001cccad5a08856d9aaf246a7ba26ef0857e755d5e29481b36c9f7eebe2bdf9356f115dfefcc9b93a77b133faa42ac0db7c63d22dd15c2c104c77e4b15dab6e5831b9ada78c3825dbcaeb403a07dae334e51d65845b7ff790717806f411c0624c5f682e3ed0f059791f9fa4ec91ce1f06a9adc79a1ad33743e0becd5f64ba1089c92ab276fdf8ae44f772d2ea16d052f8cc9314b611ebc3f7589c7b12e9129cf0be77c337ed5738e3d7dede7fee703d2dd2f84636a6b847c8540d2ae5a22047b7f4c791185ba81272a761e07a14905635112ef9aa4f5168a4fff6968a37ac884448f23558795e7eacba34610ef68ef41f71c61ff061610ef0a1f411043b9888ad5cfb3ec69fee8bdc6d6bd560a905602566233ef08db4aaf80c9adeebf36a2e6febecad5b262febbf3d9f8bd4d49ba08c9938de2970ef1a7d6131a569e34168d2d445e68debc84d4e3892796c9e08ffccac0b066b83fc951d8f96ff70420db10f234435622617297069c402d0f45ec40aeaa0ea27d80a042a356e6698eda0cee56f60c963c10f0c11380f7954dbedbdaacd5c07fc72ffe64a4e79cbc8781df23622ece4453c8711e62ada5dd59a3a8dd0eeaaa92b36421416d524d016c07b0ec1476f9d2fae5a687e67dd015bd19dec0a7d0fe7553ede876508495c307934d65829606bbb9cd78a64cf7142966fa1c1db6fb4db4200578d196dddcfc476604f26262a0840b8878a194eec2694e052cab5692c6e8f6c5686541440f40c56cbec073ee421487d5d8d933c9df4db7c53194515fe8a33cfdb6ed18cbb053f8bc76341789b4b13c1636ff23f48cafdad2f6363dfe58997e0baf7a8a7882317b0da808cdcfd8dac5922deb1eea1437e9552b0f180836d60943f6198b2021ec60816070cf3b5405de7d8b139f243be9c59d82dc1c5cdcee8c0a84003380a32c2218c8bb2cfefa590a42641678a7b8352840c642314abb30e01e5e1011164f8715d8981f72a21518a8394d2c0643ead87b3d669a071c9e908ebd6dd2c7432d0c7b1723ed3723326c1dc82924e7f15a52409c9d19850cace50938ad3abf7766df9a3a368c51035846ee1134014456e7e3be89cd2a9242cdfe2ac5db7ce932bc7d2ba1b1ac2dfd359f95eeaa6735ec7b23cecd6645fd24712e3fbd6785d0b5ee0fa42be33449366a8ac6da909dc3c4d24a85c1113c193c532a5e1ed609dc513ca79846830f5ee5d610804594525c1a2d87d60eafac2d1af637c139bc5155fd5715fbc36d4cc05e8be2be812f0f493462aa1584e15449212bbc260c0d64c6f8f85f317d5c2fb9ef43e2feb82b60462d9afc441f9efe6885a6ae02035fe5a064a13929a5813bb5417c71ffb786eee8fb0d402db566ed056d2de23ba622717563b145a7d7acbbe8d85770cb595a2c958433fc91c70e8c0d0e57c0819b525fc117a820b620e018079bbad5396ab0c074a333b8b203140fc5d5e3de8a9943eba8488707b17ad5232a59cafa0c8fcb71abcd4ddaf93380c23b5f1d82921c9a4bc438022292176158d92e6460ad12a78e4bef88c24f26e2d13fe2cef314c51dc197ee1397a6ce4b03d034c6b0f2dafd9ef523c22e84b230b116712296460e617105f0ee9ce20f0de0a2a352fe8dc3c1245384bf826e994f6ec7d51c24b67155ea58764db9ea0dd851300e3c4d3deda8d5bf1acbc331c60717483bcb5d82b801d2e54c1e67cdc4603ce2578a64c2455244d96290250407986eef4f23baa37ee5130dcf3ce8eb345e33cd8425ea7ea80d629749f781b87595fa38edb22364973fd8980a5bf0076d274a4a17a362f8c5c1188940ce0dec6cb769b64f9ef3a4849550f345143fd045bba9845ee70e22e3c244913919a4694caee185329789de106ce09b7550cf71c3785c4f266899ba73b8b2daffa8e19a7b1823b8f9683a0db8faccd11087cd3c7de1dc330eb1cec827d0efba3ee50af95ecb6d6987d24d5196c82b5b3353c7cd6d1df5566cf064993d59be8258fd6debe4151df52d9cfa53f91dbd610345a75e7ea9df8ac5b860797172d2360066794b800fb06cb7d45766787da6f47c1e84483aee72961f90b7f90e83aa2ef492ae377e23b069dbc3bad5a86a74c410585aef6bb5e197ed0e17c4591b5d3567adc0aeffd9a92a6b84a58b6fbedfe9f7f2747bb731805087241fa19ef46ac7cbabf13f0f5bad18d7c4719b69315459f71893134c86e28b50add9019f56762fb9135851ed1c7813f8e131ff10d1d197f40cb761b8793291acba7af235bc6191fb9c95c2cdf9cfa5885b5a38577a7f4cbceff9c839a1efd1f10f9b9246a45fb1a88907f674c51c1516b68c29ab3d4fd6742bd5552f28f82a32ec50b4e3e85a630fa577b12e1d4493b2e93b07bd6e0d479e0159feed27ba994cdce6686727a2b42aed1f7a87154c7f2fa8d0a82555d7ed3bbc188d4f3d310dea3499ac035b8e066dde2f6684152f22bb9401db9127f44fd8c2bac8ebe3de656b2ab608b8b871a64b027890ecc58c8f234f8b194c485f43c1cace3009a4b92eff96dd1ada4962004ac954159a8c913eb08589e045f75ed3699cd21f782137f5048a9b326fbec19be409e028c7a76b929f8351cebd26a53cb41b4a0265ce346e0c7b71cd561799c84877a1af634a07d75b565a31d9c583ec735a885da8a10a64f7b321dcef9d8d0caaad0c52545f6287a6c8ed41fe845e63eaf8987a4db71bd743583f0fb155234282c51f7accd8af8604325f660fce93ae3b6002116b249db2da23f8f2573e32d901571cd1e56f2772225d000ae63e93af9bb0248508aa14933e3c0feaaa16340c3ca531b36093a13df686cebc2ef909ba6bb0c2d0dbdebce5d30abd6b4437131ed6393d08309c4610a22d8211ebcdd4f29b63df18af8227f137b11e41a799b40a42aec941db660c531a86e6ef2675b14181e9a9f031aad365b78c87a5b10dc6fa1a7e26137d3d3b7c60a9fbc97c272569e0c641832866f97f99730d7beccc94825a44e6b7107561012dad81db814589b1fc20179a7fe0485c358da8623fc60c0e354a6bea445e5face46f953ac1364168258d0d9cfc03481b51e3a122faa450e26b1ec5a2501455b5237d0633b1e0af8f565209ecf840351fab2c98c6095bb07332f3eb38da29223f37ff77d317f281c18e7d0d2f90fe1e8d1e8f0ce9a521ea920ff5464a87649abbdca7e2ec197c2a4c2af2ac50c8f2a7cfefebf3df3dd866dc5afc688be82524376988f7293837611777ce032a3f97c0d64a5f19644db0833e7de230b8fe912059ad0cd77a8afbaa2744cfa6f8ef953e4342d84c89f31d19213bcbbe857c1e69001754cd507a11a5249e6a29ba7ac0e6db9d11e8da55772794eca3bce59470be34a1eda52a09a6d25e7dd18c98aac05d0ae164e3b9b2a890fc7365459bf8f57f8ec3c4c43a2104d6e56d1b5ce00215c303ccc4aaaae81fefa8e3d5450e736c3d5fe8bd77dee94c96c6543f889ef5bc94a83b0be23ce9e55b78baee68a64dc27266e0a47a37300922a43707411c702fd78b48af6596f706129524f0e4d4fb9d8f66d6917dbac071d923bd25a95c921d502e451089e34c0d134277a9233a95f29383132f697ae3f6e0d03a19d9c5f8febc99e9753e44927f977c60dff053d845652576fb6bbac33ffbc3ee1c6276961ec19b05028f19df9adce9a9fe5c0b1876ed65e7700dbc020fe34122614bd6ba1605ce8026d675e6203ddeb5da3fd6eeb08b728b637ce2b1bbd94a2ee9dbbc55af906c09212f838fe3cb25892703b4da064efd1716f8f495ccc42b3b827246954b9983379c8e3f2e12aa3a87dbee50ab5d13ac9967eba02d3dcc89bb9e30d2b17911ad7e5b8f9d86cd44d6c2361924dc88ee8c4c3d7b79ee96bf165d36c2938b02cba9a444e68b3bdb23cdc8a0875ca27862206c8df9fac702d303e22fcf109157ee4d3bd1b4d45deec54d8ce9f628647801cbce9923f2968185bbd68b2b390b2b4e783766f0e365f9863e6e8efc88dd76a0ab752dedca850c90bfaf3af26d76cc49adce9c9dc278bfa98c8e26abaafced682901db9e5b5148a44ca523953e2018dbeff7b8aa9c2941e116ec564262c32d4f53c9b12c15e41405669f1ffc3179e19df64048906307257092fc325f445fa75dc9b4f8376722a627aea1ba45340c56c28170a525f31c55bf8083faf6acf3f40d1983bf4e18dbc92f890664fb8a8b7ce401d56f6c2fec9c2f180b39c4be30e93e073c30657d11a3ef8aa6e63c54dff3f1d8fb375370578e7a61784f617e14d171d1d521e94380f51dedd63691323748500a11c64a0e370334554a4ea017ea016667e689e042cd99b12181f7e45f5bd5ee5ce0a3f05474c6256cf3efe7c364a05a56754ee0a54c7a287f69aaf2acb9a5f4b4a5211cc6f851ec584b8922e80bdc2c16295596929ad4d3ba62f6f40b063db2a67e265037be0c181c9f949b163380945a162e0e92517b460c3f1baf99afc43043e94675a6617d711d47fb14315b2f16bb20b4fe435eb604e5a7f1b997f4866daf803640738276429241fdd87f1e628bc997e244b0bf3419b7d05129aa117fd677f173217f29a4b19cf3174a0d60e7e6b4e3ff9ac2fbc61b14ae8d31f96badb291aa8ad0ea7fa926970306608d7f5e627e3a0cb7314ba42440639bd3974be8578e7e9e9c1e7c14169e1253f26104175e1777647f5bee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he5df8fc3c205ad8ddf97bc1e66e04470d4c67dcde09978369b913f7f92983713304ddda505de60ab1dc4fdc4ee13264824528042e281e11d0f536effef689c2f7c031ec2410b1864e0743ce644c3421d765f0be25dbee15d3150261dd392fe7aefa0ddc18b807354cab151bd1ce330a0066e0525e6fbb04912fbbfd335a61f01d34b4dee420e835bb05d617c4bb1f5ea992585a97e2bec4ce91c228a5e0df4d74315a42ddb84d45bbcfaad51d71cc3a638ccb9f4f91fe0ecaf8c7df1cb87033c227b94ad88baa80284374cb527c60e1973b89a537e840532da350bf3d017012a0f332baf65e64c35148f389d50d15915ed46afc63d6b4b04eecd11bf329f7bd4b39f6946a0d6ed779f6b411bd520316b7bdc6c3ee48a45f46b3c87ea480e2e2658109b6db8849ff3446657fcc232c19eb3429be6b91f29b62cc0cd8927964c0b96515231065ea31641446f5342c9c155768c9eea607e17215b64a40efbbd92f0a654d4f8ac5fce44f5cab1a97c717706245df0ae3416ae13dd7dd43c43cc439a3b4da4e3d29315c8bcddeda16443c379669688feaaf1319d9c883d189855e61f0e631b5521d6b77c11bc2cfb06e8ae6bf8a082ded737dbcbd0d56fb5afd6d38313425877325d41c7c8a12f8d9b23fc4648dadf73fa14c00f4eb2f6476436792be7b17c1d3559170c2610d32db693928baa59cd1b3e3309fef5c81932c2a42a463a95e84ff05d592ee1d3cc17ce904dbbc5cb42d247052b13acefe234ae364f7535a492115cfa7ed753ee5a68f3b7a58290c00883a95a49c5d574b496bd93cfaded5c66da85bd42c71705e4311f9870d8e63fce37d8201af4a0dd7e88d07e715a2b1057a44a2a005170b8471686d0674dfa5666f9e4c1810003ed73749e888fdf539360793cb3241dd32ef05326f2ba4d3c8c98f46cf50b209160f6294700de92af5febcf694bb70333a62d8dc0acac099b57a4d71909c1e5118d13baf1261490b44827726ef94e06f6e3c19c58000cbbee05854451f0610f36f5228591abb137a9614820d8d2e9cf99fd5321a81a2745741caf98b2fcc8be5072d810acc6016af4061ceeacc3fec7d7797551727fbaca08ff1363dbe1bd51899a5f04266ab4d7cf3df375961a2b934ab220f9390a1e9594c92049779bc1d642cfa3799645b462e77dce20da7ae56f338ba8af86b6920810ed7b7f4e07f08521a382644e100a82fd1383ea2aa423f42c87b31f885c30c991e1242c9c5611a6915fa268a23162b22aca674626e07a95670d15d58e61b6e93d7fc008746367810d87b8a4079f00a1117f648720e7e373ecaac4a2d133ef42104d91ffeac8ea742013280db27c6837a29b06c7498c1a7f597fb7393c143bbe332f07da64f2747c65c96ca902a6a602379ed3ff8f3f455128b8f6ae4042efbe56b3ef111e535268d7ccb98de01a8009bf25dc44c68fb88c69147c7ac606bfb35698f29e2624fdad220417ac962bae351eaa8311240851faeffb7768f08e199d5c6ae281358b8a356cab1a764051ed3d02a0586c1fc2871c66ecc77a03a9965ed089b0a5c6f9fb4486145e64e29d16df408438f6acf21ec62ad89358fa64d7ff7bb741e10a4f5979173d111170b5f5b0d1a248f21f0b29d509e288ecbee13490c8265cdbf9100ff195000c036e5a6f66416094705768c82f19c947d33e11381fc4ebd0b88f3f7049a223ae7a2e18d1c06482aa0c141a27202ddb2a2e0c7c149364bb6ec82f46a5164826f789b95fab84538e2728904d2e734538ac10e522cbb0a521567dd430c96ebc88321fa7e98f4637d9282d386897d423f0b7a4bc623397908e35ab02c5df3e0d213dd62a37d8a708f14f611d37c65b5a7676cc14eaf919ed7b13fb7044d743703dab7c303705de677e023c07ddcbef228f2b8cb95adb6bb7981c13d0a6bd04ed53f1bb08cea1850181eff36cf0c191a7195f58012d14e94baa81b38128646f5f01f0a8fd69fab98bd61ba1a6d8dfcbe6793a71b0a770a14f99000ac81e07128891a7e77b66b25181997f8b8c850fa4fda770783ed6e65386bbeb2ce77c3d38714bcd5411d89432de5770d152d5621f1f13064da192dfa62c16dab077dbdb6449308b1b8faa34aa931d452d91b9f96cd7175715c1ed7c312aa0f1dc68093b1a3da0aaaeb05744dbcf88eb3d1ada9a145d049857bd9a46f5c7bcf70d34d0d755f5b98471351cdd2babb39c204047be892de933b100008d53cb0cada60fa31538b50b05ec6cd5ec59edc72f6e9d0a6e0c1f35fa2ab5cae5f0d71bf74dcb8c830924196dc22da76ca8f292e438053e333e5326f1465097423f6c581ea76995b7a8f47dd031dc1b5bdb3803ba127cccf78c433862a624337314df8daaf1396234a4d9cb70bc1ab774cae53e4b53147c1c289e4f4d1b4cdcfa6334ee5b9fe30240fd72bab277a7ee8be61aa75fadf9da5a76252b972166ac8a162910d2e988e195a218633582455a47a45e0c1a06447f18fcefa75d7de3792112952cb682bfedd6430717a07938619dd5d2e7dcfe1cd6405cb6b26f1e2b9037f4bf6e443d53792f377c7ab2c53fd3b04b096e79935fe30fdc286890913ec0d9bb208df666d8ac5741395c7f85bf8ae2e5e0920f70a93db7adc919127b4bf0f14699ee32632d6b8d823157a6f53e6aeecafde22ee7e1ee60d4262128a09a93986aa3c29d7d968847442a0ab4d8d3e745b735ce8ab679d2665c3f4a2b3c7b6389292d7eb7c0ce20d41971dc97edb2bad87394c4a5a92a796d5d7e6afaacaf039a8a3cb513b47f4bedfc55a5b30c3ad95b64cf33b3e51edf3b5dcf262dd98d24a70f38a6e9623fe1aadef01513822b94d0ca36056e80641a522cdfc33dcd209db9c35cc57ced3fed701de3750785444f56be3a5265c72617bc12e15ba50d6ef2ad79beb0c5533212e809920bf39d83e2d7d4afd113776c6693a06b4734d46e2e0a9a05f0864c0d873a1120877e50354ffc018f4f1717214388919336aa80d39beb34b8eab0aede9714b60419b24d1db6d1adb23bc94c4a28a0632ef400a9f21ad532fda1664cca1902e879b3cdc2f3ac5b1c2c40b7f7b9702759be99ae31fc3671bcc28c66ede925a104b83cd92e52a453661d328f5e4ecc3bd4f59aeccc0dda601a8ab823e73518a8d95d03985699303a43cdee97183d052f4838d8cd8bd3dba0761279ac2c267be6a085d6ce2bd2da449edeeefbb21e7a0a3e800e3fe76f2955004c39a2cb4c167621be30f83e0af8d91077cf39752d408343eaa01f4d1f35f2e68f25d7d5734272fdc02cbbde8d9c690493624ccbc03cbdda52e46dfcbb6500c5e13a60fc8bc1d10ef19ca4065d2cba8dc49d548190751a978dc4fc2266d38e17a53c3af022b0ce5c89b77ab0dd6f7221deeb57d1f2ec418f132581040066ef08254064eae4bec2fcf5ade484f916df2af01dfb1652947f560d23ed0e203d26dd68fa4effb9c4d7d6ae1916014fb191504c55d3ca80452a2457aa8c95a3b6a94d4c18c64421c9dee66887208a7bcc18f8a52a56fc42cb9076918002e8684b50f4af17c1c7685daeb5388d6fd800f0adcd3af4b5ce0d5dc7230ab438a66ff019925aea4211e3ef2207eaf82419f7d6ae862b9abf888ae2cace2b22b524338db7de596e6c0fdc08fd2ded892ecce206080ed77c895f917c2004ce6da6575efa3ccf0a35ef6a9dda017340922b8abca1cbb5fdaf5539f8aae4268bd579a3fd05d7ec984d52fa5e0f45fa208b9527d5d226cbd148bb91310d5da1a2977f5e99933a2a9bf5c12395c7728df7bffbd74e360583941b70c20aab0eaf3fef157b89fb3275e6601d100e29f110749c6637a598497f19e252f897a4b9413c06c77e858cd1772c45d90b86b1d1086eaae0f60a83d5a13736a9fefda2e101243433cdc733e72c3eab04569cf8769e5aea6d33387189794fdee357cc8399f511060b009627ec7a24c3398a700fcebcf2fc475271e6752b930d6d0d4cd5f13e4b8ffabf770be96451141caf88b160c328dae935a67827b403ff56b27148c4a1d1f31e21fdec0071a0f00fb55371ab9500dd69559aa57056f35abd9f820fe0235184cd1d58c261535cefa0519a63b841cc0ecb277f793c02460396d82a646c871f0ff7154cdbd87cd190ddbdde5d8ca76f3f74fc13e8aedd107edc55cf0792509c60e6da2329c53f0041d831d3156bdbdbb1c08f3a5d1c2233359dcb9039911626f67a3307a94c257b4b218d765a637ed21d659421e07d2e492caee15f6e84a55198584c6eb4eeeee28249de090820c42829574ac78e465ede8af967e574dd344f9309251f306eb06a0b63be7ea7106befd6dae77a94e22822fbf505c68a1de74b4e44931e173ef41edbec0842e25dd10d665d7369e4122d4cfbeb608402f540354f702d4e97b373768bd46ff13028846855dc51c0bf6320d4a9bd8cdd64732ae288c77eb2aa985d80293c2939f69eaf643bef3cbc747e8bf3190bbd2dd9b70d1e37e695567e95c2b57651bf2b6fc7e6642d89f6e2f03c6b284397f732c45daca47f4df21b05b4c96b6f2a8432e99cbad17807face3d5a5874bc80a8ffa4fedc57845f28ca09cc06e98b6ad65c7d0e6a269969521ae8c2546cfb886682d42753fac7e406cfc92d1666b8b8565f380e644f8ffde8c9ac8b36579ff6967d8b80208aac3725c09e7ff8fc7d05770a61670c24848e112933e3db683f37a4ede12c44d1d2ec19c31cd1abad449440ee8034ec93ef2acc9d046c96a121cde14f86126c8e524443c16a6dfa40803edb9941f67dceedc9b0f8431ccb0a351b89d74221afb0ff947879241799bfcafcd102de45e74c940eace18906c4591eb759b31bf3029b14c8efcd00e99677c340552b40799453d9af4ef44dfda596777e862712fc39641dbeb0d1dc42e60f7dc2f3a13a02a64d6e7ccf9c6834b6ad391ee9e19005bbb4773de629cc0d8600407ef0ebbce350023558cea653fafe2471b1ee03c0ca3e0f0bc300d0d4727e37b85c1762940379d78d826358116ff57e1915575519d0364a2e2d2e869ba8b5fccd285d95798fa05be40a98ce5f0812ebd9b52a88e8b675168bc4c42f221e98caa0794d5bf6346b1cbfedb6b606cf75f2cfc16d85b4866e082994f7c99741b5d7610e3828a981395eba3c22993f6970806f414a331849753c53247a4497d8d92b802a8c3f14d5a311fac015280599f233e0f8f310cbc702d0853e679748d4728321cfdec5e1ed8c8731614820482beea660816e29a1a6ed362d0705568e16fc538d607bf2d47b672381566eb8a76156677f9c4439e0470b31e77fc67fef8fedf220bc82b11f5fa5d31ad1909707fa871ddd187758e9ac0363740613d5825aee2091dd0d18f5315dfa1ab986edf2d69fc136086119702452402247e3babced7abdf0401e037b54ab3991f039832abe9e666676cd697d137daa7d9ecb40afa982bc63e643ae6e0d978e106ab21dad9c5864aea7fb2af7f4dad33ba26f05c1800cc18bb13728782fe82706a85fe55d5a28b4cdabe2cc102a8098cf51893473d61125eeb1f63b180c6bc96ab352e148aab08fc8789c557707028736c142920aaa0aae72289f88a216a2794970ee6edbd9f9a476723730df7b443016aa2878797c01787e497fb20f07c426744615a2da2dd290dffdc63381bde670f275e47cf2b08b54815032b65a63ef3c06e9020a340405a1d35b33d974ea3f1642bdb894e7941709e3ee1776c751e5ac0949b685c544ba48375c2bfffb38c1acc0df52de9f6ffa71c7cf2f6abf20fa0deb40b21967a139;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h529a7732d0e5d27961c3bf5974da46e5f642f7b07c4f74838f4d3be0317322badc2e0b0ed8084551316a0788098c173a3f00cff01cf290e660c9adeaca52963112d098922584b836c343dde09895d7de9a9f3aef9fdefb54e220c97ccc174faa52a95a2b1765249d5917a93ba9ee47624817ade4f45d8602e3c20b8fd61953b99e80821a936eeba494cc2394ce2701fc52b7c1a2599f8ed37d3ae0317db1ffcf05c8610d634bf70b1ad4fb068f5fa0f596db7bb698ea3857da429432c49ceffd5937417e73df3c1c95c461101bf3dd571122e817ff45a3e8c145b05d7925bbc02006ee66e48caff6a1de7b495492c977e9b4525cffb28c1ec578304cb3bdac8678e959b65ed758965c3c2c042bf41faddbc30d08c73831227ea07b22e472e8f146f866878b162ce7ce38a0d3be334d068b25229821512929877ae53ccc80b405cb51daaba767f78bac35e142d29a50185ed5350c2f2ba772d1ea42ac6200f785b782f688be2d60b192dc5a528cbd4a7904ed3976914840453eafac4efb18d6bc3fe7935ca3d98da9669e837daae4d6590a3fae773d8931382303035fa44e75bebbde044afa8a34143e8aa270879e5c4f31ec96049a1be01b7b5fdddcaac7d7ef06ffa936402c559ccf2698985b5c07ad82078ba886b2d00da6c33c0983de4b5e76ec956693c31a4b2fb91ed143f50d592575f49207036625d78589df356f08030309ae08a06b96a187c2385ca4a584be04221af3ca8dc0b29abe90222ead4c702afe73b2f24f123605780c7ac93854e111d7fa7c549a5fd96fb1fe753eecaa87fa7adaef702d078a5ec93293898ae898cab20450d38979cd3f35c6357fdd7a566f47c5408724bc8f8e658eea743d70d94d3bbf1fc7e000a73e94366fa356b415502e853eb333cad776698f984860f0b0155a03762bfe00ee921ced48d5ffe7e324d4ef0dd545ccf1ffb7654ebfe494dff48cfe75a1d253a0e20ddfcd9f49dc096cd04b3165b3a771f7461600aef64e791a16a2a1109bda34b058632865f02e519488222afa338d900e7935e424108345b91c215effd6c5dd3d3b56457bf42a7d61e81cbf2c6c2dc942d85e0e902b8eb60a9a3bacf5009a3641b1367557df1de6989bacea6b3ad921cf79405f3993204d6694c40de187e7dbfb53dfcc2c232de78b8b4765309f90b2c33f3d89d226ec4beee1ad8d37b59b170489f4ddbc64c0049b90e74639d59bbe6bbca529dd82e923000a99d8fb034816c0c0769d4dec6e64795d0411b6b4fda427634705ba0b23fc4de54ee5920e43b6ccdd1ac32d5f70709f2423c4f018cd091d57b5f49e7159cbde200148def31af2a59c54d385519ade70395e4dd786d04a630094e78475bab205e15a33b431334669852c9e5a2da67fcb48075a24f5fcb9d5f200c7d99a280fbf3697c18f1e5265698df99535a2a3b63e470db022dc96b40b4cb503d9c2da2d6811e071a3619085e7f538bc07cf492fec855e73be8bd753367c8c21690cc1c673ade2e6efa655a981c1bdfada22af05230766fdd5f4f0c21a26abb8455c2d9f9db0b5de2d492009fc5f3319c4f443697bedf93be0f7705eeb208a430082ace259232f45805a22905e87ce25ea2db8445d666e8145a42166bf93b00bee08f1aba5d30a04d247add793c323605dca6da5f34367d370f92320352c156a6ea38b133df0e0d0090fdd478036f05e7f35d81c2daabd968159f8926d86cf12765032469d471346d7ce743d998001d4c2e5b674fb256a3e1f616172b6b60adf4e759a699966873d7c1e88b2384b32dff18a659c3c90494f744bb85ada8a3bbe39d74fe9c0e822f17e766b32736f280369c2293c103c7994d79c2ba24b7dfe1b8ee9f0129367620d191dc996d0557c260ea45a4212b24b9ad7ebbb1966d12d783760b7df52a29aaf39b45696641fcde5d3926dc696e7087983b73a5e1675345f70b01edddc611ceea8f518f3a32e84d178703070bd374637b711816522df892630bbfb638e28595297501048d02159e37f4c7ce5e329229602c6604918c63a2c989601afb8299d4761b2d35480e3e3c2aa0ccd3d512f87948fec7409a28732267ae7aa5fb7bb545143211774f6eef9f7c543855da2516feb0fa5dbd5ac68b8ae15319a7789ae640d44427085fdeab34260557d557433aac2b6fc5df7043e9db213bb4c763f9e3d9a4148f3bdb0c6e5dd7f8fdc2c3072a28bc0e3ea2442dbb99b6f65782dec24f75724b4f87ce863e57a3df5558a17f6430193d1742bcc0a4c33558ed7b0a8d9d374be0b3c88dbe64c64d2dc2865414223f2db6ec0f2b937f8f0ed73ce2416c0102a24fa59721aeae8f7a9a5d0b6f456b4622f4acae590c8797be5f4809c03eb82dea2fcf16b69f9e9bc39c16ca5156e0f9ac1bc51db9c2a8befb1577418683289d103419f893804c5393f2ec098f8c94438e150302d8ead343a97c5f5fca9fbcfa5807d61b4f47a15c08a77ea6603b62d8b5aeee0219c8947a4f72c5a1bf30b8b51451a3a4c742745851c17bb121ca59f37c4da72ebbe4000cd822d9151cc2d5d1ccf83acb7f33a0a32ab1fae2871d7257e9ababee4d717620e65086933bf4885d48a5b32289e5d535da699aec06c1ec5cdca24fce6b56a83f1c1b58c1c97e47d06f003e997d2af89f5d41502dd33d824a582585ad5fcd5789ec6605f869c210dbb4f0c3ac1c1fce5ae14f635822ff689403cb1d91ea58c56c19468a12f0c1a413f0de0822c54147389b1ced65a1a4c6f17ad3de4f9b79edb83df677a6f828a71fc81216f6c78058377a1b59416d72933523fb3fb89724357aecb5b7233b0ac8b4b3398f69e84b48f0f8d7e00e3cab39243c3083d589645a8f582e1cb11c93ecf0ac17f34d7b7e360c57ed74c5cf5a5296486947a4e3fe03cfe4617dfe82d192544aa3966c0f1d2a3afeb91bc5d00b7cdccbcdf730843bdb7fb25b4b3c0599c7527c5bbec7ed95d5a6a3a770acff6f431dc770bc5a645173100c6d6da64c9f82d131375aed177673ba30de7313a6a8029d3ff1b76b3b9d90446f4ea1579440ee33694dd0d2f32dd2907e5bf55d1e0a9ea36d4a991ae3242e30c62090a26454402a79d8cc7bd7d0d261a6d197a764e9963d3a56a05082530d823d442b2d5c8857fbd097941754bb9ce903432cb1ddc79fa0f7114be3715a7ad5327c8555b2d5038dae93d1851f7c1e5ad205d2dd127082d6a90f6f39f32c9435495e6d29e59a5a8f6c14a95a62cf035c31a254ba9dcb208fe9f65995de606a68c1a48f07d5a157577738f64a982e6c5be572093a9f969cc4a57e6217278cc6e3e4023b9262a696a358ce6eeb4b0ad55ee70e48685140deda8f8f6c1e4af60c4344ebcc8b4e943ea1d113f13d3fa8b5467e1968d416b85947c65f818b1e8b2107a14075c25f6534631a179eefb31c36145889e8e5df7768037eb8294a8202a9cb68227c4cfd2435f48e3ed574bc5303e76c5c4a4ffd927259c97b9a8b58ac5cc1426a0edd177e6d6964bed2b3b42021ae49fef733cc43d9eb7c0c7a8098e1b07db6089f9ade32efef1777094b729389252004bb5240dc69bd616bdb305f68c8579027b2e78e20f8a30105c57f19f31975a8235450d6940b5fa772ce2ad40659e11e7aabb8140640adda8ae524a3a2defb0452a589ae51c20454b4b576a0eea16f6a743d33c2ab22bd70a4520692c25c3d709f19120608478b43dc6eb96e3946e8dbd9024d13703148d4f9ff5e872c12418a200c6675ddce4df7167483eef34ae1c108ce12a00dd52075384435aac3dc44bb48fe24783239dfbf397bb03d9ddb8bc5837a19a15bc8b1c841c39ca384c2696e3988c2d32d0e8171de37f9abaac7684411d3f3ae4f78769d754ceef43fdce6108f05b65bfae24ccd7acdbe38f6ec65b447b5bd2dc38eb514915567e42b14bb5b076028ba254029ac5e6704a61b7245ea075279c28c447203ae777e655e98244db3cf30712e111b35827008a37dde2f012153c6dfb0466cdac0a737b625818ea86e21c80e84adf3c7bf59cdc7636adbbcc2cc36d599c2a1ebb000a1be8a4f1f6f0a93fd9b547d2f857353827945b8d669cffa8d6f45d9886b5c3bf56059b88353b8f6d48738ce6a6219c4f61978b36c73e267bb235cd35251bd716b7532f15ef1dd7cb7ae70d3ee39cec09fdb7285de9557219d853882eb263b20c79772f210e86f51d64656b99d3808b7d5299d9ff0a843ec6dbd51550e95c514eb8255e2a577011cf19b60146c78df7288feda2a083e487e229b1a535f3e08206d910f43130f9f1e3e0ec728bdfeb2acd60fa13a52ee1835b1d923bb6ceb6b2c1692e2d4f7cbd0ffeff00f59d52b3db13dfb779e1201cc410414ff0575c31d78c6ff26822a311554e122b159c045c096cce55365f03b01d2fa466d46605f7354f5baebbb1c63e50f6ddadba8230ff09d68a597c00565b61f687786fd51731db1b42940f80727edcbf3c225ffa78d2c2f2c6823aa806259478b576972c67df4d49706e6a9bdca7ffded2d9e900568a2408be36f8ea8d6e50fbeacec75850a528ab775c18273568d78ed5b3768043dd70c930dd9cf77fdb151f494e194daa93ff2c8756948fb6ba5d745eb339972254e6307366bad152f88fb18ec3dc3b8aa7828f3b589faf4e6f19bf453db5fe9b7eee7d996e6c232ba20d1566fce9c45af3f70f3f5a956dcbed00b9c6a311f3ca80fbb376d872ad37b2c1383fb57bc266595ef19d69111ef376a8405d1937796fa955cbcd5f7632d137c20f6a2d651e482897135750ed91ac90ddeb8ec1be35402a68409d64b78f3a1a6747fe7b1ffb295246ae7f1af8b7e7ea70aa644a7c2d0c61f7c743a2c4248b8311e188babb49276e9f2711b3f2a73ff8d89341b4a10780f9063d21af1017a70a4ec8347e3aeabc94b20454bcfc7913e7a57f5728c864ce0724013a52c13bc0da1314e290d83a1b7c0cb40a16a6bcc3f3ec43c06c30faea737cf156397d4afd94051e2b4530886c9217ca6b3f2ca929a153fa8f56ed6d6426b10e98282397fdadc5be0f322205b973adc7a74aa6e7dcd85032a66ba9e747074305d0f828924c9cf34fa18102e43b93aeb7429847e8f03ad0ffe7eb42110e0249eb94e43d8170af7f7d85d53413daf21eb04a349044242557573f8815f40cb322c999cca26a4d94da44b7be76a552ef51c4990629f98d61c1712ce267b936244c51e336db76bacd867d0f26674ed22cb8a84036d6318eae875b69188ba070895c2528c3d5e83721b337d7ecc784586835e59c54d1354fe6fa70578a05103e487b0558d5824efb1f4e2574b401ec412f19f2d59c004a56a7f8cbe1b48299cec53b284bb5549d5ecb1caeb08fd4f0415444ae05d207534691838a5d2d1996e707f33522cdb6fec1696b5ad0647fbf8c0763145a0740d0e05b7a2ae0a0dfbbed683986380b8bffc4c4f8442ec48e1a85ea751f8f93a2c9605081036e96ba26e518ce7f4c8d1d324849196e78eb315be788d89d0a625d9b55f76b13f03128227e95a8eecfda133b82aeb9eb5db58c49e91cced57276ce80c5556701bdbf7b9f63f2962c178cfc5420107a26fce59c6dc02a7bb2cb017d2169da666711e1850c9e2aba8b98f94f2115a636c8a8998995200b5ce9c22dce8fd635d18950fd416162c3f60b5efa7cb311a6fa8614b7540db9064756e3f7244522b06403881899c215364b6209675034117da4401d0c56baf3ca7888716f494815ca1d2ec9387fbc6b04062ac893090470f2fc771f567da2df7ee5a81eb4b67af82009b565;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he15cce7af6cf16aa59127f129c51cc5732733a8ea137eeb1f2c3e2b8bb3ca6baf4bd3963dcebfde905eca7e4cc878eb9a8e7cc3e62a42bdd7622f9c0a575a353100fedb3c2ff9de2906243f7d9edbdfa7d0763f197f039e5a40dac66cda47470d37a69cec0a0c60d424e796b4ded99912cf99e50c748ae54f816e64f1e69007dc4a1d156ca7f9ebcb17df4b4089985b1239ea214c40fed7d2315104ce02014d52f0f1b3faef8a2036afee4d9f5b495a365f138c77f4ad3399c69bd27f872ce1ccacff9a0cf1db0838829733b16f3dda46e958b79610e7f37e661b867db88530f69bb9ce4d58c4ffdb5783ced83bc747963fb7b28c3294445a0c06b577282ed8a283d3f1f954ac9e258cf3a2f0a45d458111936f92d2507c42a3bf9d1b1c67c0f693b29bf7456c9e41ea2dcc35b118214b1a47dddefa4c3489c0028077e407745b8687b1d425dd0b6396fd6a788df8e125fa363eda2b82c290fc9a63ae6c41da4294ab2d5016b61d6746ed53300582937eb488d19f526f7b1ec3cdf77b6d4ae070d9fcd68fdf1e33abeb89226f8815cb3932d1dfdad089347ec2992972f21595e2bfb5e784ac117302475da255a6b361c8a13f4789bc0d4dbf8beaf03bf092927a6ae545add4b6873c12466ef4a2101997e368855c218385ec2599ea32f302c6619e783897c593937a658846b57a473f2a6efb0973a4afdc15cf4ae5f44563332b4f8942f4e97aee62bd7fbb66c4c79b93e946a9de8e1f9341752ec0fd9bdb5effc325ebad9f873ae2799147292da3bdc8fc906b84ae56500e261596cbe9443baa0dbd62ae7062ec536fb7c36e068568151224c8b9a217bce8bfd82d556afd7264973b8d6a55528751458e838617aa5a838a2fb257eda614a3a93faa595a6b44d773e40abc6f3777c6bb63fc6790ec9fbddeef4a7b3a2801c01058aea60d41ba8169e3e95ba176c216a297c91a0576d74898d17ea266151b6093d46229514e1c9af7c962c0e527ee2425ec2a7d090ddb6ac5481b1bb22f96c5f8e0bd207ab91f696b4046c5cd9a98b25ed9b6ade96a85e704f9784a69423b9504dbe535d675813647253a17c18004c3b7116c520b8383a111a6c0c46b4a25644fee329b8b317d21c1d45b1a9a0286e14f2575e244a88ea2c4662973ded4773bdc102962f0c03d9146c4771c6b68b2fa1dbc72e6e0154bb6dfa90e5d51333325ab41055182c43da0ed20841c8b5cd6a412ab23982461f2abcb35b42a6b2257b295c4f5cde2f9121f55908df9435808bb22922f8108c9e1a96a6baf94174ec9d600652c513afdb20e2ff950b4eaea75c2fa5f7ed9f79ef45ff7f2a539628428a18be489575b821e0c075283283c377d736813ac2e3bdcc42669e37134760ee377ec242efca4274a9692eddaf8f29cb39a2a03239fb3c0c583366c880eb68b724f7a70934e3149e1477f32894abfe981197201dfc0cab14e6373dd96c745669039b1bd4163809f00270513c3206fd0ad98089a16e612307cd6365e27b40fa05e96342087e78b8c9286059d9d0dd8ec72f5453e4b0710031508eb1701e0f11ebdb0aeab52283b7a95c06db000f7c19d92a540104d719819f553b44456dd6ecd72c737e341578d39e4b76bbe30a8c036034bd218a022ce79d9b815cd261729ed4d8f271e2e82ba5afdbd7305e14b83ead7318125657754a1b207b25f8ec5bc9e956a49f877941c3323659d154c04bc248add0b763459bfa83747c0e570e8aec0140d621220fe9e82373ec52b293e2ed118b00d4486b8128c2e21d728a5288562e4a48b7761248c382294d4e96f165cc762e71902cb9168d3d98a8f4d1b3cfa634a8930e28d340073674a3d2e1eb82dba80afc542bd2f110489c615737984fa481559552936c657528e4fab2fe3c102e47b780e490347351ffcc29b8d453b2766401a95f682b76dd0e41c65bea2ae660fce3024f99fa50e56d9f8dcad78da1d4b7574060fcceac1606299c5adc4fda270040ecdc140e885215198518e562e2c6dadc6d6f6ee2c9ba6526b1229bd582f1d1acd22fb1c8751a753b821dc61b686216c329bcc1994ff6bd44aae30b21c310d996e1ab313e7b693607db50b58a1563c38846c4cd53a3cae698b7be9db1371f6c68e922ad73dfae6c945ce5240499ed14c2f9a782330568a33f61b96018a9007b4c7e89244d37e797b1309bb82a65b0714e8eca29c2241c466ee27b73ac06047b0ccdf21e38d6525321687f5fb97cc8d96561b05a540adba24d4d5cb36fdbde8234c5431eace34317da135675affbc74175fe63a9a562a8bb7c6eb3b13dc26ea584911ef549b3b1c586b4682a0053edb29f350e3248f9f0762c441ec37870065ca0056d0fe4419fb8461fd202715719ce910d3182acb44684eee249d74c3ad9b0263bee6a68c218084a94374c8d0dfd96e90f5612440c3c4783a12bf5c0940bcea5d632f155de87d1a6c7f76ac6316a63c5f72be634e795c8feab49fc56232e438165c731ed588e75d4e4e227b55c9b18135107800e7d3fa3f1816982d0c14aefa4f4e6f30e8a17ce9fdafb4b225b26908b09d0e441cd50c76b98f9dca20c692ec822294417cd51a53fc82a76b96c7a9de83e665f952d66d313ebc68d2a50f7262bd7edb47b48fdc26e65a76f395f084a98d7a4034360e76809924bf67ba624285c3411c9fe7f77e0ed23c86a5c1f22188e63a40cc6e33a007436c385d8cb88b46a6909e70454209e24262bc23382cdd2b3626e2b2012381dfd9187d43d55f1c70a40cd478427e0ba727904e41bc94be2329bd401dad909ff8fbb5c5b6251083291e6c37ef30bbff82271297f1bc4773fbe008c8a44a48383abed6f42841e791ded176928e446eedfa3d44b203b2c8e47cfc01ff0d65aa0bb7c6475d996ed5b5630c0461b1be57260d1ecb1d37b704ce25a74a8fdd2e46b3682002a18cc339408f7f15c592fd9b6c6df9ba4735536154dc3ab3aea2731f05b69065e13207e61874c625e85e462eee6328a53ca9d022548536150753f0e603a20972b1bab8bcd3a8d886d7acba3e7d4efba1e8d166cb5301da69715184f906361c5c5832e097469284823bd695be717dd47881a4a83df84b147392d4589c6256d11f739c3c0cd98fec7157a45a5789eb1a5c7938b0a638f7873108ead89743ca2b74969dd80338628a9bb7b23c01e36b06b95be237eee4aeb2e15dd44990766e1efd6e0edd2dc79c65528f44369579ebe8cb26c155f9113ef7764c29a3ac5474c5532b41d6d34f98b62014a8d57567fbfbfc0d40ee7fc49c1d2a99541527d9b3ec1969ef4b12e0d5b888cb6f7e87854fb6c1814ca293001334a1fbd56548d904dc0c12d8d8a13629d1ea5b9ddaa285eb90f5e30250f21cd890ab4979bd2e79043906a75990325dccc6970c02a4b5093f7757c904c513c51697b16390d718cf7b4673c0d8b88b0986c1b4edc35ea2137d01c59d7f9bd507aa032ff917af445dbdf4848f48d6f7a3a7135ae9c08964ba2c4c482bfe4dd5fa19167d401f8e77392e793cce67265cba0dfd41d750969b2f3cda3bcb67ffa3490f2f09625465c0fddad3e54093882f0db911ab6a1fa03d4dff4a3bbc64b339ae2aa17667493bbbc8dd543a81d2bbab27dbf9a5551a8d766494ae531f7b69d6e6e770cb7532ed3cd8bee7907612b776bd7572973c5320bc33d9d2fbed7a1eb172c1f06342daae1c406878e133197a5486a3a76b234a3231fb132dad596845ab93963464038a1766799786f730570560e90739fcd37b2213bdcb553aea730e06e1d7899b5e63693de0863d44b667f9bf81db155464ad0a698f2fd68429e0b1526d96e0d8fb2855f19702a66053ad6d3ae91315f5bd4fc96edcb688cfb9c681b54d5f2a412e1454287e5445bddcae816b24df8daf41ec743a136733b8e11c8d8b875683fc3c5b922e303adcd61e5e3226c0a84a4d5b53a1eec12de171be0ec3e699cbc46a13440d57ebe56f34c671913b571e3468fc4e7e9bee8f63166754ab251cd648b6d525ead5a34085ef22f2a3bb775039b33c5e32f97f552dddaf3c2dd218002f137b193a651f5fcc5d5d577f2266389dde8e97c5182e967046d9a3cbdb3af3deb2e67691db81dd23f90927e9605459ac69ec5c8b09e40bedbed0b9e81211568a854ccd63ad039f4c0eb2a02fb095ba512304f563b3a4f0099c7e038ccbbcc20e0190680ad94e2da1b3979f31a115ba88fa21ce00e70088f4bc96b74832d149d5eb97481d7ba52444d4b618f8adb4d7850c0a997586c027aa2c5b380358877f43e152291979e7d7190a72ab16738f0d10a95331c82fd44d8f4efd2688e06f3ded263569c8da1cf6b455000f35f49216291b5b91edd09339152b0b50ef3b2ddf5a94c33be10fcf54709dcffcc8b4aed6e5441dd5be36b9d987c8c98376428b982f6164000281ccfcd141a4b8d5433650d9fd154645f713fb6e19535681e86a67ff8f43a0e3a5eb69905d60d718eaf2b3366f1ad1d331c37b1eeaeba9475e956268168e5280d043ca038001e18b457c67de11cec19964d26e5d4c67eda96687ed5a938ba6ae2c582e7c52602959403dff9b7519cb5bfedeb75bac77d7765c0ce2038c4fc5a84f77c05720a629df38ff0fe22d4f8cf6e9eca5fb8d9546f9eef5fa47d624c828683cc4719ab3075ddac2b11880288c1c53902c8c6cb98b63ba620f9d31c8dd3546fb4c1036ffaa929562b492281602acfbe466e0d4033a7347224f99e7e3484ad9af9e39e812eb597b25e734b54d6af6b595b76a0f8ce1660b15457da7efea5450fb1e4ac74e23ad90f16232080f8b95e022a5e96e5121274f8c1935e5f633beeb217123369acd35ddc1093d01a753b40922a3a4403eb376faa4ab27c260c069e0fcd7f037ab130d4d9ba55a0064c1c7941404b2cd7302a429623305675531b53c2b5d93e1fc2bcda926e8bf908cbb31ba8ff3ff1f7c6c325efbcd126b8ad01d0346b17c94813fc289bae4e333cb721a30f63e2694e3bd47e019fdfd89c355afc6fb0c24e68aa70a16fc1108d779b9ba191c62872d9dd611edbf1dec577d0d72ec595358e64ff317948004f8e08fd7f886e0a7abafdcd3fa7cd192506a020a589ef9cb808252503ab942b93c37c6317cfe19728ce5e6f2e51a554a392cb83d9662bfe590ec7b677e2180d010453d4329215755879e5868abb7e9b0015bdcf7aa61375d13f9601f72339da76b52bbb7c223c39fc5b7e3c6b4021940f1cdfc85d0f97c29f1af45106d8c5d846dbd5c637d02ce6614333d26a3b5068a7ce86e913a2ded214149052f4581bd9483c5c412e9098b7232c5377952ddc5fe33f4f6ab16745925c689bc1df70b24d096ddbc1841d536c70a20c26fca67f3925a290824ef330312cd3fd71603cad9e6584e5dd5bc09303d26ffae60a9b697df1574b472992cf0bfd755da9a3be4a5f3b24d758945210532cebb6fef69029d082d905a83e2d9e664872e74a3d88bb7a6b44a73d62dc694f9fb89dc253dafc3a1ee7da6635e38ba905a35901b86b6144c545b1de212fadfef2a0e849c2011a8095e67126a42cb9c1de22eb2d83ff271bb131032b18e4520cf0c9547218cf914f3a933a4cd5db8c37b7402a665995d13adff3512c02fcedb3e15a95eb0383e721a5a79b7a4c2f87f389cb18302ca4f114877ec6d55e868d7a77765a296cec242d3d0d1992538ead8065c8c631e46b185df08a1f478e7c491b857f9e580fec8e379d3e88daa5cc92a87e53f5356fd939c34a1134413d9ca1e3931bb9be51b507cb6b13dad78ec9e7dbd9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbe841edc907e26fbe0c4e2736882ef054af7c1a9b10ed7d1d1021621bcbb9cdb189d615723153d8d57201c458ac69f04579b736af3b2b21dc6b2fbddfe2e12651abf8237ea2a8f79726669ed11213c31ff7e3940a08a70b9118f8f25a0dbf273beef5af265a2d335f24af0aaa25d51605437dd12c2044c41747f8de3dc6083302995abad171b9ac5ac07d17d08c69cf6c683fa5ad32c36339301c4490cc7808a3e9122f61a758fb6481f89a6d711c5ddc9f5205c7d45a69ecd84707b9112591a110a421ace3c4cf31939a28f6a3f10efb05680f6ab102285e84628681815cf7d6a6df2139b2cd0b63c1ae0374e01401bc4345ec0f46326bb4390ab11c0f16817268863b4be0b90df68712b2b612c77f0f0fcc808709b6dfec004c2036e7129dda16fc25a21fc9187bbca3e5c47195554b03282b09e9e2b26ba3a6f7e62151f5c3649b88d83570dd655cd67f8bcfe8906e00aad8cf73757db67e93662d813c8974f2cbeadbdaae69c640d9bd029fbaa757ea5acf52e423e6641c6285d8e5576a94e9902756959dd13cb95946216f3b21e7d76e10140e88c735b76b408231a8f41d45c9af50d1c2c1f0b1d9a1a464f4241376a2156042b3e8c7bea0b448c50f7aac04be6704836d4853e5f684578f0bffc1a94c3998c4dae5564b9877a9042db4cc8fe04866718ca6d75f919e12db593d66f09a1bc6817b198eabb4f2a93f745c77978497e798c486fb8e415bcd9ae84712adbe0bf12ff7f5fb9ca7dffc0b6cab346dd13aeb8c742da7859eea4e34ceecb1d0870b501c3ef1a672786f4fe0093c1539c338137097a4aac95dbee38335012143901e4749c66e288ca4cb576178c29b6444fb764f5e11a84e989f7bb3a2ff1b92725e00cf3d356b233b424401c7aac04957488587a15ae23e6f3bb6ef9409c47ad00295ab108e57b266875d08034a194b72db10daf640c0fb0b315527e61eb1e454f12b073894a2a59ec30c657db00e56347456cd1bd42a2fc0e88b8dbc0907d6344e083f67b9ddacc0471845ac13b1703816f299ef7938d865de2f14a626a12cb4b149723db48e10db410a79dea6dd0705df38d536b01b146ca21f61d9b33620049374a13a22b7475603f8a341e883ab3e5844d367a9f93bfa55dd4171ad5d271bca255a16564ed69a8b6339e641da8f73691358a74ac48047ea4021adece3a74189dcb9a2e282aef542e6b72c9c28a0238a329766e2594ac8b9b9f9257f31ccc61d68eaa9d68a3af29f50cf32db57b68ba24292a8fc8a3b678dc0cf3e8356d8b1d0ea1f5f6076446e68fb385a9363a62972d874b99a907b83ccf809e94e216999f01f0484b397754d20f4966564c44f2c3cdbb501c03c55081a6d01709f01e96319f16c952eadb8585950525dd5aab14870cf8b1ca5a29deb65681b0815a27f56e3fd516a54acd427d5c8f73dbd33ecf2d3f6d1f8a8f62ba6ccc39cd78312be26229d0ca228b066ec7872ca14e89802603ba10cad6db31a78276fc43e39190576922c3792d0e1966715f839004e0ad6f77d1ddfbca27115c417b5a7019c7109608a42a9a1bd86e3ec8226a09c0a130b98c07f0a0bad48c24339500934febfb2a3c953e3ec686acc29efc4974fe8046a919b7e0ae023d70ec4ba6fa42a0ed63174832ef06185195b519693fd4afc23c18498a11a12cef36a5c3078c12aed4a2254a81a2b1028c6c411a6f5227eda910693a3b0dd92285fe900049abaacd44367a4cb9131ebb8ce0c6c6aedf61c4d1e2af14f0ea930343a3fa45f198ce17f214237bbc14ea19458b9c1b2e5434fed73c70335729dd9f3a225dd0643d12175227aeb35f010ae7c7e997834de3a0a7c1adcb03490d28d2099bfeea6e03c2794bc8ed7aa733ea8dde8f5f7962877c2339e07ab29139751a3a2186c00696409f3d2d2abb5bf12f19781b261d832aa9f118b3b61c23ebe6a7d2d30a3a449ee1f5808e1f1758c38bca707994506d2c0c51d47b64a46e552539051c9a03f100d47c1f9a55e686ecee6847354f1b864fa5c7801ca4ec7f2c86d05d75b7260fb4dee5fe1ecca5b8d848aa83070a40e87eb4f35ec59aae0b0c7c5e6165b9bd74c3e73763a91e7484a88cecddece1857abff3cb81d5f932708480104c663e67d243b64fd199fc60a1c6c2e540c5fdaafb811165daed1f3bafcb699b7e7957527d4197e1f73f03c5043cbdcff5714b38dac3c4833558a8d10b66f88238c7b7638817990e42c9f380ca7e13815ef18a0e77984492c0e59bd4da09b0a3dd8e4a5f714b75fbf0a2f1692633810b05aa8c3f2f0aa465d2879d92d1097dc325d04797e97fa9afe9ff81277df268c8c41de0b9e3873599ffc1f50cd367ca65d18ed1758d99ce9f0fcb3ade4e245eafba615b81e169b5f19e4b180c5dcc383681daab6ecbf445709ed302ef7290be313745a5cf9ddcee26062c1e064e9068a2f6217c8233fb86aeb0b9bb6afc2aa37f88858740f253e5c422ddf6c0e89ebe9951450bad61e69d32dd8aa2559c0a31f910deae6e003ce88b15c71e29d170aeaaa17a47629b3d73afa41c3bf883161344df134f3b16448403a770c42174183ff0c55ad2236ca3d59d56ee38a908ed98f7a3ff34fd69f7091a3b7065ecebc48b3f1e8d2e2ada2348768fac49452c73663554d5863d706946aa458b454ccf8a3f0739291d8c78d7bdb5e51902e444866df273afcbe060ccc2e2b73384c73e6b581d7591b4dbc34cc964dba5e43700ed763d433358d78537479cc56fdc8a1f648f04132ee5edf848df936f795b20c801a32392d7f80804c6289cf1d7d10b311a173138820df07b49ae0af736a346de9815ff173d7441fd88eacd245575045db079960f23b6d91da28bc9c344ca90eb714c5923c0dcb4d1d6fcf86dc249a50bcd85395057465fde66a0511770bf03b744a897438d1dbc7985e78ff28373e79d8c20e653e2f89e447b56075fcf45647bf0872a0960db564146077de4a42752eb93f0ecd1d994bb0600a6d5313554c0948d5547c18f9226bff6aa379346e9640d1df673e9d40efa9781dbdebac97160efa39885565752bcc16aefc3c517321a9990dae67c158c2b3a31bde88e1cfcdc5dc7a10697c2e5fbb92d324cc2b0446db0df4df45016932ca2035d53890f7fec2484a956e3fcad1e9433e4ed08bbd7677170f2a46dcf1471cb821095be89dcb31b380e45279f9acccf49dd75dc157ab72688e1ab38385a976804bf614a16093af443758e679c890f11a70d33131187134a7e56682545af4c2205abd769bf385ec72a665a1151b7f1ccb9281b97de3f09ec8e2c23ca4a3aa15c678bb008857d7e31cd25ed97b6e3161a17a82dab5647e4b8a6bdd170075f92806a7c5b28e77a2a951e001ecb56c16789c613f6f1bcb03769ac24f1fc58a2653bf281089d97eac26a945458c32666d80b4a25923b9a4aa98cefc7809090ece390e82c43227ae946a4feea9afe12b6e46a421065c664619faabe80a7325906d2c06824517f1e39d6a03e0923007a3b96fed758922db415cf06ab3a1a3f92f169584922fc4fd93a5181b0cd0286b313e16c0330f534e2546f5891e67b35282d6647384652235ad4aeb5a41019dacc0272aa4bad89b0edb575ffc4725d44d562c9d02b5c545da01b90a26858d4f73799c23d8a6571672ea22885157e0eb0c8c426c78ab8528ee679ae94108036c976abd73e7b1c58c001853dc5d22fac01a08ec2143178a8fbcdaabafc96514247bcd494fcbe579fb21eaaf4817819e3655282e28de1c996aa4216781c70aec03f93ee261ff9262fcea5b8b7157fad4f149f9fdd7de38a15e338b815ed8559095c75d42d2f92bccab35ddcbe208287374387965dd99026513a94cab84ec3483386027cadf36a7f1949d1b4222a3a2c08445bec8a858e448b1080321e25323cdb9688f4d3715da9ea5ad2c33350446f8d95d468d741932213f0629edde7ad2468ce089d215c2ab1fddd496eea92eaa361a9cd9543bb5cd7baa9434f365ae9c98e9faccf948a1a431cdecb351ec8b897bb7db47abf890b2031c488f808443783b62277cb4d6cc2d6623f860aabe1398bedf43535f94a73fb4c07e02122ec532902f5782df93451e561cbea215613e232727e5755878961f14dbb191be5d522a2529be3d33b558a5bd39ad680c11334c78ae01674999a98b7b2220a2892895a30eb72d5186f60abdbe2f47f3ba126b00d599838d590d283f7c8af1e5f6cd0879739e7996284827a66428d3f8edb4f840feae279ce7f7ffa3f415cee02cb7e02496070811f5b3e03574575a3135585acc450f6dd7c48a97f9e4a7df8a73e343c65489f510bbc66698aa31b5437ef88d96188218b3ed9645627c72650d7c5b08f5ef78025b7a70e7e291c2c6feb1f08db19142e65e6749d934d68ae368b2e27406f1991d860789f6928caa6eb54bb2ee1cad742e2b90e6882a166251b88bf213087ecd479c93828a84014609e9abe178de0dcbf019b0cb7b82584ade43921c9a544347f248a345cc0ce4dc17cde5b7d646febacb466925ef78f64f78e42c22f765f42e7255dbc6f213cc91769605a997711517e7aa7fcef756e01600a54cfdab048df6045e86a8e84bf9309a7373167aa0b912bfd7ac2582c4b3f1ba5d4268f61d1a33d06adca70904b4a5c8059245776099e571305c6896fadaa6c828a1b286b56305466102d3aabdc299f2ded4a51f6396c1617c12146594ea377c7905f41281d215091ad20830eb2f81ef9a450708085c1ebe054d3ecaf9047635faae9d0f7c0a1cb7a1ddb9206c7682f94cc5aacf5b316ab6171794506f3a1fae26a26f7ffe27dd184f6a93031ff2540fdbd7086ae7128d50f176d14defc74108f7416fd895a20894ed4083c29aa98213bfadead97048fad7aa1f673e60c7ccca2dd7b28da94bab34e7c8f46df134c51d39709125a69e31b198673a8839b8dedb1d328c7eb4de19eb0ed61eb98986d6d367323fea1b4b4955e68bfab2afbb834b0a9f388d068c9d0e25efcc533aa412f97226db4e01a615eb73e772aab34c1c743b0c7c60e7cb968def44556e973c3630d0bc49d8489235ec921a9ad15e0bad47380661c55f27e8599fc62582e188197a84085db2a7f2ad5cb530d07f335aa56094d486059c07399ff13a0e102a740fe68bfb8a1946e15e0a2cb8aa6516ef3b05fb8ecde6b3250e0bcd06b2f3fcab3fe65972dadfbb06e72fb019a0f24ccfce978d91ca159d6b5c2e59012e248c41ed173da958114b1294c42c1a45a2459e639601416ee3558f1d20f266372538cc1de4be49451814b9aad47ce93c91244e29706ee2d6ea798be728050cb8043c50b24848816fd899175fde3bd8cc38403e1f5cc5e3ccd724ac2c49a8de1fd0dcc14b9d53193ae2d8325516539ca5599bf9db5f93b0f8f1acc40e9589c7ff7d2c719c82199897072d3d9b34103505b3d1279a296c6a3b5933629cb4c9a1ebed46bdc5f363390b795e33d00dbd82af39f9ef078a616a86551e8df0a99abd0459e5d2d6dad19335eb0c53c1d9eee7cbeb2666e97831861f82fd2b65d0584f59699e57812f9f1245893aa3481f09531f313875a75f5813d0378687f622c45374a84d74600146f4be32297a386175dae03aeaec9553314e9a00f7cf9b17e4e385cb712f8a2f6cd68cacded5c7e2e1cdf49ae5cacdd460e4cdefcd41f7e643bac649f71f64d927f7d6a0c07b958d765a5602cf6952237478a93b9ad6c5f65303647a83882b334de30e6e82dc7573b55d97dc679b11726e4a98a5770f0144e8b5049734b43b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6b38e167c274ae5a8675caf52560a63193159dfac81e6834e9cd7d029164ab36761e1a5d0daaa3e23d3e890e000db966c04de82e8687364f47b439c33f9e5f80bf7c46d09d7ebe6000f5dc5bd5e786f7df3ba46dc4f450c8913232a5c32dd4d5b0183e8a7f1c9c17919f07e08518c46c087285c7360babcd17bb7d62893fedb011e106f15aedf4e525278e19a9eafaf16621d1aec0b86ab5144dffc23f89892468a94a5244e5bcc6f895104094374fdd9ffbfebf5e6fa0407557328c1132769f3473b009eaf6cf3053c9a4ef0f173f679d587fe6185c041ae7dcec49da93fee6f9e7639aac8728f183aeb79c968e0be15eff948c0827bb0f401ddb051d5a29f4ba8fe13ca2828eeca5324c3f8cfda2e2e3879152e21748f1ba0db97cd4fc6b2cd1f620a887724cd00a2cd625062d60ae44e83664e7a3b1fcc0a4455d9688b7b952627abb31c042c78550d0fd7bce5fa00e2ce33117722122c818b2347d2eb50de5c2b58c00557ee53ef6f198f355a285a68439a19e380270c2bf9bffbcdf1fec9b23a43d5b73b85867c5db27df62db5048b56e74f3f2cc399f4cba35e87b211e7feca974756d55770be48050a674b1b3bd7f08a9bbe5213c1ed0f9e825e5abbd371dbdd762f4b4ab6eb4e6be3da136a06da61d825c2e5ed4604f1c4b2fb8b848665280a63faa64e8fa8d355bf15801d6227eb083bedf014cb472f5416badbac9069f59c0397bbc4f56a4a16219d5cd30686c003cb6ea1dbaef3cc3bd25721b37a100c7c4983d2afb74ae9b6c07f1e0a6a2b69db75571fd49d5b3a87a0ea3efe76fe176571e04d47c5e57bc50c742d369ba56d0e667b44196469e2c5608d3eba6efcaef5c47a23c0c6e4c1ba19c1a4a3b24892618ddcffe93977f00e233121cfd7d4f23d21afeb66f111327882c9467aa3d1562fd250db233f0c7ba0e59722881e3914b3e0d139e7adbd2cdcce8fb97b226ea2f690f0908496216cffa07cfde8fa28c15f80e4615b36a8786665bbaf3a53b3a689ae40af58169d8a0dbdd234f92b4d480b6fd3f1d54ac2e18b096efce36b195e61d14fb02a8fb5e554c333c60aeae90181aa842d175dc0ed6ce4a03f7dee435a0c8af2ffe08d3287859f9bc4a92d9ce395c6f4d6f432a0c6e8669afe8004e36b979e84015b2891a327e3abfc66f40834002310f41fe964b35746ca5c7e3a955369aafe296b56dd31f816be0152743a2f91b1906a4b91ec40b962a1284fa801eee99eae6cfa25c39138ce9b96c19b8d07a7c22e88c968e54110c6409df84abc0a36b99756c2e052e020dafe54a20f4413508fea487994fb144f980579d5c6bd2b1da8f25b271558cc1a0249e3101240f16c8dbced6ae2d340bf43ef1262a4cddfc3d28475fdf90bf44d84239e451abaa0b98212f8e6140862d2f6cf1b5b1b17d90e0b16a3d68d469e19ea425c511e2b8b77624cb9d3fda9dcafd2fd4bb678b8cab2e8ed6b5b4948fb9e0c8d5fc8e36dbe1a0768b6ee941f347d6d05fe6854ad5d36743ac6ff336e6165a76ad00bdb1df365b6c32c19c0fae09e178d3e48f06450e4012fcc18a84ca8a6bf9d1f3bb05be0e2bb22552804ed270863e851185b26376a0f8abb7d17c6a33fbffd255f53e3e7843de0b9e69dc4640a7d05e1b24015450299718f16512043c661c9469b1c6d119dd687e1a35bcdbe94c3f91ab8e4a50650c559e5214f3189563445b0d2d38d47d7b570ff1dc91b2e46015e3821ae043514ca01f133c3b415b7a81730529f296c21db5ddbd8debaa9bd3fa7b78d66bec358d5455a17d02f92a4fce411b635bbd5a774d1321b91303775732d15ead8b6c90faf424f3908c32664d8b333d5ebc540a0763f435a4ce46c14905ce2551698b1eadd5fab3625b3226c80cf34a69aa6b9f22af1829053b40cb3ab8a3d8da5259ba33d543f8b4dff4633746e80418fd34eb817bd3f998819d7a774c645a32ff9f669ed7a3b9a5638e04df2d78e8bdaa17d6c9b5102ba317217c0cc16446a84000f5ee36af3a3b9b8ba64b5c103fff92eac5bc847267e581b4dbff3c79afe5f940afb5a52f4163de8cb57ab85b950c7a4fc5b714dc38e9e18692bef5cf3a20b2201e8140f1655fc7fce50aaa16746e68462ecce82ef183b135d2a9176cd7ece96d9c6a0c7148169849a0e553ca23f1ebc17f78443d37ad9500e02c09bb2d9f0dd227a5e5a86c530fb3a86f755392deca0c2c35563641c522ac0498c759e6632f0b3a7f940a6a715e01e17bacec4d8fdbcd9435d504951a8f6e875704529e8a25cc7ef5ddadf3a140f6dd60cd3d916411cf6be783454f406d840a2d6028371868bced10b379001d784bbd537ddec79fae637fe5e23e496653430a601d5fe623b14765379169ca4f8c016bd52e234813f17f0d5d45a8f3ca379e534d2ae566b7a3b369df4a3263e6c37fea6f79ddad9ce2aebd9451a3f4ffacc510ab4eec10d971a7deeb2e6bd4dc94998e8600091894e5cc316c51d25ddac1424c825d5fd4f34e5df16ee196bd35f8a77d4c691f96419a93fef023c09d731f2190cab9164b94caf90416b7cc7a6e0d5ba076dfe2bb4253a97f0749cf0b9be86c5e65adc64d8bcb18371d00f6afdd9a0f6a8e488b125cf85a19842b2197976733ddd50257edfd24d5307e5cb0cfae0110992f4852b642a1bb4b29aaf56160cd8ec9ae39fe5245cb8a821dbe5b0cdf26ac793e00cfc0bec4a69980c96918ce23fd398e3dd92cc24e0b4a5a679b71b7595e4b6819d9a34865eb6742c52464a78afabca5017ed480cf1594617ae665b224114fac71975fdb8d0a5eb8b7f36df2cd2195c5255969f7919c304c55ba91ea28b1865fd47e07832b733b3fe8e7daf09db6f1b5b5ff338ae283e39849cfd15bcd8ec22fe9398211bb1f883da0793fdbf6c024389b739f191988c73d750e665616730113fa05cc8df24c0b4af3b91645ebea250024c1d2dae037cf99763728742b032d649fc1aee5168a8b02a0da1b0554ad72ca7182db9a2d1c7624ee8b5f19730d35b36a1f3615bccc00d8e59a8d3a2f261476eab9ec517e02fc274bf4c60a0a3e89e3b78c075e7af7bd85b1f2302e2022eaf6f7b290aa73e39e97846df40483168f7d17b86cfc8336522b89986d21626b905fd423f88c332a033348e74cd468ece49389670f30693933e95f9d620c98f3e601db73f5487041c9be736f48a261745e76734b46f44031ff15426000f19b170898740bb5d1dce75b47908aea317b86eb9fb917d31bc0b5f6d46fb7e84bffa86da21267614b8c7c82d26824bed351c1ecd207f76c98c1ed77ec83ba9e8a0d18094b1ddf130a7298e2253c9b52abf86c05311619890c2905a5aef5b8e84ef1693fd957a470c2bad4ee031759db13f22a2a0e29b583e09647337e7140ba7953d4c201f9ec00b9f816e307bec17cd33fa33040b2f560c5d13ad4a89b341446766a703e43c16aa9910eb77a441f637e3e31999254c8c891930351f3ea8af8b98f7c224ddd24a13568231cb431ca6fbc779f90f4623faac2cfd726df7d58a5730127f3962454394b2cd767f1d9806af1adb5e1995a96139083b295a057ee4309cfd3292a21ee30dfa380992bff775cba741a66ba2461f239f2f261d69dceffb1fa2d61f818cbd358f999dffa54e977bc1807a421c477c89ec278a540dcad00d3526bbe54725c88902d944bcac8f289acb7a46b2200d5ff820e20c7ae2cd59b845bc2c660799769cd77881a6a2474e33a4cb9d9779414a943583f04c7adbe70953d005e26bf2b74e57a2055754f6330cb0d94abd7720a395f46bcde85bf12ed942b715e2a1bc9d78d5d4cc4c1a5014dafa7546c26a5f18ee1e59462b50d02b6d9701a3ac1609e9b500879558a1837c9cc3a8fcf19becf466a51d9c81634d2dd8721dd4003b6e1007791500defb7843058a383f1b3c0616a66c4b3f7172fa97550019c72f554c682fbae26e4afd589fc35ffb60842cae3213aa35b6f13009d07033ed65f4710c2a73cf0cbcabea686c031643197e1583333e52f97497b108a59b8ffed77b94bcf7306a9789a13a7625091d1a4faf10bb94b36b1fa34b54958c1c8a8ba532e28b286baa03cb33362df42c9a7b0414fc66e5ed210ad9d7fb24f776bdb542f136859874353a19912769c9c0b1997812ad82a59cecd88058541fb6102ccdceb3382a7ac28bf44e5e4b3beb9151c8e05dda04672305633e9e8f6c903d86b7782b68782ed1e1a03906ff738592888fc10e0ebc0f55dc0cb87df083ebcaae4a046713684b098f9b4fdf3e7802ce5eb21903af6cf3bdf1b6fad78ef4e6f1e9e08e3841cce1b332a2bbefbc5b3b87d3b5e13f7d43018f43e693cf346fc6de0b7e36af2e0fde10fd8752e422dd91e056c2d24f45d2360e8fee81a034d66bda8443e6f091bfdec9ec4f222ffa5fd56d33e0617b97f5f2aa5f07af68efa25c1f149b0f76717aff30e3c2586851f7150b302928f7820dcc87b61d742f26cecdb3f30764972fb693e07cb25a95374f7b066e6d55dc7414d14d935830d3b1ac83fa81dba454280d553cb2f9ebd5b6084e9cb292c4be6053915ed18e4ef620df6458d97147c5de3868d40ecaef7fd2fc24d95dde9e0cb1b360acbec0ebf9771c6dbc1a3bf78f98d33cdf09c05af8368e7f55fd1e6b3d7af112f148e5a6bd035f6cca3daa95f8e3348a56d9fd608dc017aa992b52cf26da969afc9ce8b96dc1c45385165529d809660f4aba19c73d01e7f253a05f86e647deffbc6ef9159f5bb67cfb6cda132df135e19662240990e2633aa8e87e152123d7075ef8313c54d7154d65d31750683a067e0c9dad6ef89c57bcd9007734a007138230bd064475d2f7f8bb48466e003416475ea70855af41e460ca95f1637295fb4b2394082d39eb07044f8c6884a4b8802ecb80db704edd3ea482f3fdf62c01e67d69be2ae04012f2cf44525b3addd56f5bc4b58d01d90ae65c7b97b794d0c11eb342351b2bdd50f30c34861bdeab42c1c216015700f3dc6cb0ae87b0e1f0256a62d3b6ee7d9e6dfce4f30f7972f91de895bfbf0e9b8ed930199094c401cb431e0f0627087ba57d723a2555aec33aa71ceafe9af2910e7311a0be7101ca12971120e26454e89a3aa45702443c8c5b0f7471a1f6fdcc47487b114b7827fad9e830335d2e881385bdf560d12ef76d42477c329106797a51156811a2b7b9296b9dd83d3e762a94dd6283bee086a8cb42c3e3c9807855c82635a97b1085a923b10447eab64c39c198d7e7206e146fb5f9af3f27d60e2b2c10cf5c50c9da623f50ffa4bce0f42122fbf97616757c968eb013bed2dffcf004d60de471a4533fc72f61c211e358493d20048b5d73d706bc658602b1d6c9168c436ae163d080927ffe7123a2430ef9cde26684090e8affc77f82abafbe2573d71b92f6388158eba3aec7aafb9614fdc373e2e8d3b042c133337d9c3dc7600bf5fc69efe8df90b000e3e482312a4e58c5ed5de4eff863986c4594c409b4d663c3ce75c0952b796e80e7e27efa046f7a3593d46b6d203cb2a9efe2fc672f4172666c7057d5657cbc5e68f68766879daab3c5e9ea5f097335c09668068f145b993e26b62f0ce4e8cd94b04ad8abf6f62cee9f1f933afea13ff17c366bc8d35e940754891a37ac31e4b8cac646df5b7fb9dfae0945f7d19d382974cfb8d23f05faba8323b747db7de25c2d4ccb41d0e309d7c907fcbe0d8781c654b8547a134e76873ce8de90b595707117049b8aa6801cd3688ae748d67b08e3b6f7679ea7e4c811d002a5f2a38814de1048e7f9eaf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he4ee9112a39c6070bdb2eba22cf109f08210fefd42629460124efdcfb7fc431ce1f1b7e825a3e058f5c959a94312dec9bfee1d7367e8332cc7564b5236b6d05c2fa4d710b181f0207aeb471959538abbe1850d9912f8457569ef6123b3e3426a21813e6aa125966f34097fdc44cdf084dff788211ad69ffda617f8e09dcc6f3246f9b47175d01b4f4930c83f3f31664a453a9f0d06f2d4aabebaf603203ab4325226d5d74acb6cc4cc962a6486081fc3f93c8688bc0af487d63b1b0430de302dd85e610f61d5a334a464041a5d62039052a6d483d9fcd3d3af15fcb343e3c1b5b27cab020c9a7f14de78db869515986c6f3cee713e131e636276a01d0f235bb8b9bf8c69003abe8a3b85e4dba6fcb65120265b4af2afc8df1cf7c3c775b7719818bec0912a655105a4798a0ac585b13adc2eac0db3efd6c10a3b26c3af28687e8abddd4d4cf244c4e76fa1e2f4780676c0992b0b7330c49c6182fa59f1932361f7da6fc348641d038c928ac99a33d7d87947ea1f718557fcf3f4481b3c9cd82aac053ab889aed20578af6f68a848b0c30720ae6984665cc97418b6000abb9ae2dd95f3356828c91922dfd03a8f665f5e7777185fdfca0a6beffe43a7372dcac1d2a544d1da15d9ae6db5bf11032cdf50ad3145b26f1d8695acc22f03722a4c106f0a04c5492a9aa1241bf1864ecefbed1e85ff9addd7e71d4ce0377874f25f8852a350016d58a9cb6b73489068c847a0c96d73e478934ac883647a6be79c9278b06e27ddc71a325a50e622c6d153b879c12045c9562d576baf5daa110f089db4eb3933ec097284310f70a6c55b70ed3b8f02637cec62d8f3101616d87fc14f4b5ef47301fd9bcab78603c6f2dc78e15887ddad73bcb6aab3ddf9f6b50b3fb17a01114f3a3116771de6b591fb9f7dd5ebf0c97d46f8fdf3315eeb1d3d583c35af65952c0172fc46059764625b99616bb1259609b9ea549e187d3d0234012c16697a648bf7c3442d7a2ad85983a53bc1ee725e0c16bec65b7174f1e4491fbd03962cd534dfa8a4ba9c26fade0318a054408c4e15554202680d3e8324188465c1cbb31ef65c5a6c82311e04ff5eb9111bcfc45185b898c60c393f4d5f3e2989d7d7601f088cce8b14ad680c037a7cb30a0762b54ad85c827edcf4ec6644236781e25a7c9f2c50e82767ef4324c64ce1c0b3f7e26e4b5ce4a430a6a1c3005cfcb9309af7e5d2ab2745898da37677f896e10d7aaaf023720bc640b879701c55bc3dd840fdc4a32722fe8160586ffe7c5ea7f166c8c04a1130af44e2ba0e28e78067eddd0c4a5bb602bbcef2f84e7096a1194bcd7c1a23c49aa4fc2e5b61f2ebd9cb8651e640942810584f1f18674d1ee3a07f216ae0472aa9791995918167c36861e0043d026cdfc3efcd48b26e5f83bf86acc327842f6cbcc062a85d6d76e04682c0b77ec359f49ce850cdb4fde4b9f72f608c3aedaacb76dde0e873bd220a10d3a54e937b0cb70697d8061e2f8f1590605d324e2ef1347bdb3bae3f4c958cda33d087aa08883babc8618aca26da67169eedaf5061c1b721c09abe1ea6e16cd23eba90931b745c2855da83baba474d82df57c5c45e4c74dc4500de17b6667b3806f03df5f35e8a3275322f1587e84740e383b9abe0a5d10640dc3f6d0820683c517862724fa872dce85e1ea970ae453d6fc5986c33a9507229d93116fd062663f982881b1619895ff7a81598b65736c17c31a1920c9402a9bf38be564a25c1fb822aa1a3e04fde479b861fe6b9eb7e219484f3ce0d97eb6c8d6b7134f5865725942eb0a5da300c0a400f80e7109e3d0c9ad73f1fb7954d91c9d890988f2d95333257e50ac3c2d2cdb92d63c4356b4fd560872ecddc35985873f967293699831b73ecf5e0c5a48fcf99a611bfa46f9fed2591ff9e94661ff921aad5bd7c51808277483020f40161618d4ce045b70405265dd561bf44897b1cbde7017d46985907ab7ed8f09a01a27e24ad2057ee402fe4ac9e0e843a12d27685692ab8a052bc5a8a868fa53922cc951d3ee071c4075edf6c25e083898012d1865607f9b27087fa5877423b739602afcbb2e792c96bd28544b97cd0a0ef757a7865a1a400f7c6606e8483591997bb5b33f8e54846fd291850ce755c9284ab80e704fa453d10e2a11fb2160a80c33d13927278dadd9d3660f9176e8b7be70c2338098ca3814a0e5f849c364e58e04df016de551c4ae02d16b5ecb728e5120586de4048aaea0a57fa635f41ff3272affca7c568f736c49be9e982f7ec66330eae318eb14d9d1d87ba81643666ce82dee09bf04bdc294b4fa5b69117f70cbb5a5b02de5d22477f6232c5793515ad0cd64fdcf866245d5e02bdb07b7ea8010a86664cdfe67b9b3bd1607014a324dbf49589f7f0d4e2d292ba5368b668aa329ec1af80c1ca2bb36166d64b6be8c31820b76e83d120f848896d8d3e6c750342b4bdf43a99c06bf689560d80f151050c2b994ee424dad9d388a0c0c2f8b4d013a768694a481f9b1fed2070a037a577e2aa015103166d6cfc155e878ea6ae3beb9432ac747747be07a03b499d810fc65f2f633a41bd1915779ac38d6179b2dbbeaf9621bf64d3fde47ad0c4ddd064d7691513ac8be020ab8c4ab2ab4b7d16f5dee556ece38164193875166b39839eb57faa496592808462ba9ea8bbbda260e771e060c399294590e654c4ad4059db76fa140b43693bc3532f82b121b4ee254ce7fcdcfa06398cb14f020a2364dbcaebdf623c29067a00a7aa49d6160661a8c408f1c55d2195dfd91308c678321c8380dc66e0913f609f294d529034be2b315894782be291df2cf29a06b6868571c7fad61515268343a860cbdfb5a344eb76d7774d8df226acd7389477cf3ee9a6a843a112092bf31f5d88293719bf82e9dc55d2f8ae51e66a41351cb861e8f8af7fdbb5886cb8d79e9a9104599480ceb9726e8b692151fc139df7018203520fb54694fe5d31eb88b6f78e684236dfdff77def8665ee0126d2a7c24a43453fe3539874e0ee4fd6fae3011ebba96f4267ca03c80cbe8a92f1bf281fd5dcd6256ef933ceae6337d3d547338f9f933b6174cfb8fb85e78f0e7d1338c13c3e9e21df7a4e0e2adcdb86295f1bd7e6cbc321c6944309ac62706ce8ff0272fbe758a3ceaf61dd9057c42909647f585d8f031517a3732c777f51f2d365adbbe375f0404a73fafec51bb2f2c8005270efbbdbe14e99f0e8c8188a504cce453d729cb2d36524af0e03628ebba527bb1d34c335ed863a86bc8c6128d79dffdd74848e41d27c0243f4a08d3508f427ae7bebb84504dbdc6d5351d73e84c6a13176129b6d07f9d7930a548ecc265d81c20a0d790d7d3d5bcc8e9656f4c3ddfbc7737910c9d502c73035d19bf77d65b836bdcec9e6e1bc697ebc5bcfb629aa77fa57d218aad9b29e63bdb3e3821b2233abb180c36e8a6185fff79dd272d351e45c854b9d5900c128be214a3e6110ba12f0843b5059562b00963f3c3009f5302d86244d2e2aae6035d7909f291c221a058c4b6295e9614ab0ce5a43c449eede5f70908dff17e4f38554b3ddb493b024fd337bad8ded84278217b6429b36b0943468771a68f847917ef86e8fa106b4458de71fc30ca31b4051e8d617e4a84eeecac762751a32a1e5bb8244f590bb2e0d7fb8b0d293b61dcd8e286a2f07a7403375c25e96141b8cfe547e5b95291b41455fc0bd555f2bb5b5bbe6b9f8d2d7bf2115fa192a6f483cda53c24e98bb5a9fe8ee8ab04b1a093df30de644dc4cb7917ce6e7fd5808ce81a341a0dcf90dc35b61741714f78ab87a2645c9341ca6307d85d2eff24c349ce21a6cedd5f578a2a3ebf6e17e8b4ac86d699aed1e43dc591491ab94e55402206e7930a13b604acb764f0144a3b0838c342365ae6c4e08a6a4da8fe64b1c638e3763e54208a65fd78359c3f0fda51c7ff6d1c51fca59abdbab670fc791d1ee192ff90ce04bb590ec365f5bce4456a0cc39987d7de4cc16df37e203b8be9c12e46b3268c8d95758bf74ca67446758b5ec8b9a63fec2a72a40461446ba8d4b76418bb1b9e0d9f3dc4b933e1a808e999778eeb65cc68d6f030a35b42f0e89ba8f1df74bb8224e10b9ddae2c3da7793d659c9022f594916eaea148465b4e0ed7160bb2f4498bab62ad6a72555e3ee703722714e8e9dac02787c922d015b6a2faa5d361cb7c86b300b66d0e0c03989f6294ade7c262fbaa1740de5e15730e184857b416430b4e504c5a17677a289fdba32aae95487a8d5d7f0a2e0acbd0f0de133f44f5c286f45f61eefb30ace5b8551140810b5341c4b7e9ce7c9db20b7d6bd83a48f1b9da9481875fd5a0f4be89257d3a4667ed4b2069174efe0c53e41a764834775b32ad0bacf46e1d93a3da72bdf4a02370a672dab66c137ffbbc17d343ad7e59f4730dc4e69e0300eff51430599d2810f773c360abd1514955ce0c4df66873b48b7339b45c08c01a171442387f2c8d126011e31ee4e92b7c43fc13c5181f71f3bff951aa21265d6c3baa3df9a267b41e77ec0aa0eb1c0d8d0d532a1d915afd13a3a3cc487552fbd074a1e4ca9aed18fd1bdb209f7f56575c5bc1310dd0a96d87a83e74ca604f1e8a1d1034878f253ed353359581b2409410a098c58668ce258010a4d7e23f7f6bf5f53d5a37928777a24802c48f9e5cbe55166d3dce6328010a2c80e0ee89a8e34ddb97818b1c10f7e6bc96bfd5c6e3a45f201d766f2d5f3b7e2b0c568bcbb147034cc3c882dd0d70fef21079fa8fceda4e14e9847fde9a97b199cf43ea84870707ec2f93f339481d956bf81fca2c6c34a5a4878397abcb5dfbc386e7c334eb63c736a01ba98f90af39ed96c08ce112cc1f55268aa667b02b7af44248bfbecddaa77d35bdb756f32f5ff0dce7a0afacd17665ed3e4a593f6fee601a5522dee86c4e7ee058d86b046ecde64bc31d67cb428fa1936ee26a1306197da90cdd3bfbedd3a741f5096a6bbd006641e42cfa6ff48dff75e3ec696f0a2216f61d09096a717a4bca949ce784252e5ca857eba32f3c9822bc35b92fc325b35d0a5f08729ed73ddbfae82ade3493974da1d8e4dd76d7587860474bed53e873b6e2cad6c24de0c2fe94df72b92e20a59113cce6184dfff3bd0c118e7de75a5c34c7c678caca878f4af3f55c6a2b459eac619f478aac37c5820f642d64524d7baa2d224aca4f849663e01ec7e31301a5fe4f58d3e64a90bf10cfda25961a81b0c4589cc703aa909b959923b2b359db1e5342cd645a0ad48ee0fbe741c4b984648cab4a55b18edaea00691319bafc41e4119e3f0b500894b2a23658fa316b301e3476820c746127793431a34516a7e3268b4b70a9dd8e30a87e11e749ca3e2b23f9aa5596511e7a900fec7e5a64ec19a648b61169c1ea6fbc88b8d920e3ba4ca7362f2b40f0b1ede5226e7a0e7d667d6cbb426bb91b6527864e9b84eaf8ca33fc2834482920faa512850dbefcdc8a28b32917352c027e111293ce380d2895ae57e5401221b9b3960859993b9774bcb5808fa9bacb14b14c27fcb74cee7442f1a5e6b8c627133be74900e3765e81ee9aac1abfeb7bc9512fa54ef24c20119172ac23eaa29b7a92061755064e796bdce123c3ffa33363540316b9fe4fd1e1768cbdf2a5ceb937b54332e1ae1cf36bd1d00bd056027ff559bf7cac2d43f4e59653c627ad457520fa7a38c968c43f9e8f923c18abced1d2ba1a70914fde550e0c255112e689c4b1f384b72485a6cdccfefd34d868a9faf35e77c90e320aa7e306a74decd730;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h31c22d20bd07dbb499722ee2e60a1fddbbfcbd5cbf5b44cd03a3b954e7b9a8294412d8bb5f0f343d19d1cb30d7682acbafcc24f9d55d783ccf7b103509c1b855fa33ab7a14cc787bbb96054449202138b3f03b0a686c5aa5067eb688228e652f520117a9f6a207c83181c213c66cde7902029b5c6b295b1815bab25e3c9ed07dc5cf0bcd5d65c2e85bbc9fa1d5227f2fdf54c4a48b78c2584874cba9fd24861db66a7a607e5cc54704c4dcd1ba1180428e058fcd9dcdc8b493e09cef04330d95c2955cccb0db298a33f346a737ba5f5ab231263495ad7261a2150e5336589384b7e607bf8993ede1ae94ce3eb1b6152e8258520047667d33c39ac998ec9f00ed55d3abdef5445c7f32a315efe2fe983b3e1b85d56e2f8fc7a0114ab8707590a2a3fc600d08537594003780c4ad10478de23011c8c0684d56f1e7cd798252adf9ef1e6d6a39f773af5f13bf28638ff6c8af26ec644d15d213433961e7711b67c3b861c261aff94a903356f77a251502b359c759b22620e1eccdb2fbe46b05258fc821d978f85645e544f20c9638ddd51c3e4e7e9eea6bd32063f5128232d92b3f5a79c5011150158c805d3493c96eec9c7cf27246d95ba086ec75b29c83aea381211aecb5b23c42115a87ad73164407e08055dfd0f96b2fc2b598ba1e90a61a6728b15fef76112b1671f3f4be2250920e419aebafc9c7085cb0d1e5ab3edcfc6b9f75f9dded364d9d6cb90f00cccd2094bb15ceb88cf41448f45bf415421d3e2a9d0f3981d5f3745977aa82ec7e420afc7f7efd0c5a4956967999a8cc89ca2437c8d7334a8c1ba5aa8e568c29a534db21cd283cb092f4376ca950260918771f91985b5d6b4e195d5d477182be395b53e05d1c832791cbc5f3652d5c2f333f3ad61bf038e41d4b5d8921aa8dcfa122f48e9a867801e377f8c24a9269adf270cd52f7acac12d1dcec56afb3c54bbb9e55518d6291703e756a445b02814f3dd68d4f563c27922602d6b9233ee1b73f0bc8c123fd13094a43cf637ec1b83205f249e33b7162712337e244befeb633af33b7118361b322e55048a8ebfb4c246af200ea15ae30c40bbe2dfaadb118020ba948667d186edbd4e1383d2c1b1b53fe033468301bbebcb18aafe03ea47e8201805451ee06ee9da0543e6ffc19253763537604d7057ae08062787735fcd2bb0698a8c0dedef69e31eb0d066a2782cca7a5fc74b671cf8d75b0063c876d1ef86a34ccca5b82b4b33f5098743d8803404844889104c5d164422b8e7fb128feab1a435c71ece98ce496923eb6f83211f368f1cf48bb10f68b2ac7ab8b6a34b4f0b1db182ad011c5f052c2ac40ce6102d8c6a26d14455d8d3fde44c3b75d5968037c62a9f10dd4a17c5fe9324fd3f3399c34a87bcaa66a89cb6b5acfaf33922084941c77896205d94a5b5f4a6d8afe30d5e74453e1b26044ec369d1653170ca3e514cf0bf35bd8314daed783afdefb413e961305bdd90231ccf7f63f3ee107cb0f4cb6baa04e330b41522e81214de92f044c0fdec580b96f4119527c97c71ea3a32586f0107af9dfb4a351fe5aa9858922c9d14c245f7deb6fc8f3248c0e9e0043a6636011ef8c639c48fbf55ffe04f253294f17f31ed10a1127e4b093ecb50b12fc713209094d68d40ad6e7752f972ceca4bc638be2f478f4cd9de8d69780953f9a528923db0dcd28627cc1140673da4d6ef1d9ee6c1b5ab4df8a655409299b1eb1e7a0646b18f2c50cc65aae31e79da31f363dffa7eca7dbac8dda3981ab0faf050f866ff9f4254aa57c6d50f5a1ca0a7a7eec9fa33a3a5aafad82babd20b9f9e2de8e9824220e770ef9d1f664ef51c7c6b57d2fa9462e1a5e7b4d77edf5b9d2dfaa6ea60e9c8f7414bfc92ed1447e3b56cf02145a3253026ac5b1b91fabfcd7f43308f2d1f9e1ec7047e53ce8a4e382478a9660dcef3d983d71b13d3245e1f730dd99e6935f30c7437f2ffeeca98c963f7ca825ae33a16abda33997930283bc27ff729291f5667351fd24e89f129589d48059576072b534ae394c938dca2617e752f730d2141f6028626d4b2263ba4138851f592d1b67f197fbb4e792babb6ae125b7cbb50e89aa9acd64884005c0f93b4ac9d24faa39c03d58706ff4a631436d740e18631dda18f9424c1a11fa09f8cf9bb8cca35fd9ac75292acd9c65bedb35390158d3465a2e4dd1aae8e112623101ea10af78a783ec9162b79fc30d10961e8cbb7e8d5b249b87691906574537118b321420d2b41684e041d9e89cd83d27a8161b327805637a7a3200fe3464058cf5bcada2491e2e0434a0608cf028ce0078cd8902d74b9b087f9f26a2380a587d8edebab4f675b2a0385e202b79c2744b75595d6672981b6bbf832480d7506a722931bf238dc0c185803897439ca325a48bc1c8c1983b0e479ae9a07d3dba01f3b17249a415aeaf40fdec3a463ec27f239b53e4afdb5e0b52b3b0e495ad4ae5b5ac492fb2ac3b9244b64721044e8373a6ffceba20d9e678a931f27b63e97ca90c61dc715238b0dbab136ef32258d2aebcd4cc8476dd4318c6f9cbb270553382acfd36dc3832af56fcd1c8a40a49a732952b67e8712f4e46b214c1ee246311205d985492ae94fb7ed96afb564412cb2f2ba5af2cfa6992393aa1725b268f905fc92be2f860451e0b17c827cf8684032ce95ba49a1c103d402d2822510e4f22db642e9a174b43808670708a69dcfdb70b7a4a4ece7d084d533e718074e7d2916ca0ed74ff14ac679b8acb07d9e394fabbd6d3663c394d8ec9b0fea6601d706b3ca2ca2a1071c587420d5747603d4c9f8784a1f6429594ca1dafdb96bd49f5af24abcc97ac5f66d917d4cd43a411b022963250a88c979d3be152adb76a7744550daa65d42e4d298a72d3d7381bbdc7385e41ccbb22aa4b644fc315e13cb9acd70e1fb20c78bcca40743cb8debe36b850fd05c99fd149c8cd2e3b69dbabf780b3e39057fafa4453c6d18c2b45eb3199f1a9c6fd134a804e1efc25957baf5f093d1bb3f63f66c9d0122c43bd5480f4559eab382429e91dcf748450995f9943a5dee8ea3314f6c7137cde4817c1e966b296d0a75603c5293715bc6a44a62d936d574a80f5db327903f26846ea2d90ab2802f00a051eab595ebeb518750b9972dc7cc466b949812197372d4bb6e0d8961c7850e761f71c2f116109e1bc43599b4a896da79ef140d66c8c353b9590958fb1f3f0a121fb24afaf2f27cd0a4899b1d5c231c2bfcac78291321854a04558e0ebfa29dfd9727770669b51573c86ebc46398ae2e4efa2e1b3b72369d8a4596b478cf7f421bc34a3067cc7909ad68935fd03391fa108decb98555c07e84fea925bff1c58926897a2d72077962d2ca9132b0c2d8bedb365d8217c9e0453ceab3d91c45b90ddb108d5f2850594fb0f35966047735471ba68115eb013d6518fe5a54494a80795c6968503b6ec954ad5f7c9a73f804d67229dc75261a53ac612fff196db92f2e54ce6b4be8a1f28f1c15741ea0e737204805b7f1c6e57ffc4f6bff10f8208d48aa3b973391e712d1898a916e4330d5395582eeb5a17386486f4240395d11f9f5a78e3c0e7b245cdc1d5082dd2935f0adc64cecad4eb56cae6b4d75e802c26c110f25b0773304c50cdf91faaa4c347854381feddb1be1da2feb3156df65aa09691ea10cf1fcb0cee1072b98c369aff380bbcd5f1cb945c0c4c941436a83b359b00593eff4079fc5f3006026e534efe09da4a8455685433c6a802d990d355af3b4ef6a724fd462bfdadd6562709f7400b5553f277f77e44586bf362474a0ddb8d98d5f411550cff947e8fe3872288bc3ce8db4aff398c290562a90f5d1adc1d3d3de58dbfa5f901e7a4e0be0b98e6326e0484c2d7ef779601e425dea183bbc6b6711cdf69dc8631b9301f5fb677c2964d917b90a64e7c0a9b4dad4c6b04708046017a1c1458cdca0cbb00eba7cc52ea03940b315cdba0b5420fb492f343a93e3d4ff9bdf59fba4d2849aab95cc53939ff690db400e7db6325e50c6a8e3f34d55fbfb950663545510f56b92805604124ae987d323d80302f2de70a6027fab403dec6d1c6bd887bf8b8c2cb95b11b3d827a9a7c20c45c4b4e3a937a2def1009d00fc4d21dc60be2ab0a405dc4d65e84f7aae59cf3d69f4f743a4de1ec979a09f45935deb47e7bad6a3c37c7ed4acdedbb9673d9b9d428dbee4eafa28915f11731f038cfd4b4a78b057a9ae0696d38f5f4905134ac49a8b4bf2fc549706444b36d80a5f2105dc0191edde33182968fe25c30a4aa99067ecee2e3a616139f2b9403329bd59e381494278b7ddc52804088653b1df7d53a49ddaa27d2f76b0c02bb5bcd62b8b611623b5638998d7c36f8903889f4b919587584d0e9a55ec9cb9caa5c1da17547141b826f5fd9f5dc283594f12e5ed4b36dca9d901aca71ee8b5ab5077a17c0c72e94afa730ada384e017675a52adec32eeb405747cd226f5f6dc5f4f110c4129b9f3a2112faa63036e33374f498d5fd7a38b8ca4ba52723ed5dfc7e512042fadedb639b6b869036f152ddb2305557f219d7a7991153a18843e3c231074918b26ade3518d25675484e1fdc9c3efdffb3acc1b820a739b94a544e01a800bfe2a2205fd58079935b3f407e49e70323c2cde9b6752a62cf9ff320240edf7dfce8c9bbfab7a6e7d9b8a218b16d1387d131402ff751e5563f90b751445540db52c2a7b23a862400f6c232aabec70022647d0812c606e82a3bc46299602663f0a3ff48b8aceeb57f71ce239fbf0f504f45a122fae9ef73ba1aadb7963978c266211f83e624054d214bce534f9ab4954e3512eb71e64fe9104c32c50cf18ba719f176405c0ece81660f361e4cf3f366739357395f3cf9f5e80cbc8c9c7d21423e4ad80be533040a1fc8081788dbbefa50acb3f8d5b60ab69889aeb1c4f2853f378a23cef3ac9146f916b07b102549700d128f27d0fd7b9bb147e77ae68f70b87127006b357f39ec36697858e4c0b82702ab1ec071e96a06d9b2f3799f2a122ba761be0069eccf925f7b5cb97598fd570f8ce6787111903efab36d0ce0d389a3d20adc2f9879f7aa07a07c5d1681535a951172b53ea479dd17ae86bb3d415bcded0dd1b14a70b500a1727e99f9e402f72cf0f250a557f92586a93b11842b48f2f9c3a3baed1f85110f1d17bb63fe89ae43931cd2c1e9a2399e7d54b84d13f38f0c676c8d81131485ad5faa3b8cff824853423b91779a1bfa0f446864ed32cb21788befff9c755f132fe64fdc9401fd7ebd9667cb150ec564aff6ad795b7dead1e5c5df314427980983b3b07788e634d6133183487ebbce3ef8f230e3d32edf79022aa4552a6764759e78d5a92853a207cd9134b2e395bbb58451142613b6470df428a28acf63a670c081ff9a627d3b87b7cf1a213ea27bfd629d0a60c866d00db967e63da47fe84325fbf0ffcdac322c61357da9421c515f93182509475a1cfdc678eaa8c179c3f1ec9d574152cb36f73f0b803a1e08293abc527163e17983ecf9232e13bc4097eb85c485e645a9d8d82ebb961f0e57979b2a3bfd9646b6c0079736efad469457d00296df6f624e54456a0b0b8b678136d31ec13ec03bb918459b9bb37711915431d29533344f7a5f72fde49ba5340a2d815236132da5391ae8df8493e00dbe96cbc6fe8484ebfb7832ad8fb4f980dd8bf3caec8faf34741788179ecb4c0dc0bd02393ff07a86c27bf5254579d8839ee4c6ef702d2ee7d73740e94bc4e6af5097b0d15f33179ad1049ac1ec884b8d3a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hdfb6886d884d40d643fa3abd9649ff0625b4fb37c52fa743989317d57407b79f489682281e0f8353fb6a09a7e2ecb84940d74757f2e3119f3d5540f3058f20589857292190c8a7462341e47483c7fbc24c29eef53ac4eae6f2199c134fb75a46583800bb6adb4a17de7c4d0b369e70e32140118ebea29cfa468a90e5a2fb65c04ea36f61800156cbf981c485a719029450ec1a1e15d27f3576eb544f36a646d3ae203e731029214aedad64679c689d6d2206321b78e2e79d84b2c347bc69471e02ddd9df914f6462d3c1bd8065714477629497c5f3a3418b6002321df5a1b3999190745cac08425e0c1b54f36b471756cd0f0d4ccf9270b599e8bdea127138eb503c4cb56bab4ad184e339e63be50305b138a03c0db55d15aadbd6b5d148480bea4392222d38a5ada16e8c9e43055751f0d69e4a0edf5d4920fe553dd55b6ffa389945c37d1b8a836c180de287dddecc1aaa222cbf180e5667bed6c7273535b6686c2666ebd934f64ac79602fd35e1079fdc286309d363751fe1ba37df2c180aeb71723db0b426151342104afb7c32e698e6a438972592df8fe4bc7dd7cfcb309309ad01e395bd7b656a7e944e5d717e6d43fa330c17c080c255c8b879af0fc28fa74cb1547f701dfa39998289c6d20aad6766240466cb50b961cc82c5a6bf889849d6a0d2c6d544084a94f6090188e81361bc1ff4b85b20b531c807b86ae9bc39d4787ccceb01aa81e33e378fa63ab155cbf1066c20b2c8f3e8448950a86c744c2678ed52438e58b32ff5f2b282e5c22d3d0c86cce3844d25cf528027a415b28fd91c50731a399039369f4d0e7d6af4f129fdbabbc8b698cd1e47e0480de2483e00e2725e426353ffd07ad00f2934f195f6480e8d07f379c2ffbcc90ea95e5d0e2d9df65c26335b05b97ca67ca3464ce6103bbde5fbe3436952785ed99cd660e1216544ccc325e6d91641da8107aa2667c5cd5e44ffde90211fd3c922b5e488f4f76471e43547800d7532a230ebe987ddcef374243e7e41466dab817be24ce332b12037d7b73eb9a7340acf10283b5471428e7340b9c7abd5a4cad21f19347638cc95ca018a63cf05e4210678119d821199bed60c06aa8bf3efebf2fcaa87cdc7ecb5b6ba62dce478ff6a75e84ced9070da2f69c74937c0f29390922d3e21b0fa2e437105390da30bbe83edb0f6117ef93d4891e924bdd1feed1d08f2dc12cf626db75cd20561bfb665100b7699379d1ba6262f266cf6aa6c484f9e849482e93d12fc5c9bd1ad4559940ff0b1bd7f530c867737b76568f381903e74817afadfbcaf5d70d993981c23f855a64d77950e4888628f7e6960f379e6e83e18bb0be633220882d5e711e4f1b1fc66c7107a51d33525b8973e88dc7178a9acb048a52e3bed3347d58ced871bdcff7c5218dd0135a480d8c5db6c808383b39f79f1178bd23fd06d7efd0fe26a1f2581ade71be52a8687edda6fd1e7501ef715d0dca1f897245fd37b81a3fa93bca2bfff7f95aafc381fb94a7124400a45215326b3ae8a5c37c76ea93f41b1fa7850ef87911756b164645167b62b528e993eac52cf71026338cb7a96b40bb7cd191688a81e3270aea5aa79cf5b8a5d65f340a4f06a4ccee1a8f5e64bd6774107c0d4a38630bdcd74dbd90938a489a9e94924c531344102f8185165e649485f4ab79173ac9287e9f8fa92ad9915c7c2f225ca4764c3692c1812ce21f48bf638329684675cd801d96076278eae327e1abef0818cbe38c348af54c5622421f79f23359115281295ef0eb1f559bed5220c9f3688ac139a6a257e8528066fb215950cc863e159109437227d945f6d5daa6a852f7cb677234f417c6d254baba08447ab45821c9609878417cf0b5a20c7774208e8ecce0fff91ce729c2ba55289801df381af0bcafcabb68f44b629c4f4d8e2cc91594f7d402d1df6cec823aa69a8e0e1abc6c3e3f73bffc9d860d2d5bbe69ec1d069944cf9bb0e3e952d22cdfc8014677f6d8db7d87d235dc6272b50bcc27eb9906aec593c94030cecd9700695b210b14e8b0da156f6f91997c32dc224651cdbac04bcb65cf73de6961cef068582a19c40035f9c5712ea0491828d8b722bb1d5b42a91d08beb78ef820c5a92f75f8c0b38473477e1ed8373123d7823f1be6a29edcd2d124be284abefb378aa2e299cf5012608aa93effb41e23ccf1445593f9d7be5519d9997f1ace39a0ebd0ea6f3b946ea7c3b6199999135be223b59e6390c138508fab7a1b019448e17828237a6066ba6698c288aaf6701936b72179dcaa9981d8429bbb1133c3fc296afa30911a82cd838c9707889be26537af6b9453e8088d74997f1b2c350fea24491d1dd38a3814b3010cb2a57561672aa25d0857ee2bd621068c27099d693e12fbe926783ba7e2a368de86f72e715c80462e9551e488a087f8a20f3a95f46dd1cb91c1b149857a24e40a9b03dcc0065e0054106df474e178bcac902897e89484983f26d12b4ed1b7f12b6167509b3a7720f814cf0a20865600bbd850f2ff0404e890e183ad41d53efe1173a643d9d73cf6b8092ebe8cd3512b2c3d799a01ffe001a106a259379fcb45171f6ccde7290f57ee45bd0552b0e2e9a58307da560e6d5dae6417888d3d1b5a535799cf5fa3362fb323b6e4c5b2afaa026a880f5ec50b9ec3c8626a213b296a9ab5c65a6a42a0b78dceb774b7515c10efb450e2ea1b6606242cfe0caee48523f7d7838962a7ec3f6e301941e693599670fe53fb3c25bd098530012961cef5f205bdbde264659309891683d4a77ee60b5ed959baa23244e977605ad72dfa9107ebb4e917253da1180bcd5dcc1d702da7fd7d3db48d7a834a79da637a2977955706445e3580c8062307d6948afbb8f75f38ee7abc5427b31f4df023116de695d27e0d0b43e3792165854ff5dc2d704be1911670b3f024a92a09573d9befe59de9a07b87baf63cc5a69fd69ee7a8e0f61ff685676d21602e9fba2bd0367d6c0eb187962be1bc4a777707c36c4fc2796e77bda3fe787fa4a23c260872b4f226e4ea76fe3b38386550a5565c64b6ae973807279f5e8cbaae031dccd8af16572698ebadc4bcafa29e38eebd10b3c767c50148343c2795674676319419628060aebf7217fd8c57ddeac58ca8d547bc16cc3a7546ace166ef22f52d25a0304dc2141f1f07284f670f629a7ce6f4c8bb67a64afaca41db1ca754abc1a8fe9168b56446af2028b26a48e8a2b86c0d8352d335e7175b05137a03fc5efd4d6e85cbd6cf7892ef103a28ff93b05d236aecbf2a15fad1566968bf71e9c3fbe1954674310b22f0949814d8feb4bdf7548fb222ac675b402e72d260dddd63aa0704b34109743effd2c1c0e8be7d0575222cda79cabc378cf9423c1529cc2f9b57e12947181efbf5bc27c227d424817470a9cdabb8905f72c884772bc890122edee5d2ea0e98343010bc88423c041f757026ee927c205b25f82ea377be98f559bb780f7bd9335d5e71e1f6ec69c484c2cd5f3adc4625b97b3882e89b30052e722d63f676640730a4a2218bfb0105430169933b4513e5ad091d8524bfa504c7dadb1c8d6a4479668c3714c9be43e82d5146d0b7eae9d58449bfdedae508cd232e42c8965ee8aa7a1e834900ab69df5f01eda0654bbb76e2c8be0cd0e274cc0611138288a8a9145d2ea59d056847e3efecef10b880da49f1826bb2396cf0aa45ef5141ff6ed4feb527d3fc21a6232c3bb09d8e3bb6798ca2070228a86701307788fc82052953c44b7522397f0a3d8b9fb523c75b64d018db9494474f687da8805dab6692037002c03c5e0d648272664f5a25dc00b1ecfea4c90351c014e674a8121ebae074845023dd8f79398525a33be1c49dbdb0eb492f6a364b9bd84e509314a621537d096f972cec5084a1d539df0547fc4028f59df594778e2a101d474955aa0deaddb986d49d65e1142914152e697147267d32299077e3fcc0910f90213a5f1be8b0ed42aa34775c1dce34f051cbbd0760ba9f742ba6f38adf15ec6f4486f6b034fbef86669d7c9474f33fa0333b095f9c8ac69c4ac8236443b766cabf95a6e1d470f51034f0870489efb2005d69d66ee0f4aa9d7248e4756080527a4a6327167f5ceb3b296daede10c6f4692cc4269382c11f8216859132b67cc1928f2f51cf3e191bf004f937aea3fd9e8104944871372f791f66723aa3c18ca6ae6aab0e6b6908218ad058ce271d69192a47644de9d7743ece481f8c7c81b4614de900046e93e3c8f07903c21986bd6c1bab52a5e3c89d1d98af76ad938a74fec2c7a0f1fb21e0abd4544e0a202fd80d2dcd85957d432ef1f387d6727b768ed5a6ebbbe15f65fa7d3b4c996a9d1ed46b19e0c79c493dc93df7e952e0a3911297a5ba0ea960c5399824c28e65cad4ec85e9ae09437dacff49a8b585899e1719958569c64cab8fe1c88b9e7257dc603ffce6264c9d75f806029194dd0aa0a22113524be7f9b51875bf2e5abd5b6108810fee2ed0c84712222592e294613995633e8a5240cb5d24de2294734fa77d97aa4466cac62f8296b8b562917574ff0ddc1c4fc3f71bf5a58cf91120fe42e2bb2ee1761eb849b3cdbebd799a78f90b34ec0c9d825802aea72c76259b9abcc70534cce68b0a0a13cf5946474967c7e2d8615d5581c4d128a982a602837f49b835bb0c5ee0e4ecfc0f80f409d0a64c7cb6a6f5945dfb8372a96187988bac39bbfbef17e0c2bb9614af1b36e24a3bfaaad468bba81bd2c0d0f95826dd5bb80414cdd2c78028a688fd5da0a57a8dd45e74a8a3831793e11c0de5fcc3812b59611807bfe79b045ad079cb18c2f2e4fe69430a1420293a2401ff0f741c8fa0f8c31ce934d639211a7a4cb77546920091013d5a0619a4c64de0f14d34f9d6d873f2bd432c5d2824413064ef6b4f821e305a9c69edbf4a162e16d09deb0a6c90cb53f3a4d77dbe70b891821587250e0a8a0a2ecb0fa09db3894f60969606565b56a2249e84ea00803b568d4615a463b3ea4dda893b392af00df876e7338af4828c3ceb0cf77ca7747f293ead39eaf603be1a20142f7739c2a0e2cd51d68148bbeb5610714127acc700f17fc711ab3cc3d8f001ece4238f8ea7e54872656d4e77ec54a1c62c41d3c52c5622665fe323d7156339f1f3fca37bf643599a9a3b13278d1a10e09c2e8048c7cd51df0285d35d95bc3ecc2e3cfdf6d158c4d6ff793cc7b4418436b8cdde76066ea52712e195b828fc418e8b7f26045e769e469ba5bd1156e5ea412a66a9e8d64a2292e52c21523b26b5db6ce035d7803193cc01ca4d819eee1642cd0a9e86fbd24298ebbf3e04c7a1b02a052bb4bd59c5b7db296c142c1b8c43b62d476928832eef523bf98c58c77bc61e9f6f8863f0ff26d44fa9467519268cd421541e8f882c0936feb62585b65628d9b2bb88ab7f0679eef45e6ea1aefe11db9470dc83f63d0aada1b3a5dab2e9abd4b33fc3c9a6d295e80c8b5464065fd3c13db6c5a7a2c850b33bdff4fa82ac325914d2bd4eb6750b6efd975e2eef3ca90707dacd939f04dc853b91d2f9bbaedaf0060bd3f8ea7e5e2b637dd672439438cfe7418a72400265976f024055b7eae98b5cbea7ba60aa198e915d2ecbc03704d54c85b3f708036d3e2eee06333767facddfd0c15afddd02722a5289604f9eb6eb1eb14fafa4802b094aa6938d6035863dd999ca2478d4161815d7f1ce48cc1e1f0dd7acece69cb20ca67800cbf21313cf32c9b30111c752ce5a0ca7abd7e3b2f07cb5cb4d523b5b1510d59ebd9cafaa44f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8acddd0f422f929ed6bfec1a33826910185a97f5a18abb13b4a0151c8bf4765dc80a726785751f54cdaa1c0eaf8b833adc5382bb5494d4f7c35412e9e2242207678ba350684aefb564c9096f1e08f68ba4d3b54fc4951991fb67f5d2f5a89c296ea9e70ae461fe8ee9e69bd4784663480d3cba741d63451b2435aebfdaf6e53c8b570895bbf3e9920ee10b69ab86db732fa0d189befa5bf1e1945a531c4cccb34ac71ae6ae456c3363f090609c0bca07f3612892328956654b7a121831ceced1384d19a5d490bbcd5be7a14f88cd101f137e60b4711c57ef3c543a8d8696749d84028690b2248f5e8f3586a45dc28786b26c0ed6b5db9b7ea4e99e51627a5c3385570dd73758d79e94b22b819eca3efa136069053c0937879639afc3e4ab065226ce05ff66d4ada0c2672895de664a25076b068a97e7ba710fc9791c68c40ea11b0d62d9a34fa07e89aae0081b5057e8d29b6b9d392a667a6ddf1e41307a011e46c54e2df848be0dd9e13c239eed70176d0a0ae541da6d2e82ef6403a75f21f6bd9b9dad9920c54ebb9daa41cf7566ed119b7b949586fd8592177d13125a39c6c7d6a927c5a22c55f6302833970ed26ba185836518f46445997a067de453731e832f0290096219d5be44d204079d054fa59f2355ea253f868c366ff6b6d3ca35ebd9506c79c0d96dfae7360f9ad8f848ec2cc8db210ccfb33c78e5b2a08782534ac8882c2e3e18da94d934ace75c33adb4e8c35ca92947d45bbec56a516da4575b44327505f5bb3b4b8a1cd4f81f43f40741cc31049985613b4b4c0f52ac9eb1e06e5e563044df5e5597cd6e975cb62cce7b0b422f6873bed30b668c8996ea25e400a772f138907224303dc428233cec6c6fe1df062b10adbb1f63f6202a2a89f12353a8bcf17d27cbbde8c5e5926918a0b963648400c007ae15dae64547e3c9f6ffb9c5fc7a4e15233a24db4baa27cc1d2a684284d7cba3d91282ee760da683a7a5e06324aa77705fd0d0138f8e169eb24f98c95b604adb9532b04bd827b4e22d339f84358f6236af1bec4b1d600bd48caa7a60a01a24b5606179f366763fdcd9154d46f4d0d8348bb35f199f71813e48a34b87f863c9ce8907707c573562ab41bf9ddf825036e6805f59cae1242a25e41daadeb733ebd52e115e933432f160b448fb44c685e6ac7514a00ba01839586656d6e47b29db4984381adaf619ed04d7879a1433691b6dfcceff1b37cd8fadb392da5f397ffa944632e4015baca965f67aca8d4e110840a748f9ef3ddcc27ba8efa28b16d2884f59a29863c7bcfaf69b9d7cf2a66fa9d67902f7e876be13afc7c2049d30a85e55d330d55002a8ba11d0e5755a0541e50ad9f6d478db24e01f14d939281baaf9692445f13b5bfde2392244d053d9fbf4a07f2d1192d83e8ea0382a5a75fc20fac251ac3da8ff9e8312aadc6ba0dfed92bd8b9c9f76f847c679664def5f97c25d7288385580012c7cd86afce7972ed871d72633f901600300c3dc9a89e5ede6e68acad8ea837f464fe50725f4694315f088390a0d24d652ce64cb943a0f9073b6458ebc1d75a5b3bef55de6079a051a349e440ecc06f117fd263d16240b91245946d73513756c9e22b18b11ef2f055e5fc8445051abf3976c870e2959bc2e554b775713568c49ec5bf9e092213de5582a7b95c4c6e55bfa6a083f019928a2c9bd1045c899db0c307406cf7f6c2c068e2bc9313fa8f897dfcf445958e8df363f3fb0cfefb5209332210f67e4670b1675b573a8315c9dd9646e3726eb66b20ddc5c45734baecda688e024c67dc2ba3162b05944b947f382866c0383545c43ed2c8677172f5ae182446d483960e4d62062d006088ec3ddb5a61a5b6c284423e810593f14b9fa0f37309c7b21f547edbbce974af1bbe3d68610b0e900cde214f51f4965db0bcefedb1a2e525089c29168354abe8d9aca28096d6384af286f1a5c9b9e0f88352bc808458996dc9b94ff884e4e66c9a7a31a34d6d641316cd52b95a8fee8bae260894e44479e82dfb14f07268db950441d34f208a53da0da3608fe401ffbf0ff6feccc775409f6d045670b2c91ea8f7af192bb620fb2e41edc3bf93b8ad92b4e46dc445d07c60e11a086bc85b8650861d1d345478c44e3e2596015263bff78eb363b9df58c3dcb50dbb466dee35c13df126e9eb4b8636ed01ce7ed32fbcd13b65e95d267fc3d36524950eeb3ce4cde0ed27a48ec1e061b9fbf1123464aa65d3c7eac42d967e0178df104d6adf6f84b72a4ee1205037bfdb3d11daada41fcc9a75de174f667a2e4a890a940efd017da4064530447d8263812d0b328d9dcbd2f7e4b89a682d16e8ca6d0c827ead1905de3fc5b3750e30051881d6796813fe39c59193c768169fea7e85e7f50d87b438dc9d001df05ed2a91f3652f1bfa1e42c2acafaa58900fb44dbb2bb314d26c579899dd778e3a57f0226beb5bba0a2920e5abe0bc292688817c8e1465b6125fac5e058b2b5762f7e38d5b8215b20b163612987ea6af46f52e1878ec551315cc51be88db96e0c61d1314f54070d63b4db3cf962b51a371aba3161b3a6ddb27acff372469af3d79c28e5b0cf938a74af73e58bf9ce40960367805380de3d0aa99a092a3763429590a9b55f841bf364c1f5f257237f084a23c770837d022489ab674c5fe3de73e545623b43bec24d3c4892b8c0176c47f09f728681c5ae5ac1b959d2e9d91ec692a674b81be3a31eb4152f91cd9a2efeb7300a9b7c0a57c7e0b5885aff676abf39d9d8dbb5443c47d35f9134ead2e8e992c9b2d5e4c34f1c73ecee1c775067cafffc7e5aa67d806e19430cab3b720a54215969c2041d66f2c4757e19c3ecfd2c568b9aa9df652e4824f66a94674b982e87c9027db39d20f0b95be1a7b3b3ba86738681837722bc36fb572996acc0c3a2c179edf732b991bde50dcbff832ddf504d90ec75b216efc68a7c2378fa301e91df376ecbccae54d6cd8e83b3156d9fb1b366056eb9eb0feb1ad91ff9714f99e18493da1324f9e5b15ccf32fff9c4bfebbd2e4f49748ebd2c58924efb79ebffad8f5dfae56ad31882665e7b82607aa0ea68f318d7d6ff294b5120fb16f2d3c071c820fde5e5a070d62135534bdbf9023f8deb36a6c2f6f8c4915d2c109dde0831c9894a0dd9c62133faf219e265c92fc46d1d8df160b1869555addd6c3b215af717df1c2a84ea463bd18662ef8ca920ff4cbc8ae45cce00eca22263ed381726422d1015ad7e365b44884a6f2246f96f8d07dd7812f22fb40fa3ed51d7f887c2d230f424308c67ba7b68def5803a9563f84eedc1cde607da5be368a739713397970e72cb9eb0c9566b245bc341dbe2443de11d6b93efe3464260c73cbcd9f826f7600da9eab771f98b68be342dfda2feafe225a967cf90c82a8ba16ede30eaa676bab32299aaee918dbdb5418fce916bf5eb78e10ef4809dd3c2f294aa4347c014a2329a2b3ea17b15b32a0f0c06c361972beb5d7d6d56c451ebd6973c59df65fbf12fa2551b743343c778e925b18d9a2ec9274d07fc88ea8de33be7e7f856d70350b139b0c6e75528f0921e756c1a42b1a456baa213338af022dee47684be004703aa447d6fb9fcc985a40381ebfd57b5ef0ff477566ec27e54f18ea3f8628c621b40b730b1b4c95648d517fa88e199686e98335ea6e6cb2b5f0d8150647ae235e7d9bcfceb991f9c0e4031e63250c703a98d2516b788882c7edb1c70d42dc8b212fdaf1b65f3e5563513a191ed25d55bc44dded2a08d4de3671c70bfd7e1fc47409878ed3dfbbf11a654554eaa4d1c4335e7a20863a5c1854dc55b76bedb381c43becfbba5e45b62a61d8d52b624fd6288d0586c266a4de28f84a4465f5604ab1b4352cf20a256db7e319f4aeb29f2dd045c43df05ae72efbd36cb5b3d77daca5e1111f3c16337e0817b359e3f943d42e2fd22c58af6d5c479e30ef4315d38b9d9a70276bfdb5a4a097111e9f1e889b5cb939cd6a8af526257dbaefaf26cd6a5714e8a07b5630e8f5e27e2bf65ca663cb32409d6ec7fe4b7440b67195730336a5645f98664ad5205beb9c5c354d60f5f3f790b8641574c229f781ec4c3423422232d4de71a3ebd26e747695a4e2312a3f3f2a3b977a968f94678cacf860c4ee1caa30d4cbc608b6923504e3cbee384109afe6b581e25c1375e90ef9d848608ca54f9dcaadba06e76b6702e7591103b33cd74f091c966677ec520c3426b0feae91952e237a352bc78558cef47cf65c2aada5b63ac42cc855a7b4e707f7ffe62c8b23c37f6567292885dbc75e1f431883346a4a6211500eeebf24172222feea92fb79700259a5ea9c1b2047710c314c65fcb4ea377ce1cbf470079c94bbc771f4865cc4d8e9f101b5c3225eb59f047b8ab3240fc1ece26b24c3f985cbfb904c514b41d88c9d4ac5c2dd774a99ccaf44b1a204a64e6f1313c3ac7d420a6f06d403b0f5ff32ec07d37a8b39ff98bdb8d7e4aba84056f020f1ea00d696c75a5f5de0c5b2be1ec05ad853cead43f1b1758ba4a2a7f4a287f54a7c75877f2413c38c217162fca6e749b897968605ad85c101d7b4968d3ecab8fd98ba003f91ff2dc70f60ba03122ef231247b4263bc70aa8628d0177df4ff628fec28d638a5f36da570ec592d3254c21a72d84d764389d9d12d3220b2092182567a621573ff9a39f2e7fec953e29753e75fecb6c5e6e6dc43b4109fc546243cb617201863fefa97ed67c9770053ac11b66d645017be7232d523b96f5dc0315ab156531194e5a9e1641f5b0e6033afa7fce8e7200a5a3e9d1cd736b251b330b3780cf825cce1047cc77359ba1bf736f060d0a413641ef67e1c1a773fb5c71e2668ac20c5e10eccb540631ed14dfb3b6a17ffc73efacfd7939f1069e1fae9eeb5ab67cae6f2c80039aab218c617ca1b6792a3c3963771c2d501e293f34cd68e866263e6d02c96622cef761eda6d9a0138056d160475e27be894989a12e5e5517bfe42756d165a5ff376658c23ba1e9dab1a188b3d3ffb903a8d4327ac2f20d9e1dadb7681ab855375a9652efa82ca21e6ffdd19073b41940411e33785638667d5c02be7c8d727402eae83429fb300f7ff1fef724d91ed690dd32923c7789c4625e815c464a584d60efce22d0ca92a34287c8b7724055fbadbabf286c235fadd7b0e38fc658c5e88038df69bdee3a6b3f900df0e5f9d11b634e3634fdda50729ceec482eb73ff696adc0e33dbe153e3bc3bd9776a68c6e7849f8502a39ba7b21f4590184b4c3232c9551826f1b80a3fae74af7f3fb81549a7741fa79006b6569b51edd39a1ef076ae2472b864b7c84e6145098503ed45fdf288b978b63c19a6f4b639cb766926c4cb084158c9abf01b3940fc4ab8f3185a8a143a4641cc84a1655c199c8daa30c4a33bca6c3d34683d50a4c74722d6969909805e8262aacfe8476e42bdfe06643f5ae1e2a016aed041b3aecc0f1fe5c1d706289ae9db88712c2d600ed9df22c4348105accdc4e741c56f636d5d075c34dad5361a3dd6083abbc0a18b87ad5cd21fd23836e8ad8a0085cf231b5f34f3ee4c2c65b274210f7f86364aed7aec0bc4f082dd1e9078dd83f849b8ad2528d442a7b5e3f8189b9273969dbcb539fb22aa01ed6532f6398efcd66568b76ce8fe532c3e17d08fc1c76306f061bd8e9aec4346e4e3c0a3c85d4097b6d6f13853bfb6c92e4102e1e5e866562384688b99ad5fde85105d9c10630ab784e3520c610e5ddff844b79a15b00ea5fb817336fbba33607b143882e2a8d3e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc19f92e5ac79384a5c5af5023b102c6e8abf12f47714221b73642672df00945620b57696e38ac0d299ac8222e6c91070b0d108c527680f9ca91755f7427efe08f0e4d19dfe720f52500a5c5cd09149f0727e486a21b36a41af949f7a3ec8e9276ed302ef749bb950522db05976c694730c446b69c3a62ea7cefeeaf2f9317f84c421567331d94839ed39365f0b78e4b3b11d54cea9f32c657e9ab045a0134d9af8e6bce4d0fb50d9b50563e88bc47b8ac3f830b1c08629f18214727536fda2b91956c14b3f5f71c6be4042970565225bc1bb2a1965b74581bbccbb10014acc11321f2bf7fac0f21f71adc0af2d3b06a05219da7bd03651916e29cc3d7c83437f1fc763fcebbe5ffcb764e6a5d3a3c639f32ccc427d515b5aefd1e79f0072db824f8c1d4f0f161ee75c8fd14e9e8f745063fa62ca48dbb804b6ae0b7f938d795677d917625091b4c6da65bef58bab1cd449cf87abcff2c86ff34934449ffa70a86f195955ee4fe75a4128c0798b79e77b65971f544c0fca543944677615009411ad38c1942e425b6725723ef9dbfcdebf331fc925d01278be1efebd09dc9efee948d2164203ec4563f972c31c30330711066f2ea5966361ec28800eee8ff8d3c3322bd6b2af93a11f2ea41dc763c62ce21a41219ca3949a8940c5c20a3b1210faa500dd5e4ee616c9c5a1d4c921c9cdd3b92557dd4944861f35106de864ba0fa04628ac1a860896587e76fedbd4bd8998e1149a2dea42898255e748496fcbf85756c376d256ede9a13f17ba9b952c6246e03be8d79abfd5c0b68acbc403d4d9b3bb71c54e148544c38dfe6eb96c4c12b613f0a355702f8fa5086ecb7269b85706db801d13f45361d067d073f16f4b6ab3e1be4f0a3f6983ddd9717f401ca0d0967d40402d61027fa5d84b1ffbe806fbc2892f1d5dc3205d6669353f50a633e128b7b0aae2e783bdb1b75c347ea02805fe7cf768c1443c23c503b0f8b9e4f763bc78a01d0dfe2c953bac9d7f40574135dd01d4232314e753c16a11c73de2ff5d0b5050a768ba7bc24846ba1727272beef0a167f599f824f5f507f3a60d2c46d4c949a92150b6a81ddd97bfa22115f5bfad0fdfbdc7d19bd9c3c21f027a02588ee010c588b74b809c8c1987baa32e536211d7f2206e75ad32ce76bcb61280229abf91f4134f7ce5c5b046e125c9de1ea56e749e7e7295ed29b517dd720e0e811b084d1855e8dd3cd289c04d31a51e5a30bf1713500a4e3105d404c5674f73d076e731aeb99ef9057eb2ba1ec1f5d249ce0cf158aeb0502e0c748d8d8b1d8a9ea6ff7f76ce284bab34dbb28863f83df43089aefdc109d7669a1a60f6f0958bb1a69c6076a10362d4090379e0a295e78537164b5f74fa65089f531331f12b5b9eef7bdad196c1797d9ed8f006413a9bdb626ebc2bf0a670619bce87f0642bdd0dbe02b3d69cc01f89882dc00176febe02abecba72f41d9009364391ac1cca6197d3adeb0e2f7b7f830e4604308caee00986cfff6429d95428d203f81d49758cb0ad1a4ff2fdbbe8f95080ad0862150abab4e00916368998250cc977e56bd98d1952250252b3d9ff57d3c73060bdbea112525b1f873055ce0792a18239f9884d6d687b9102a7181d40f232ec7fe0e4f39f76006d9a3b83a0539ce90029383dda3a49ead26ae841771f620969fb74ad42a5a081cb4c40d5827b1cb6095ec9eecba5765904a717be5740df9d8dd30746cdbe4c3286cc19be77ff40f192a68ccbd864fd0283b144fdc184bed694cee2125a974f36e25fdef59609440d706e78a2e701366522c152479171ebe6b6be4b456488dc96cbc789dfff76fe34de291fa53ed54330ce2af82405d9509bfa7286970480a27df11145cd85c127c05f4c03d21ff18f343ef0055b332cd8e135bda0839afdcabca6801104c8a8bf6699b1adad786e165a6fa2b8a22d2a863067d2143707e96bbdd25d1a3041ede4a8035a511c4c8192cb7d0849961bbd1686d1c900047e24d560aa7ca42503875ab4795b2b650e8f6af95732e0483a6d896a408e723cf7f692db79954579c404ba959812409afc27022224a160d15571248911cffe6b1f933176bbf3d3a8f7c03c82a988fc6b4af62c1641802b3fd3113fb673e2892ea227bca224983c98a1bc801fd4d984aff669166a666b70d0e28caa1dc701a58a6e31ecc527a4103b4b7ff34dc261bc6920821afc7c0f6ec94fc8f902c816ad9d1fd1c73866f8c3f6a36d795d718d6d5b5e78d62f60b361a419c7d37f056ae578034c204863e44626cbe96d54a2a870c66270736b975ec2144230577f58e9060989aaf580bd07c28e91d70a5ebaa83f6a3d1a6d0092e63d2f72f0ec4ad2a1b5c010a87f2c1ee74251e0add81298a04794349cbd576716512985df10baaa09b0c59ba4ffdd9c40be60c8675a2049dc4c8a8b37a5a7849b8f269856dc1f24ae3181adecacfcaeacd3a3a7fb05a2474694f23a01b3e7b3c6f519adfc0f492687579fbe45f962f43758b9580f2e68bcdccfc7b2f6cd13d0dfa0ef21ffdc7e439d74dffac24d9592f6c3389e3e6c74864730ac334663c636474166177d0dd8c368c6708705e93062ffd0572b3a06d9d6f5eb58352217da9be1f357134bf9b5a1eb2db831d2b158871a07103b27ac25f671082aa0a2796542427aeda8a60785af6e9fdc03518f11df797b59fe81807b0b3aabf81fbd09da383fc2a55130e413198d1dacb9c73089e38e1441735391c788e43a9dac68ffe19c2edde3d032d54dff4974eed5c684c83c6b5fe3d7e8799e0caa8533a9e9489a072b1dca6bd77dc417acc1f8ed26cad3291fd10a2e6fd1e9e9c39d7b63410808f3ef485c8d53e7dab8ebc2d3e148b12e88ccd1c877ae07db937571529868734a198ba929116ac20133de03d1a51e3bba95c1985bfa1226a555f37a5b3021f951e77abec73a1614ea15e7e177b0e0f494655c1124837cb528e62b671ed2886d1b8f226d213bdc0d2b5ede3d217cd00fe34c3f274bbb88184011ecbece61759bb5b1592db10f2fa8297d4ddbf57c89cfbc4f5c768485a5ddf4e0daafeea333193e5b98478598e7f18d6868645917a01672994e4d26d07a3f8ddbfb5ca18f311c9caa363a009ebce64f02e7f09fbac9b49fdc93cbf3e062635eb3945e3849938e9b72ce24ec2b58208c73ff46c692815c069e1839cd9ecd542dde6d2ca9bcbc9a3cac12db27f7dc57ade140b212a0202e8ac2439d3429d039aac4bccd7072f66b6f06e175759cd9d51bb285d670596963a399e4922f59165c52b953a5e7bfb780829c32248b78400971cbe9534be88af5a863f57110b4202fb88f923666be644d826445786c2240a8e39558ce778db15dc7fc8a73a63060d1d16c6ef9b39092bcbf40069ce6dc76f7e594f07c99cc990fffbbb6f43af71e0ae0bef22b4ad3efa0f8b414da70eacb6313a4426eedb8090d335e513440c1ab7cb2cf85b47842be278ec133337574f1e6a7b240ec1c8b568650146a86f4c8326c1512a433a71547ce7a7211ade06ba0662da67becb7fa42b604573f62180394a3501d7916c652bb3ea2cc1bf719fadaa3a220968363fc961cb516e2401b9af2fab4ea958742c4c64705d68cfbe487df7669c28393c615ded5b65499c917bcba5f9f64c3846cf796c563ec1e16b36aa85ca28ae92b90c1d8289627eccd1ed65f7980dbd1698b3ca55a866b5ded4b6634772d4d4605dad142f040382a08c97587a0eb657bf1a722fa609e616bfd0689bcf23c20bdbeaf5a59f3e5294ff6fc67a42375da0f2b21394fdfe0e9a995c360bbb7325c569f513f93aadfecd8a6e63ec68dd2f417c45dd4d064eabac620150b3019042eea29798051122fe6aa573145620573ed5af78cbdca98274b0e6b2f9ddad9f5c8f026e37ae56863c950316c152d6301a24ce89be577c4d40cc0fd784dfe4567991a3f40036d9ec000ea3b63e3829bc1ad0edbcc69c1dbf114823c6c4a94b9720d4377e89727b8dde466e70e085faf5569ebc9947bab4bf9a779141a556fcea2d1f40dd7e79bd95cbb8d8922d793615f7897ca53b45a194b6ab7941f08c6c53bef9233a8d4f0a76096753bb5dca13a9e59cfd7ea5b1ff310945eccb484e0454a65015cea5e0baa6e77f093da69495b1b650ef3e104b1b5c8683ec6a2d50b21062e99a6838de6b4e3a7994a38880a5d80830c7eb832fc8a1e177362e03f6d3c2c1ffdc4a812006c6d2770757a42fab034ab2df4a926477d70e8c828730da6855c939db7eff382fb1611e61b55c372a7cc3ac5b7c5612fc04257603ac70aebd6bc1d8e57c4791f3722052fa6e6dfd6c801ac18373bd7c18f7127cbc21f9c680e725191033c211f3843ca4871e2dad64a90e1eb33872067afa98d0fe8a4c0ee26439f9e3d851e6aafb0f85a5e9f051e779176e509c3a3242b33de5d1bea6fb7701b56c8bd5799c7d4f6e5ad02b06cc48ef8c9b5c70692230a1ff7997b464efc28e1f8424f09b0e7892249fba568fe44be2773dd42309a41b87e62cc787e4e244d1b94c55761cd2fe01af56a87be441d6f93e37db3c2f2c2679cc0d3c894cc0fa3546bda6e11cacdcf3ece9bfd723877408106ca0cd217e9ce914434e1b2cf828f0e0310bd0fd9926a6580e3a32b87901784a176b13f6473636b3d88395a925bf660586600e9ec97e6d546bd3364c6b1c2d12d62f571c82601700f8524f0b6f8b4e4e14dbe55adcec604def6dc634e8cffbc97fd5941b927d7f37ae20f4fae9f628f5972837c741876d5712afa59139b9b99881095d3502a2ab9752642b6c0b970bda3bfdc283e998544bf2d6d4977aac78ae6794de845b623e47a419aa3710f30cab5141d74a0388bd4282296d07b571dd93510dfb284e9784dddb8392ffcede12afb4889506a8e1463e05aeb5c85b15a7b6e9df88275c39103e6fac2ad70e81ae9ed0e298df346e5f09217a96eff1ebf45f0e8f035116c73d21f14cb0ce09ea5ee156297db8b7e442bb3e3d42b796d4d9bf34aaea8bd75e65fcc1e6ab9c654130a8c6682b1f28956f0f9cb01e17ef19fa874a82860f5c738d836d87ec25b1f918d3562eed2737d2765221257cb8853edc9b4af9c3f9894e3c6d8fe60ed4eafd606055dade5eaee1ff26c658f5d736efbe04ff79a63740e7c5a7c9e4634688547958a1bca94c23f2376d562b29059b569ceafb577b88492daca353edbb44e98a67c29356f351ad10958a1f5ef6d09c573bb86d0df79f50d12d065076cd21501d3f25afd756f726469c1b7d4fd27d202b3016f3d5e27673c184359664282dd5d9bbd16f63138f6dd0297e01eb1df0affeda5ecf03a7127a9112336726c90857002ae52ea43fe8ce7514438c1cc79a385b07f6d64220cfb149ec31f0804a57e9d10bcba390d8ed284ef5efef429631b65c2fd4ecdc7d0a3e56ee9185e1047e1109532f36200289d486c2fbcde3e6872d2a710fd8fb865ffcadff01cac9c164a0b942a13a330d81cd6445e81573ae8b7e509376566d52da9d9a6be4cae83c74a0a0fc1a8b0f219aa663833edcf3945085414b18bb53b28605e660bb7ae8a414e459a5d0ab9d7e67100ed4eef88e423747df9444cb5b539618107562c0220a26cba058c7bb18c985edff43aef59317dff8f00123926cad4fad3d0ab4e38f2d72d593f35863759b661f40114d77369c570fe975c6b09284a79ad128e6d95133078b05e9a37483cf3c7257cbd1167ea0fd45ab143bd72b86e9479448098cd8d9d8489a320642a579d1b4ba4074fdb30b3bfc24d8b99a9d4c88468b8b0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8980be86b5ac3b03f96136ec3eb58ca18e408edb72a2ac6692125115f6c62efd33dbda4fa954848531fcbd41a216cfcece33e38aea65e49d17ecb33ad0b7aa2e0dba6523a5485727eefac559522ca782141b836c08dd4e9540199a4188fcb48419d3f9c465f8d8722bf0389ea5c6e4cd273ae982a2009fa06dc2f28dd65816043f97ab4df84bcc6bbc1cde954ccf6740ec04a9d537ce68a8b169db0e3aafad9871b4f032a2ed60eb2791da58825816ccde660dc9e9a5d72d9824463bbd1b686b7aa571536b54e52293b2ff7744b5c21cd44448c86f4163915a61ad0a4bc362aa04628192eb0a9619669c36a2f9abb12fd8baf50e1816153e4cb22cb7a8794719ab3589973efcce005daebffd0b537363dc7974460232cf54adc03f4416f4ecb604bcc0baf07476f5e47b3c9fba74dbeab48abbbdd43ea166e81d7387750e86e8967619e737bf2277db055ca5d367c22e1c47e1a20e3a3a311cdb12a36dbd4eb46433ff527eb4ab30f25efb48b34799f63a28fef568766c6faa95257ef7e16b8b40569e314230e8c5addff80e8c921ebcfa0734edba3dfcc4aa8cafb68d0af8ab5fdc9e04b2dd410af27d888bcb8aaa5939c78ba728b069c8b3c2fd0ca4587cb59b08e4338fa45da31c88cdc0cbedc80af78cbab4101d87b267ccb3fd70c57a23c9c7820adfb04aa23e48caf5f2e9385207c6e4824c2a785f7ff12774ec2905f39b1213afaa582f480c3a6cfec8103be483c7067391266d9105d9b15ec5e3449159a3540355682a3fd0e60aacbc5cff55e837ccbee44e5e04e835db89a1fe7738500c7f4de3d9a760251441b04999aec9f3957a8cadcc6a49c19dc29c111026f524a257c86f9e51f3d08d4ce243f683ee0434abb128b5abcc7f6a20a533e36dbf32f804a425585fa84514b7e36e3f41afdf6e8db166586623d1aa708ae74f6f0c09a5cc76f262f3fae6899ce2aa18826fd46b992050618cfcea4ac0433adf4db9342bb63d8de5388ea3ac5cea1553dd31d6b7df9e5a1be70204d6706b95e9ee591cab9daf83e6ecf0899cf0da60fb5e71dcc364a21b6cd8a2d9083f7740511b2e199a5322b793a672d9238d47445c5e063999d63654ce18fdd9fc4bc8cf38f48fbc020931a84d86fedb3c0ccd5503262ab269ff1497d9fc6be18f63fc3ffe85f4ee3f73144dbf7dd5fcdb87021b1223fdc88f2eb0f0760c8247036b7196cdcbd325c66b560b143ec2ebe2e1da44025f33d503f7c9d60dfba76ca6531b49be420d887a7133eaf9ec0653788c5fb9fa378a51f220392e95896ec8ac413bee477d12cc0cc4581a54cc4ae6b3f22f8de95bdfbc48287b4796d87cc4874bc4949e1ef14358138cff4c512c30cad9f4be5af4a0121a886ebc92a55a63b3a0a60c8d296a66a90e5de3d9699ae1c019872a7a6a66a8e710d71f9403ab976e4211a582c082f22c49065445d41c285e0c5c5c5f1c8cfdf40d260248bac5707c66307f0a0ec9f311946049159d1e28ab58f1026cf73b901343470b403b4be35a1b446b36674e86f30932bab2c5703ea3eb790073973ca1908c37b49614cc14eb92f2d29bb73548d99d1b67fa08bddf86e3dd811122c57d71bbf235c02d1408f7148a87c01ff288ad8fe5cf880dce51831f17ba7d1df90b3b881decb59e2eb362bbb9db938c48025e774842346210fb12d1d47c7c515df94c71c378a925274f0ac0e2b86c46678b217de168f79f781a011236a453da2e28429ff11811d5710989577356b7eb205a4f864cd2521e54f3725ffc932c32472b97a40b9208068c9dcf4374166f91f963e8b4bbfbc21b57948f4926504f4335996fdc0b895ba4eb702156bbbe1744c314de1fcd5d6d2cd62374eb3f1ec277456f9b656668607a6e3a1adec6b2d653d3bf0a0583e7c25f75c6872f7e1f5b1e1a7ada731d7ac10049c4dacf6c2ae8281bbcbb2f6f263ad7557bf368bd600ce5b4523da186fd5bc91f624556a663ae1e7d85b5ea8ec2fef2ef57bd8e2d08b5906ac175ca2610e80e7c53190b17792e4311fafe6499244626c6369e82ab25f554cbd9c64e37dc87d05fd5a13ee815e404b41ef31c5b9290430a514eb6f9697c4cda01f05f4e8b721538d42d4182a5e31a0bb98d6ff233a429505eff1772f3696d36f83a22b9cd639e8d80d5b8b88f2c3f6e5c8e7ef755ba64d3475445449c33fc1de7e52e43f077b26d78697e7d9245b6dba778e12c5ef0ef9eda95959f9e2ed19d69e8c3a788a945a56faf16b84b987ac5373dcc9ba4f0c524086f120f4493e2d8ac02cefa301de97b2022a3e2bdc4d4c368a3089c8b3b2370a3e4c4d03d8e7cb84a12245fd2679a98faf395ff9e8e354eca19798a3b901b44241ebd58de2e5b66faa1cf4c0795bcd8e0b59e87b3b4479f41f1f62edf2b3852e7e9d6ac4654cc9cc4aaefec66a439d6bbfbb3da60e997edb97fd9dce25add44429d718de388a054c503fce446df9666529569b553395093959140a93c944cb7cef52c154f1ed2440f1331bfd514c42a7dde9874bc26c48101c3154712f377f5a41edee38fbc24b0ce2a5d044813f7a683366ff44c934537c5e22ec52fece7aadd3dc8181eabd45c4c00d49bc65353283cc949fdae34b6a66a03dce11b120d36f2c528b6628a0c94249a7db77d9ae32c181a8b9b64d393c64f368e363b0605c6114b911c68ee6dcb416ec1650e1318dd2ee3d8010f647f8cdc34ad41181a6187aaf2f015ebe311b6c654df07af51abe426d54ee8fb268501f5cd7bd855a7da7e96ddcf54514bec1bd0f976385cff97c5f07b4e157b74c26101286004c4831bf0887186c158010d65d93f220aaf2bb3832eed8e470659e1bd5634f57fa2308fa1d86d08893560a56c44d7537d06f2a731ea56b0af4f3838794cae2ffbf79c9f51669bf6cb507eeb4d277a2be29dfe4a3838fe452d9dd2ca6e2c67680e746b5a3268792bb31ef37dbaeaf7e6f4f78c9cf1a46f893c8f82306ca537a9f15f3a56afe9482777393303b1668ee860b4eb65bdd808c4723214d2d3cfa8450ff1e558422a2f102693c94ca5328bd089afbcfebab746ddccbbb5aa8c969ddc33016274bf82fbeba8afb8793dac1dbf352e64abdffd092825be11d727d33c6bd2b159c5535820b66eecaaab3f8b3dce5339e06f131d827064e1b1defa512ee6174a2d6c92811c7f671396878ebc7d1ab9b9fa6b32ab48eb8f2aeea498f8270d3d4895bf04b5554b41793be2c97022828b3fab7298d071299998b5361e77661523277f31ac8c8bfceb2d3036003d1aa2d25ac5e3c1efbeeb74a6ee6c5ec3853e4b9bed224ab266d5c5034e89bba729709ce398620c486304c6f070cc15136c79fcfcdeddb93cc095f27e9e2cba2fe7c1b4bdbc3f0bb2e5325b8bad3d3eaad5ac2a48ca6d278eeda42aa053d4a878eaf9813a72c4316b0e09d2fa0f4f9894e49372527e0a7b62122800e175fec9a2ed690a50d921fac6ea5e11a2148bd9f2efdd4cef6dbaa9116e563383373b6a53d1234b4797434e7c282b71c95449628c40ce4acc27dc767df8845589945e6771d882dd09e736e51235fe92700d58ba08720bfcd936e40333399d13dc7b303f6071f8a0c65fbb6aeb6aec503a6b8f6cfceea0129c28d738a9ecff7cf07ca44a067866b598f858fa66e65cb370ec09394afa64697ea05b71427336f1ca7e8b42a6c5856a12c9c6c0faf42c0f0277edfb8f8ae2b5fccf8a2bf46e792289341d610975e2222b5671cbf025375852893bce864aec35bdb63b30105ce706e18187d539e74fed06949f6a4d0dac3a2c34432bc52f4510437ba63a24d39a543572d85af7eed8b1f4d73997a40a605cc2dedc33c976d3b7ee3cc44db3ebed9f09d3dab19e34487427b63902f190800538dd16ce683587c6654570e992153b29f9425e2af99cae7af1a7bb2814069237561759aa10df1555ed9ccefea5bdd5538a2bbccdb56ffb5aa7b692f53530e9e44d1fcd466ca0f548d689d601f0ef99f72849637d0b7c538d6ab6b5072b641c2fb04d1fb75cd4d0d36caee29ae501bb8137813fc9ce1857f321254723fffe39921e96d43353c5ead03dbb0774239c4d30095eea0358a0d5599aabc39a2f42f04799b8b5f044e7ed50203dc2cb6ebef1596b035fa0a3b49aa7da5ec2f744b2ffd45fdc7b1f7c7c595c96ae758eb2036d44ff08e5bcbd4dd8bb95affe53e1eecbddbc691f9171c94ffc3648414f88318f204a61b452d5baa590238446c33a93ff5322376e54edefe5b050d26dd94fd68e978a096e210609bf6df1421bbdf7fcca2642d3151d7c6d514eaeaa90ee814e3645c3cda48e840e28e3d9011095f7c9af284ded407f2db449b70ccf0f02ba9cfff89921b56f2afb437ade92b8b2300553eaaa9e3cbfb869c3ce256ed0e14a489f2fc43ea7af870063383a113292b7bff7d10f492e4528cdaba82443e9afd7e9e1e69f813432d9a79b666b24c25ec1a6d9b070fae52c24297c67ff8ff1fce515c8315c3f06bc9c0f47700fec67e87ed9c010ccaee93c188010a85cafcc50504cf88c67915874c7b6a49ee85d5845c8307618ca82d98e687c5e29e28e795ab239fe176a0463fed53fee24d3f41c56b12bb38017d45fa70ff1e60b98cd7b44656df1ac0a8e257569e436527150538b9f00e46fe476947e0dc72f342dacc691f06c49155b7f147ed681100e7c43aa0bb5275a8a66f310e694e01a17e40b445a42656a596e226014f73fa6f92f3bb91ac81d19979781c22921566cad37b7f3e5590ed7b133aadfe87c1f3a218c14aef33077c190908afec6f7221cb7e2d702e0e340dccb30e09a94c41e1af890a2b8b9b862eea320b668f6841b181ca4c8a3de55cd6035374c18c510d580574988634cc9a55f59fbfc782704053c4f5ccccc2bf51abb91ed882d56d1dc1a7de430f504e26bc5947a8b3ebfc9ca03440bc8ddae78c3b933e73bec2ab8e0732f7b26d5decf1e9ed0a108d6c48a88669c426284fc10125f0988904111bc732ee472382ded82245ccbde8f9c6a7bf63ed5be8e49f2e80279456e21177620f789846bf04a78d426bea68cad4ceedc04b2a1df2856fa0b979c4e4c7d807dbadb0780fc563fdf65fe81ef182db22ab063621d8caf945adef67e59010b87f1206fe2e10573e8dfb88e046f6a5d443d6ff033dc3f79902c30768c74a6cdcc3229e196507538174ea905bd4332752dbdbe04c13a326a929e7f244191dd9497dc098d440152569204d4476531946450b14ec478bda35021b6d2a87cbf9f99e01a4ce0ab8a67513293f155d415ebc62073fbeedbbfcf8ecd1aea61e63badfa7560d9651bec444ad0d2b99b839de5d756d0920f56a9b1b614f83eeb2d2bcbd92782478f02226983ef0c4f3fa58f798003ad747522beb3424350260477e223a04956ef64561fa960ccf96c417a8f7ae0057ec1bc35a8ec9ffc12dd00f4f046c27db3afd35afce61064f3b0ee94d0d6806dbe2c2cd3bbef95fd114c89e146be8c3cc42e7aa66a9a008a898c854a9f4fb1d5339dac38e3dfd658912f0a56fb91aaa2c449d2f3ac81e8763bb750044ac03fdc12bbdda1675f0b5e8fdb97ab263814b60962ac968b7ac1c62d0b60dc540213c8e2d8190ec0808b8f3fd9f045b210cf856f1f06fda57265f033a92ba18ee9a28aa0b338c958484be65397a5ba81c712421dc9f7fc52cedfd665ba6fb44bd624481a51651fd3621160ace72e892dd332dc9202d6dcbbc20e00ba0405a345b54f5af9958ba3582a029b302881677b0c17ac500ce42401c56ddd03564a9810c99279db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h26f10d9ab3adf5cac5678d238a67f904e55aea408aac9b61c069bce993b75891eef6b07ba74926575bece5215b9d5194725a491d3669dedb207545ec6aab2d560f97b6bcb12f32aee3fc1dd9edbb14cc359a5c3213ad61167ec5872242998ada6e6090dc76733415bb85e0e204b29d0191e94cb3142c742bf24b458c16a5839d9d63cc12c5516766506fad753372600b091ac7eb902e5f89454d7a543a4d42a97e5dbe88f5c64c484a02c571bdb70368b320088ec2743a0037144f77eb380326dbca32d645bfcb363e94ff0a410d7b7371346b4031239d2ec7ecff80dddcfc4a73e67875fa14999f4cfedae90f43b2d5170395cbdb21f242244e17c8be31830f489abb052f2322c3ff9beb26d56b1e6e901b36b069ccf42bbd8eb40db80c50220520fbacca5dc88dcd05c9b66f3c3dff8c7f82951abe2e67eabcdcf17ac0eb632350c6a9cf39ac033d642e63743dd62cdfd0262c4ae8be514b23d531562ead196e882793307b8e730b5d406cfeaa3a604f0490986d99af628d6256ecd521ad7a8b113712c194e1a50f112cc1276875f1cb8b96f7e356f705f8898068ba14a1f233d4ddb6a28c51f280ba1da2a44a0f1f60bdd93df5679c8cdedf062a3ae46c0c2862c95b3bafff0c33dcf93cf43c975d9909da6f66103f64cec1f4502ee4d93315d15420e9ffdc84ef56a32b9166c6d59e4fb0a44b71280e3e22a76be583ccf6aae90846a2b1f0ac8a5532680b6883be721fb8e8e1a05db75c83f0b8a5e0db2977966293693d47c8368ec7fc0fb9ea86adcebc1cae9c842cf857fd7eeb5ba0fd0cafad71d6bc4e75a8b5d21490bcb25409d6378efca6026279b820e69f2c1f94c929c5c4de3db4ee177cf5bd4622a046f1dbe272dae2f0fb20d087ab10c960edf2de702d3dab78b1149630fa676c00ecadc398898c4960f53cfcd9e93bde1bcc84027b10ed498725e7b88bba0b29aaf309d65f187e67aa19b9b44e871974fdef46651314314d263aa0dc14fd1c6835d0306c7b2e69fd7690c776152f59721a582e3ef8355a1cd075c6a4b3740d4c9438e336915426b71388f289c034b62acccddf6da08c6e7c8ad4053723ae19b22f5694f0ba2487cd6246f40432cbb424b0cc62c7c611044d82a9ab6d1e2539cd1cc98465079fdea2e5a932a0c91def0c199b0eaefa9478833d64a55f7b8a7e3ea2e5d17d738647dc797f2246f408335dcb70c158f3a7b49fda0e24b61b07e2148946f86c14b8b0523a6e416f179804075cca331abeb48aefac46c37aecabf2ac91f915a6de9fde77367bc985ff7422bc2bee8eda5f14e222d61550ed52428bcb90395576b2ae0e4851b1e7fbe681c6ca327bdf4d2e7c9aaee6da0f5955f4e9f4bb8ff884cf02d61da9468177fb6284d8892e7aed2b30bd1347e98aa890f7aecf22196179ed1c024a2ae8f9f90c03319c8ded568f61815f0b4629137e8caee0bbd142b45617afd5e9bbb3623f2f2a9213feccd192854bfbea278b2e9e3d751c91ffa43a0664c39254a2cf346b9eb851c2c8da696a199564f35255a58dc4513ec67e535cef564e6e6984335a8c225116de6a6f8017a38a807b5a26fef470881cb5e33edb1c2535ab8ae7d1831c93742bfe1581422f4ad06c03b3de22ada6936fe2cfe84b9e9149e578a0dc7477b081266fb911aeb94613b282d5513380f8cc27e345c7e6d960e65bef45046f0a2513091bf1844de50d997044489e757972917181f2b3178235521a2d7837bb6384346806225e0ac5c53b9e783361409953be07c11204592166a2e3fed501d2f8f12508767c657342c7c81183f4ecba65ffcd36893d97e0549549ce7a152b15e178f79332b99fff51c252617edfe76b15c6ce8cd03a6491198a0701e971d8fcbb611e111918bdf4c4b1285fcec254479d437009281d06ffda3aadffed16c81464d294b51ea7f74bf5ba6b51f0105ca7cb1b1991b8719733427a5112dc45d7fc38ca7a2b47bda29cfe456b2a688467cecb394d5d27d09b41b9726def014709f60d23e3b5ea5cefc7e2d4493d9667be87732edbeb6c30c0a2b6881ec34591f29fc0908c24ab4eb97610a1337e26ee6b81de22a1e314e669b99b6dfaf7a41907d5d589786994036cb1cfd0d76d9bed84d5a0410c4d35497b946b6377e65042738c9ad89a286c5e03b0c29d73d4b6d71da5948b19691b07fa3c80379c8a0d35f8d0ddcaf2215bf3517961bb02205f7d7684dff0693bb811e4ac72b142643d50c559cfa0066291dbbda2b57088b213e9f3790be7bf0cfd898e39ec69ac21c0e0303a633a9b6c9063acf77bb150c790a8288c7bfdb10c0741600f87bd3a3a85f264ba7fe773079d8a48eb3316f9803cb2aff632487bd7aa5c5c69ca67212168c7b151e5fb724d249446753e0f0aaf472e39ea660e338a598d649d4e81dbb205cd4138ef3259371fd18c6a67866b40ab2bc422e4ad58ed1000ef6bc146cbbba20749923a1c79c1910cbcc0138480c8e4b5edbcface1cde44f4f6caf5d8df1eb146eb87c737ab940a471e8db54688540ae783817bcb48b53115394b025d0e7ee828275cd80dcd5099fd1dc5eae54f63595e23d389e3f6d758e013708c6b6f6b019ff5b45d41098742c8512b3d00e48fd01ad4f2e84ca1bde118d7449e2419a6cdbfa85988f2e314a34b8ed80616ab7445a25fd4e830ea1e014f5efc1ce89241ffba41cb286ad29cf932b836b11e185673d6886fa71e825db52920a6a773ff13bbf3dff7d0f561426d9e2998964c0cf83a4f72854043cbc7f553174878fd230435e6e8d8cff8a450e30be88b605eb7b6b2764bfb3cd11c2f74109e147520caa268cd01ed91f7fa8639897770d0fea34e058ca35a892d380bcde5161fde5d4a3690bfdd8684136d188a970057fb64abc418a675a32513965d5106fcb8d6a68811ce7595d183dee962cbff2ba1b2f67db8d6a01e05a5a9a709b7b2eb8fee968288dc11a026702cd2fd3dc7e61df3e699472bdddac9349ceeef19ca1eaa27bb9e42a7a06e7b437345b7aeada50cbbc24ee42a8972f43538a87faafb5c54aa3ac39ed66235a1116d07f79955c49e5998edbb8aa34c4ebee8ee3c85daa75a024020dc28c23133af98b3e007e0ae5b31fbf82b8eaf168c3d834c9903d0504d448ac7d51186f317dc324b2dfdc57f673d9a693e8f9885ee316a1fc3eeceff300aa7fc8bbbcfaeafc1419c06607696bdf9ea91256141a7159c16799612d53bb6feb3f5d4c3617b0fbee176fc1dbc2d5a3bb8a9158159b5e9d715b765f7dd3b5653baafc13e8820d0997905dcd764e45fd1d0ceb2f6e52ac42a93b85d107c8979e9548fa81523f2708f50b73c2ed7be2cbe23c21bb6db7d76840ca52bd0d2698d0b5f60116d653595a180d5a3fab06ab423bf981aae1e12fdd371f01e5e10ba80f8ce8905fe1939d10ecebff9733cd86e0a696d282c08af789a7eec8d715762f08935b09c2729fda5d6511b562bfa0859a35fe3db60b7bfb747df34b61d9ab432d140619142f1dbec81645ea97c6ba4ee630e256009fbbbdf2bf1c9fa6f0db4ac52aad7ecb895f2d0a3a2b0b371b454445d337a0d025aa14a7649967026f28d91175b991054fc06283d70a0549b34e2f59643fa5fc664ad458682c95ea9ad32c9c2e01d92d3fec87d82ee2267a695a7b1dfde60bc671eebf71452f728591b11a74021d456d7564c4485afb87a055bde0b9130e73c4d20cf387fa96983311d948b52fd1c6bdbef09743d634dfce1f41548b9bccb0762898e205f54d8330e760877c93e45afa7004c43d600d31f894dfc2e5a765c096bbdc441b30e7a51e31740740332c1f32ef45e64be7aad5e790d2130deee75428b1b7b760bc97c1088885a08896e01c5c8bf6bb4e613ce19e12c0dc03c27d71380dce52486cfe3e86225730bdc07af9b419bfd7dc5826b55ca40d7d6905aa22bf950ee104b3742b423a20a158e41338d411773a06f042367dcf2abff6af93798c41bbcb302a45ec61e6189e9fa0d3d92b580201df698fb55360b464b17f44a1e14fb9d30c23e81d0516f56309eca9e988b14d35ddae73bf29614e2bdb84e56c59692058e12804d0f5033d9ac6c1db749cc13163ba9b301378b0ec4d0c8e901241bd8c8e65e70edd1668598466e820308be93c9ea9078619db87763d52407a3c56b702bf75a9de9cd86c7da598d788fff6378d975ef3c3829ad49a3293550b9a64b002f0653b5f66ad7792e7dab4f75031935e90a69154862b7f870191492d148ccfa5b4b784fc559562433e58b533f000abe977bb6d5524bfb72b600c4a94a4ebabd56b7f68154c597689d25e374921ff908ff6e8753da25f37902ee7c0992a212a1392cf02d512505c1b63aaa85e68609dbd75c8234564ab6924fb8b5acb4409906adb072caf8927328a466d39426c381a3ad4e6dbddd8998a2ab4c370dd076b19b768f051e257e3e74f2c0a9c450b9a55a861d976e2e7699ee81699eff35f7c2335ebf6338d2ed2c143137e694a092b77616a430e61319ca4d987f183e3bdf3314d86d793cdf1b302037fbfd1f3d18a746d412cd8ae5fe2a642fd66d0f5b4f8d94c0f2e082374383051eadcb34c0c5ebbc8470658579a08cd7f2a505e971cb97e074dddc69874a9dd21b34513d66b0941a61d12b8d94665ea9b210607cfd218b981e4ecbf51170aec323e3bbb51b305a48b339be5b8fa18a5ed8fb6e3b25ac21c6625681079afb9f2a77bc20fc82a1b817f412fa48b4513a87e309e990ff09924d3fe00f6e315942bcaf45d78ed936ada5ae3441392bc222c495edae699fb5091213c80174d3353542c42badf24d15e9f23b158f3cc95c40c54cb7dd4fd4db229bc2e7b9d5448d3ecd2ad3e68c68b8fd3900937611f847db2ee5c7cb10ed17e53c0a8fa9791fc34c2dcae2cdabe40a275878ec59a886b18b64dbb1276a394c7cc0583f3b7d383bc66c6ab73ff7c10f1e6b8737b3652e53aa6b3451d43a0fb8ae90ab0f9d5a0675b81eec773c571cb3759bfd32f24d09995fc0dd5dead070a7225b34d54aca7c034b1ae5e23e1e7768c428a809b7fe0d7470a404828124cf264631c3b5704cb75f762f570318c0bacc63b4398eb8c92ab669ecdcb8aa6ea102f1b22486e9d704c17de57e443268d3e88bd0b1d0e5be681fd98003c5489215306a0a34639d1f47b6eb35462a4296b693b05003f1632fc3973047a91837748fd984e1854e71536d19925f85b3e0315ec9e396fad92d0e9a6d81fd105d2867e85f02c242be7008031e359ef4dfe2f3d2c18295c9e4ebdbdd6545043aa8964e09b39638d5f4c1c04d239b92e46c39dc1734834fd86d19a8b57523f9e6bc2b4b522270abc3c442f3d9321094628fb0d67c4691dbd187cd28412301ee7e4f99e6a91c87034a5460a04117df67e75b99f26f0f2b83e6d258c646bef852848f60066aa9ab06c47cf6d5fc09635460cce65192d8aa195cbefcd5f048420b42750343150e746e5c209e65758005e0d6f12921c45c3406dd931647b4da7568383af3ec23682c8c3891ed4018e749eb65f45339f23921d2273ab468f031ed68028cc04d6c323f92fdb70cabddaa02d80d310eb64d689027fc30d8b299b00dadc505b8b97c6a5a65e63c8a6881a1df96e619c2739f7d7485a717a1c060d2dfeaa52de189c1a3cad2b6f0aed42d505f97571ee81d2bfb41d461f42de53d32ff7fc400ba16f81eb8b5add5bc2c4a450d853ff50870a245fb2f2967dd8ba1e8939464f52cfea20e0938ba0d72f3b4ba9db86c4fbd7b938d6323d3da8945043ecad3a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4caaf8fe0252f527d51b0ce35345cf6534452fa5cf5a2c5de419babc8241d69648817f575171540d6416c26cc2de4f192ccf89a45db653cca4fe6c051b76813ac1adffbed77b9f6796cb743cf4c818f86359d2db3890974cb6b855778b169419e136e2e6652780af51532b5c2caec34f0c3cf0aab6fcf22b6553ce24289cad4cae54fca1f0278ef8da594ac8c182948dc39e7871b227431baeb41f0bbce2690b0e7fb9ecf9ad5ca2a44b245fb71fc513f33263dc2ddfa11d3236cf830aa0102d7c745954c82cbaa99e30321b1c421dd1c87d7337b4042890d3b2a86e50224618cd15b9fc1bcfb66fff040fd42e483a2a48af0a8eee09853923862d05aa4cf06d1d1ebdf185525cb329896935ec1b1a05605b63b31cca9ec191c7fbf50b9fc84477c56c63687660abb337b8da16810ec8b5e602ae1cc8c7b5722d95b22f650614203ac0198c497db9454dae3ff51a61c3d0f8732f39602ca134500a398bcaaeccc30a2ab1a7f0e710f89047792aca509d116f59d7310067e0f77a60bdaa7ce7041dddbdd71046a0c6b4f119121721e58d896e00431074c2442059dc7e8e414f462c5801b1e6be7f059938bb22eea50a54c23d2ec8134ce212c672121d89e32295dd83251558e34461b8264beda57733a92b1981941c2028fe6cb65c6d1b132043d406f605425bf2a2da1d790d02b4f85a5338f253ba42a0d148ce7870346740867f4291d80d8caed62aa3117f1796cefa78d354616390a056cdf0c8aef777f92e8c430dfe1be1bbb1f4dc4b8cfff468443644f86952f1a6c4252681da89393c1ecdd98a7e9112f28d6dd80b92ed539c2caa1aa2f0cdb07304469b807deabe4b0b0689c713acb0a040cefc5e3ca697b41c8b58b6cdeb68b612b23ca0690e9e47202a0cb23bcb5073f6bfe1746a4a3cdcdbff55d3c554b3c5ef040582a18a8c793f36a8f764960060e14d715fc4da4da30fb9ab37f6c30efb37e21b7c45f081bd8c8eae06e31eac93b0553753d7a8f93bdc5e11696be005afa114df54caf0ccbbd7c56f16c008a4e170d44aca21743236de7615a898a04f3c1e9d6c6d2d2c3eb7c7141c3fb1a758acd9a6c957a6e3ea4889eae3449680dde8c98fdc06c4ae733945268c92b83dbfe8bef086a7747da82312dd1122421d4c15ec887452084cae0aff5453fac624b134e2b89b2e7a26c671ca8754700e286735fab795996ff7dcd2385b10e85654ced955e907dfcd19c9db598643b2c221b23e14fdbc0199bf9aa28e0052cb5a9bafa5a40880b74f18255b6616594cbfa8553bb088ad200e66152831f8aa0c9a7d2beaa3136b2b60ede1fd82f0618cb373f0c3e2c01cd3e62878610107dd727dde8140e241de7161c593460e717de166314632205be2efcc27c3411e7582089b28baf115a39d1786397d14418d94fc38962954fcbf502679eaddf118e73fcf366d55dfd0dcf39f2268a722ba70333f8706e0ea875fe6b64c93810c577f530aab80bab662d079328444e8dda7a3beba19e6fb40dcfb64d1d52622573d1f9092a81f785b34f1e7eaea90987a5411bb966bb31d463ecfdcec1d676444e0528f312c1e217cd9e5a04abc10a18da4d1636fd68db4a367b8562a80b26f0f557a1bbd4412c4170c260b751da0c03736801d0da452430386334a3b9ac51556a22cc88da52fa897e41584bc3b365ee4bc07f07f000427ea6a009405b8f1b79dc23b977177be63e182d17bdfabaee932187530683f316726240d2072f80c2a1efedcdd08490548fd7c93079ca62c1ec0e7825e92517b1174a25020c9c16338b854e1dd8a8d5ec990bb920d1b6810ff1d905bf033640d08a79996143b23cdf5c2721c13f1865f3b9fadbbd3baa7022207efe1e1fc0f5307fef11174da787736fe1baca13e67d6993113a7a14b71b5596feb50b6d39cff34ddcc25239d26225884e7004cc957376df3a968a576ce373daedc00eed9023e4186ce4a09a16cfdc9e5af122e5cd6003940030ea95acad931d4c74ec67a6db4a2c36eb1ac35a59d4007de594e44f16a78a85e159c80732ae8b68bd178c2b5b53dfefece469bcb1ffe031826efae0bb5bd61dad0addd6ef18f06a356ec994b5fb2535d222b1318c399c5039be371d51256c0681982dc91375fdef614faa8e220008874d4d423c20d7afd3f9d07a564ffa3ee83a934319da4646beecb382a0d0b8c1de460316f24b6cabf73a75be219052f6ae01dfd358389911aa833bc7893f34c6c4f0e2506d71ce91463bbf82c888f3f8b98b3c5b5977780d65ba453daa6ef3b4933406ab9789eb4eb8cea4893cd313ea315a6fc889311268914c982fff40b6a82499538936f3ce7bddb19cba620c27d654d44140c436b81d376a62f2f513c36519c842038dda6a28b908f7637ff3208d52d5519dfda9f114dc03739773f8ddafc568f7bd6382e33be3238c737fa078bad867417e1e3f6496e960e2110e848ddac3dc4807fd88d7bfaacc125a29009a79bbbda0ba25fcd8a2df99a57fda2a1ad1e48b20f53411453fbb2560f2ac868a40ad652de3a9c6449a6d1560f7077868189046f4bb395f1c92fdceff20348105c73cf68c2d100ddd9b85ab3c5a45fc0e8e4b1c9474f6363a75a6e0b3d5de38499ce559b3e7bd84409e54ee33d92e4fb97c0b0b0cc5ba1c4a55f78df476f2154610c7327a9cf80cc9392d89878e8996b22c8b0d1ff79d74ef85bcb2fee6bbed69b1bb076fa3f1814a18e5255daab948775ed4a49a1baef80cfc6991b984c60cce07777d6edbe38dd9343818b10e493873ea0cf6c9a25d0f8af242948662d32e92088a687ac0812035fc5e65b707164c64b460d6db3ffff8550df62f8869c357f025bf88660b8f4d7fcbb15e73301072a1a804389188990028ad4be28694ffb3d87bc12d9d95db26b8823272ae782d0aaf5d1d89c907dc604aae7239fd65f7d7d5f9f445ab39683053ef58d4fe06ffc98e11a6d5589ccce274523fe0d2c1805416a76ff71fa7e7a3d7b37435c7c80aa16a635fdb9c12826fb599ae61f1cc7d6d8f9bfc5844fe1782238fa0bb7b9a4b9d43760a3209b2cfe41cef7889eb6bf7ff1d7e9705360469afd3bb3cc351433321cdaf261446845915057aa7bbf6ffa1a3b8f7cd5f4bf2f23a8125abde257c43af9c19634c91d97695ebebeaaafef44670be6d767f5b2ce101c4b711fa2544f9dffdfa93f90ad4a0af092bb3897aa705a90a957f3e8008bd64d912f8edd9e698c82ddb21f503108ac1a1520892a9de173080202eab51d27a9d20b2dea1ab3259d376a685797eae0941a63b0109cd5de6d96fdec5a34ea827c13a1103cd3b080194e72bb2042c70393054745c3c3d1dab153115cca501da94fbc0d8b9c65908ad473fe8b8b418ff4727951f41ab6e4e057a532cea35ce0f31e5e90e1e342e24242a0882e786d4522b368cf3fec25614aa12e2fa81a36b6c5b145961a9853fe6361b688c1317ea23f11c2873e9d5192b297cd5ef31ee67232b2d001eecf72165ae2bd8930fe6092995015123021fe3ddc3ad8bc662f2311aae63617489600bd824a49922dc256491eeacc6d6d011b0f1db6c0bda853584fe50c4a434980cc8b956741256faa3f02d0b099c36c0e98ff6aadef57fcb98b4f61aea2f74e7b95e32fdffdf0b92ad67c7c771117b4aed3ac829d29598fb98b868be159fc6c6bc63a8a54ae6b1e6303ad8c93abf6b521bf801486ca109ed43a773fbf4f9e72a58804be5a3b23a11c7aeab6e84144178dce6e0b77542d35c7f9498af1a20769d85ce84bf70289df6ad86ecf2402f1e85823ac1ea5406084c46a1058c1a951e065ed6861e7b326d37c0b6481d07da8a800342bc92e9468bdb67223bc40083e9fd97efcdccc92cbf292f72b9008bf7eb7ac97dec5fead30024fee78dc897b2d07dd5eb72af79ad02ba00d2dfeaa964c4e73f0567e81581498ed8d092c3aa5fb4d8e95eca942d5fd7babf0a2abcaac37b9e63f9e80d63066d4a91e678f612d64df12f9ec0675978350e6cec5e19163bba849f836ec597fcc82851e3489d3f66eb6a4b9a5c6dde78e84a569c38e90fbebf365f004960d60634873128d9ae459b523432630333a010e33d475228ed0b81796172194374d83f1f5573adb09067df3f55ea35226dba0f25654fe43e8ea210f02414f54b397a6a147e3e1b3bfd9f0f3f269774801a58b3201bb47db8625042331b47c618390a41a173c70e6130b608620a14c26c422318012fc404642efe0f781a9e44d58c12de7f15bfc52a8a5ef3fd66aff9dfb46ea02ba256d54fb9b5f3e0a625b9740b20bb9427b7624e2dd807c3a32b4d3ad3681618a14cf7a2f6636b1c23c7570102eb41054aecbdba122cf57b8e07d32f0c69fdcafbba4c9ae981df8bc5eb057b266d60f9dec40894c3f898def0565566d0eaaa6983210250ab4698846ef3c40ddd2ede9c0c247271bb0288aa680d1cc0a6b45fb4a68a975fb8ef621bb8c37639570c5d96a6d5374944ae4f30ea518187490906d6d33d531adcb71bbb2095206f2d303be8b218ca0b1ba5735bad084c744dc7575c39266ffff3c46e186b5a0435f18e0d304677f3434b99ed930da0644d1bd49668d11b96be7c760acbdf98dc8164a380e4e88a801385f2ec5a19d4a5f73ae0b2600e22a557b9e85d558ca8dfe5aad942c5c6021f901c306ce9b51ccd176cf4c2b5ae8d3f2af0ab3b4e4521a0af15ff9bb1043f1dd31e357c3ac237f181ca1d24c36a2419cf4c247c958614e118f35827ccf5359213a1b620433e82fb8aa886c3fad8fb5dccb63db29b542301c9962a8d85aa058b5d47df0a28aa76e19bbb728edfbd2648f6c2bb79fcedf669d433ada0012f193219bd93956a11e7f2e4ebc63ebf0cdd8a452394a18bc1929563a152ab294392f159126d10a19005751bac5d7a92ed5ce66cd0320d5e33b3b0bbe28502034a800521df9303669cf0d0c92a4713c6839715424547e7d848a29ec1db5b9b4eefed4aa661187ca69a3b0ea355b63c04a17060e1479a6591330ecca000440858594ab1b2510fbd4bc8f32452a10d58e6c26fdd3fa7e4ea529c117c5424669755045cf5044846dd7130012abfc7038488824ae2a11b24747a61b396a13efc32230789b1c3873ebd5b7504dc69035f332d21354628f8d5d02c3dc8d57c4fdfc50a9f398132e5ee361058c7bb738c2e8c18f07d175334c274c3cf8c1fffa6b5411941a731c7ec9ff1ba6f2ebeb73212777943f2ef2c4f98202a49efce0a766362b9b495aa3bad244517013598baa3b7daa476e88b6e1005d41f7a61c4a1461807ed19e9823c0f9571f65ae9e3f72662815b00f3a2a50a80bf4068c47227aa6d6547b7f02cdd9e8e5fa9f81d857adb3b45264b5939002f18a2ef66f0e47419b51c2ff5ed334dacdd4889dc6bb898dba3afa22497af1f6fbe841dd87e4c1a459ccae699aa180e95846d4b96eefd965156044876c2356501aef361982d4fc0e1e29fc5e7377ff5118e043777ace711f1a35276b414c2b006c6d3d4bb73fcf9298e66e294114122b4f90b8a914ecb40f90967d2e48157d92cf3988f00f1154b93f5db4e43d385ea0a3f793a097b55fcdac9d78d46403795880745ab0c953cf2bf9b3f5020df485d183191071b91b23cf76d9cb3788acc72825289922f276ffb2304738e00a1bc790f6321efc92015f8ecc4d811bac03c7f699fc2ff4bbdf1f0bac4a8f3f2510a28ab48d5316384c5d907e8f9ccfb7b41816cbf4b41f2da3edd870e23b615d0d6bc82aa9675278e9e896ba3ddf9c59aca8d14ed61a5a4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hecc7bc994f60a1bbfa91eaaa36a559e36b281dc1e31edfe285f1bb2ae4e5dca763ede08108cd41a78e5df24bda953a12a54c64e3049e01bc64d1db336ca73daa5584e9da7c873635f4f69b3863a533219b16b04180415095d6af08f01a8bf8b2456356ecf592865e62ad2718da8caacb80de4d1aca18553391f87e814d5f2376acfbd137d1308b1f92f9c2575939c66b763dacebaeffbc68232f9ea0c583497bc910023ee3cfe7123492db7ba0f09a35b4717ecee5d851b993f9fa314da870d1ebb96c1d65c55f84fefff13ce6c224e1d5bfda9d6283cf3194413a18cfc091d5607553b8aa3f9f0c98feff656af180c0266ddec37c643aee2db538b170a441f2cfc14542613a6c66d909281caba65082a1e440533cf923b6c02c1fa5abc4408d9b2798c20a01bca13a0189bd4836794548ddc91c512ffc5218c384877966cc956d8f5c631d4b62f6713efdc880cab8b46c80c80c41cc5345d9f0c2b915171fdc6dda7ef54b8dfc9080d9301bea60ccafe6c8bb4037e6fa43b17f1ef5a1fc8ffa7699791d1962033b1fd87a413bd42bc2c6b44ee3dd2d23798f5aa3c1767529b76cfc1859d1f09a92585f3166d657f6559397a6e3c79bf5571a9333116c884fbd04ef2fd34bc102f40ffb2697cf617d371756cf8cc43abc92cc9cd5b442bd776e1efeff24e1113aaa45bbe67702b34da26cfcbb1cb4646f4ea004fba36960c7b2a814c95289a9801428934d81fbd50d9c51017c83d2dd31f8a7a7384be864ba3dd49eefa7c1e087a05f39741eab7bb7e8d9fb88cbc29a48ab3b3864abc6ea60d63337cca751aa40fe9f8cad8dc9a213963dca3ebf95449bcd4594325e80b266e537a4931de3033c080d57d6afe6e1e7eca8d7ef162b9ce03b686553da49e7f626d06907cee26ab5a768b897b4fe8fffe92e10f392dacf1eaf7c956aa07461dd4f72e1ca6245eb7188a602b0687b26d0f9f7ecd5c3ec8ad4f0c4a805e9b123f0d627fdc3e393a84ed0dbf7680eb4ac19bd808e6926ca1e610b4c15c159020ef0dc43afcb28372010ac29500246847f960c53f54b46808234e969cfbfd368774313fbbdc99ae2ec86695d3a6bd7df70a857fa1f9ffdd563d7242c98a26da8e51e1579a4db515cc63f815097d7066f9b97e3bb66b149033e6fe8fc5e56d3943b4268ae838c97ef8e92c319b7d73b7a9945449ec9dad04cf49a69039598130c33a746c5b8d39ad203000bc0d6ce85976c69caf79f203be2215d115c141e4b185ab04372be20c7fbb7426c4da0fcc40898f83f2584b72853e7c6c64706a1c9e2518c0d5e95d1789d2073b3b8a5b30ebf284f8f67878d53c84e6c78fddbd5bd97f4084af26be7ded583dcfee7769d3908eef2fab73255c5f1f09794c03d57a7645365a3f37034df106315b6edf1e7e66ec707ae8a0f59e917fefe9ce74790934caf71a2bfa317ae728c4de3716f281f792bb0aef6e89fffc69293b0a7db62a1606cc63f493443ee0cb66fe4b03c61ab95006b56fcb69d865d35a74af30462ea1cd2793d00ab58e14011a0e6bba02c0c51f4089d2c0f424f4d27332d4c199a8367382c9f76a9fde4102e38c9f70319934a109b74ae24833abf83ceeb8f1dd09006612bb8e389e9543951a8a5b631ae646d20166d17ea2319c5978034a21a73863d4b230fb93cc96ab326155b69a9770e3d8ecac8e5e69163e25bd85cb083bad226a2366118e18091e5c6204148cc42eded654bfc29a85e3d197c90d6189bbf77eba2ca9c6377168e67535f71b34925a7ef53f679917d3f8fc341d433b148e45a7b355ec5ae6807b2fee49e4bd41551b787582dd6db84926146495af77fd5a78e9846ce51a0bccbe0a49f569c4946c01a4a9f3aaeba432f3e5b2cb6a95138990e0e90f88469792e92f1c8f3d8e53fc6a6a021c1ca9d60419e833e33b8a8bd6e3a5140d3c578657641bdd5cc20d3c7f8bc75cde3eabe470e483aa58458e84462a29183b705f8f136f1f9609d1ff1a923b1ce56fa9ec6a8898c1de15606f09be87dd85d92167a6b10224ab8162100048e7d89414e74ccb08fd1a9469bc8c28a0a8918bc0becd5a17eacbc0b5689aa479f17a929df67531f395d5ec1198523bf609f19b6e90cd6c8fe872192fcc5b102fdb731e677542177617cb0433a14c47de51ff82f924d98c60f647091a0bd30628a9a354afcc5b3ead14bfe16c6659f84a0faf35aee7072e6794b4f4476e5d9ace3bf549c32a90b321db3239ece4bae1ae5a6c6b3b289a709a8667207e65bd346e3f3a50e0261ee5bd3208ae9fb65d3e6a44c29b2f1101bf25e74e2fbfb4b9d47a299b56a3d6e3a67791808e5ba1d0146005aea4fe8435c05cb332a52d570f17a73d6ece12db1705a4986ef6f899f860c0abe49fef0c5f0137ea83a3979ce26a8950856532abf69ec66b72c858bf76ee6b8c2b386d4146f04e7b0482210dce336ff495c0382c7653326ba9590dec6755e882cf785777ec5e7b4c783842ca2c87673765950ae4f6c965dbf40a39423b69f2da80bae36f67a6fa85bc0306f22388a905365cd0bcf2e8172939ae13179edfba701eb50050a4672fd2cf81d599e78ade237d438a4b4b73021e18089d97b3e43e94781fcecef6d65de0cd80e6efcec4c5fb01477178c448334d025e9d817129c4cdb86ba7062be7e5fd0c4c5071becb8b07a5ef3a7983b917a2c0cb91bb4bb05eb649a45e1e63a08b8ee708cd35c0385456bc4fe5972f447a269c349614ddc3353582c16771dda9c23857b0d707800684fd2f26d824ba594e9ee4356e10c4e30d5b4c4e91e722ce0cf8ea4a39d5e16d872f72ce2b418f98ec5e251251ee262d54557ad630227411084e7895e0e1cf51e5e6bba65d46878181b3f92f4ad94c6edf9642e975238f96269880c54446370e8d796e99b1b80b545bdee958db5bf2a215d38d3494c52050f56ee000c9d35bfda8fbe27bb76cc4473b973903b9fde935847fce540040e6f8d904e792a992a861a864a1a968c477e5dbcaeceabe73d76523525569db244f3c4f43dc17a353cc46d87f8368b364957b03da5c4057b4969c8acaa14106fff447391056c02f4a1c5c998c259951aafd00ff451737597e9f542ccdf5ea06b34d966fa2ca410238d2d8b54ce5a4a43d7d76667ccc73e0f832cbef71660b3e42271e98668905115d9763a7db0b894d8e94bdabc5e070b3329e0a034a8eea1d3a8467841af1bfe83ced9807f344afe51ec63d8b70eb77f6c9b0847cd874263e324b7cf6132b4564703469f595157d1565e71b1aa878fcd04da8a4a6092e88e3a0b5615a7b76441aa074896a468ce022f3a95c1d819251f9fb942c3be0c857951f5e22b473003eb9c2d0be005b47097876d196edbf625c2be624bf93111056629924b8643722fd254af74a0f245f52a39a7c18c9de8ab6802825b181b3e4c4b4677c3e1585b0c94899aba380356854ca5f715692d38e41ffa82b3b2286cff757ad06edf2638cc030907a0dabfbe8fbb4f06cfa09b5d73cc9519b0657d2251fdbd0e74922ff1946898f9eb96d3f36291ed80983a9dfe949cf2efa46ce16941e2f8156fd397b800f12cd3eaf58ec4a4350991d735d9f2cc487da1d7d6b1a9b5ce4f06e8f60107a8733bd5c324c809963942e8b2b73c33072c29a08ddaece3ced6af62727bccbf0b1438f7c30b1385d7e68a30d5b0f90b6d76372318138c5c3bcfadbbd8f61e9083e9b313e0601f6e8986bce14683ed48a9b61e3af7946d1a8e48b7cb22d8b822d476a1ad047898c8f55b5e72d93135d661286d9127be10d03ebf6b9a9fab628bc0078ecf8ca3da80d78da324934973feceb0beb951816a0d91fc12471f620d39174aa470027679cbf871bc6d40985ab7f5b6dd24574a79267b30fae27e999223f2208a045421df4cf588468c2af0d7f5fe1c2bffa3255d6b1a95327703a3f48d1902baae211149b1ba8905667b4f10216a3e4d92cab0471a99606812536404be43199748b8e75d84a42837ba8a153a5c467715dc10a0cbf0a1ca31bc86e08a6c544b368ecb1d96aaf7a5421d680f3f272c3b753f810115af6ddb92132a6f2adc49b3cedbb74b5f4a0608460cc0cba649acb37c741d932aa60028bd55f003228044718cbb6f7d65cc209bbbf8a78e530a22596729b34d08bee430fecad78379772fa07dd48eb6cc594c64c000bd9b246faa2380174c6eaf91f460331c731ee9282c5418c5e82628f24ecc37be51641beca468a9d072b44adc4a1f7dad29a9054873d909d29b4cb9a473bf47ead0ee50542d11eb8cdcc873036c7cb5447687c979bb23435ab80bf9381eed13579d8a09f0fe28f2d7b7d66db34b3dd8523754f54844e6a11d14d37fba3ab11b751907a7819f0712f55a8c614d2cdafa168ee7f2789537583067685d72c5e76121c479bf0c2cd3bb805ca68b938a62068cd96c5fc23a669c6da1827743f4a4d8c894ef3775fe222feac5fb7aea5bdba45e00bd95a7913cdac70e28132b89f50ed53997c39a869724168561edb22dd9f38b384ce09926252fd18d63c81e0c32fd6c819836efe3403282a464d137e759ddb9b1c9fb2adfae0615930b52739e58b553313685a8bc5a9b1f46ebdda56895215cacf8dca96f63dfe345cfca9e26c24eb10066f2aad99901f1d4428d1f851d46e050fba7d5725389ec20d02c4973343307cbd025cac098f6068a6981df9570b03deb2dc5e653d9d20d3c178bb64ed6665c547ce64a19407da8e56f529804a9bc660a2d14bab2f38158cfacb1d7d5d2277744b60d0d841ced466d270812e935d47767ddc301713f051442a0bee51a3b16a09990507ac744ece03f289fc0439c5d29a1c528cef5d5ec9a4a76ee2b5003e557f65931eaf48b694af930bc64cee9f19127fc98b11831878c28494268ede029f2ae9fbf6878a23fad8b21ae8f0512b1985435de53e2d5b0b57e7c7579f43ddcb438817cacc62e44f17f55b141a264030ea28f8c5263f6884b04864752e5755c6687dc1e095763d59214a2ade3321521e2ff944672326d8d611bc85fbd5a396ec97e4ec7f144047fa838af37297079b849134b12071523bdc56e109b804f2a602d2e3e42126c42f91e78c44b4a00f16dd0e13553a8e3727bbaf5d37739b959e68bbd69196d55d0bf25066f4a022cf2d80e0df546f2f38f49193982aacb5f80482649ee4490e16b86366050f22dcd9d80e8d9376c36a1d6568ff9ee11eb15196fce58f940e3c9a7e05e97a194e2ee74e80be26ca69ae1f09afd2d99c85d210b5fab01031ed94dc2bb8479efe346d537852e0cee366222e354505271706554c33f75efe96b9c903c425dbf7227bfa17fe88896b6466c01f75d71f99fcef812f2cf161bec7bc8c3f9a79b1e54e3df0030840b832fb2845b574ddbd7e0ce0a6b72228fccea37da952b55d146fc5e90269b8da6f706fd44cfd8c8602b92e1732185d7ed0d69a4444d20d292b5057142217fb65a9d25f48105a99278a84da01eac6e0d4398d19ad5023327d5150cc2f799d2533be81ddacd2dfa889a6b50e4d1c5634b449322c9c209dc846e1a3d0985d237711b48d10379b693fd325d490ae397228c777cfa436b434cc638afc1567cb66104804cfd7973f2adca1134b762284791a9d4f86f40c5ec30fe5adcc75cbb837a04fc73728488817bf881c3bfefd7e80c028b52e2ca770f1885b86ac6e09ebdb1050f50dc25534cdb792b56476cbf42f4bad6c1ee30b6162767b10c0aa3dff84355b68bfadb6ec39ab29afa46e27a89b5447178466cf0e7569d53980f22f7f3545554;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h840fd3f7e4cd4e45462a9f6e7e85e934102f940a4b13189f89d2b742fd1afe06d88989740951eb848c0b1c7bbcb4e1e3705bc2c216d69f7e1d8ce40ddf60b66026e7499a3783e5569ccd3389cd1e5cc578ebcc3d2d4968b914057cd24461d7d1407ecdfd6ecb7f314366e68b8b6ba7c4cd78ca26ea50d321e11c3750f99109043ebd528228947e97564d7c66f39bec1cb9da02b3a76e847c2ab3ff733cee14598e764f067c152c71ee6c7be3da7622dcca38b3514bc2d9fbd59b0fb78af46e00a4539ac3d740af30aeafc6a51478008393ef34df0d98741f91442f5b7eb7f0e07d66aa49bcd90d95914615c9766e18bd0738cf0ac139d04f0dd184aebd2665566d929f24b15242502f6113d325fb8aa91a523d9c400da247d6dd4f0f47ec3357139226b9fa371f2750abbfbdd5cbe8defef79ae5fa67cc46a9c1dafcaea4c07d81219514318112d0e1d4fe1425e8e8155b3b335eea767b2f702e64ec6a5dd85f72089d32305a804e43027c04b68ccbbf86d18aae66bb76909ec5108ed8dd592ad415f79d2c2b36cc7fa8f097880e52538aa2509b6574eb7867cc9236f9aa5c4f8bf2dd0954050c47768f3292152b59f704dc0a0cbb3798a76c44e11cb9f921a794a4c3aad0de6ad53954de5adeb3e4230ef26de9a1e07568af374835cc94afdbb18734fc1d0f767bd9263b0138d4f0e2a6c55e8ce53f89a4782c6b8f1aa1fc172844d9a21e24cffee0ca86205dc0a96f79ae2822ab1a31340531010c77dd85daf8de2631bc3cf8ad073461034f4a4b494f532039967ba839430317949a5f1804af848682b41cebe83adb3f72be2b870a1ae67fbedfe302e768e8ff5c6a11fe340ae1166f8e371973764ed57d3e568e4f2ccbeb59ccfa5ebbeeca1c6f898d82f56b19a45d04d403f6181c1827ea917963914f50f475bb3775770c0e0af55ced17d800518920950239e5dc3c3646e788df8c9862c0ef71a6f8a1129fff4763b387c94107689179d1a4233078beec1cc21db555ca021467d025d3ba3f554abf9cb84c2778a41905c7d4e91b65ef3d264cabe00f5ea56e5c3a59b8da6333dc08334c2d818b8381595e4c324bcf37533c0fe8ef12b1c66f71aaa081bfb9ad1ceca4cc6ed5db41d544fd9cae9dd82859768fdff071b390cdba9ad984466808848ae9c90b009648277276cbbf21557dad39c06721c7bcdcea6366ce4f72509048e3baac0eff1318a94190319e366dfb5aaa353fbf7666bb9e90bd80db414f522a1550fe16107512423b17a529f36c20e7e8b781721191e2287f8176fac3b66fddf05267918044ac2455b23a776174078160a18c2c03cf665a0a1714500f3ab4c802af3836117f448e6ff9fe1619828aaef77d69beaed0790359f5d3cef01eb1d178a42aa198b5d6e3a957a1b41cdedff3d81d255cfeb790c2d8f80a4610e2d5578919ee877e6d1573330d521ec17e9999fe93434def8434caed6368e255e10847062ac2e5bcc567b506dc2d81f416ded56f0bf43233b597c938bc7cff264f5b61e216ce038392083c72ea7038940bd2c065fd48124ab415aa72bbef67f3f9830a670d3fd3e17b0cf237883f814344d108775a9fcc40d7d8b8dc912725b2a64aa4e95f304ef247a87648e1d728d7169fa6e29dafdf2e17295e748ed128c2011a2b31c5da5aee4f8c8c615d4469b89d349c1b889854cd13ff6222136bdeb3da549cea6efb8d4fb07af73f54b5cdc68949846eb0fbe2bcdcb157050099b7fe081d51f6d30fb6eaa3d6810ac6e59f770207fb97fafea9bb99f1ae205716d23f7802a6406f29d262124a6452fb282abc80eea4a3a2cce9d82fd0b24dc87014b9db2b5e181aee810b41060c74fa02d68fc24f80632331b3035b5467652e3291c086c92b8928f5da161fbd60e0b774a3b3a755094991c67a01aa2698d567d2f35e90d716222c70d429980e5a13ed91b8d7a086134a3b2ff12231fdd7a884da347766aeae96b47923a076b5ef90ff179520ce610571fe45dc096e73e5ec9567b5814c694ad1c8fe5c7b18cf717c7f742e610c52953a282b333e9637f9a6ee49a6e2d70933c09d7afcfdca18c76bb08968bc9aac65e744229eb9e7c036794ef5fef23ea45c43a62f78dd9e7829e913fdaa6cbf544367e2cbc8f55a7a19911f2202e0d40a1c7754836b2ec1dc6d37d183a34008c2788256aedf49f03423e78be8d29c867d0a9c8680080923fd6da871d78671debbea3ec39a7e3755be880177649ca2916258deb7ecfb4ec9f8026eec9fc2f23dc86789322d636a6fcbc07f00c59ea3877a829db5dd0831b5fe6746d50969e803506e0201b0142aa5980c1b700f2c6f0fe7d8e9bc28814af464e845ed35a2bc5958b31dd3a7d0946c16e3db7d4a707c57db06d24ae02cb918397d2ce3e7c59acb2fc27fc24ad68072d2dd5f6942bd51f70667c0f536788aa00249552a5bf5136c3cbfc17d89e7d19360ff16b792dfcc6054e7848b36b88dffcc74f836a7a970cb88c44c3da5e2ceaf0a2a19a79e781ec294cf015c31195626e5a0414e04c83742c40ce5b753ebe894de3181c417bb8b53191e5cfc1fc5a745713105ee2a6fc51b5d5a1e737e2c74e38df0f993cce5d3f18df6c8ac2942cddb28be71c68ca01735865225fc622d7e7fadf48b141b3dd30309ce0160a45e41ca67d9872f328e8e1d8a181dd99ccd1cb92915f489dfcf5b1f2a7f232c0c67da27e07c5102ce3dfdf36cf7773aaa66e2886c74aafa3d04c438007d0481a3830c05fd29b34e639fc4ca2dd6f40fefd65d7eb89383427aa24bbbc59f03dea58e36d47c36070d88d626b4a0f9b2260ef07f0daf6195681b7a0c4ed8519e0d642c217709494f5a383834e8f5805e987ab2c7ba67a4d34fce50927c6440610a1e20dc79768f259ffc8b68632ef87c8fcef06c9bbd50c6398fb358cb1014360f189845e1db41a0bf3626dd83c7f866e20ad9fe8fae33ab7d3a505c42dafbaa862da923c64502962b4d35d4f10065a9ea085e5157525a1b545455d98c510fabf54b8161b20f3c17814d2b2dab17330f4f0f547bbe5d949caa3e87275e1fbfae9a8ec677f60dc0ddcd7b38dc6e402c5cabf9438b159614eb217e4f87e7cc38f900fa63c0a68f5181bb7344274946e035dea9281382c1c6b0e04d195f64f6db260d1c8cdfb616796a2e7da3ce25e251a157b07690f9c2796dc5a07265d202e35adf8093a5c5839885acd4f94a6d40379874c88b2a3b429503f546f9126f89e1a940936de73f102b6bad1bb2fea177188d1e1f84e3683a6508b24f30a8b0a83fb906dccbdea7b16f9ff3a26f9a855e459c41eea738d541594e2fda138a115f821c9bf74b0b1b2c71c75ea06320eb26865d964b37af44ff434e58bb7f54525d94722c59d7229db8271a73b7a8d516946bfbd7c9c784f208e50815943f4895056ecdb6fc9cdfc1683366a70a9468ad30ad8430b9b56b5ac1a4ef1c684ac4734faa02c7a7b7dd82221afb42a19daf706793683a283e89f8ca2cd16638136f08637734efd3b589c9c35b2214d23951db528585d1d43b23ab749201822090496e2ccd53afc28575ab2232f81a60302c56ea93ae4bb22b71514bd968cfcddb41e82a2901373c0fa92e31327097f10a428c0f33431825c7fe755ab9b7f84e1d4efcf0375e27a66333b894d0f1c0f3625c3f88a430d0761540d7bd17863172a8cf1cb22127496b41accd03ae227945e8f9a862a809a49db46aa544915b7d2376276499052295a1ff34a381c7f3e7e961a1e1dd997dd10c8ef790e9cebcd6c64b39a9c89bfd3ae06551cd085a42176a2f9641b3ccf1ed2ba9e93173b19feb179da5f8700645483401e967acb79adb648f8977e2398db5ff4cd4890ce9ccd64db2c1d348cff5e3409fae5827264eab8f17080e2b5abde493d1c27204d99bbc3c3928d4b5b122175cf49211e866732974a4d0191d4724b2698d7212314cefd2d7142f2dc0cfb6c2147ee223f736c871528a12c10cd1e913be5a63532478aa01b94173ccf935a4adbe8f837c7dc3bd2948442036b847728a890c091b48294e40c7e55cc8fc4120fa312cd63b745b73f8727a3cf0b75c79513ab76fea19a61e1633cbd350e742ec5210852a2e6f549afe13be44b00bff712616d4a23a9f4d9c78e5146206cbed7c4271f678ca8498b88eede130cc521338a215fa14ad3f72322745310ae1d842095dd0e905a9480dc2609382b409763757bd9647ce5d0d727cee62ed008aed3a10fdd0b8be6db13f5221c86ed5b79926fe31aa34f3e5e82c24265ea218175baca9817e93e987dc86bcc960d89c33e119d5a13a259b1b75c1e0dce4f2e35098255cb2b5f0ce3031225da55b4668b9b98ee0e85af2ae65183fb7972f7cb365c1bfb9a364bf58b3a48a544a57c5d390b7d7c9239918689a2dc5ea1b4fb29bad2f54740ba578ff35f42ad4e2458fe75842c49750259f74d0152dcfea88acbc9660b692eb8f5cda3c68868d43fa17b273b4c6d62b5d68d0452add76bba2c789c435e0b11550c6b95ff909d22ba5b62256189fdb093ef73551c3a43f44c93190f88c73e6e642debc76200664f8d90088949f31e9651202e2705bd808c0d24990c016a4ded53164859fe1490ee4e3ddf596295274a7a3662fb65d514cb40e4be21b84a9138c150eb444c020bfc99a05e93148a71ca5d2d1f6085360330a3177b13dcae2b0a75d9176efc97cfa7b681791f6f82ecc7d478da262885143f7684c76c11cc045faa176c1fd9266d2de7b765fe11aec48653c5d0a91f883e1eec721818c17faf34fc59dfe9d72571fe29169101ed68c5747da85b24d1c7d1b193dc87ba9e273f8a794886bddf645b93434264d51daac5ef96cf043218bd17b989156424c741350f8106a62372481c1cd1abc73d0dca39ee099d5e5f50f9ac4148c7745986bb7d4022292cf4ff95c5df0f0972bf7061192aaa1392f491f7029ca9d89f03a514d69de338bad68fe608d1edef6adacb146ed48f202cde37ace7cf929285ffc28e7cbefc73855b9125b620faaacc6ebd2fb89a78cb5fe9d78204b91b664031d3eb2cad0346df409d6abaac879c08900b74d99c0efa036e3fa5dae34d1423efb201097f217abc00eb90aaefd5d675fd9406e792c835c855a02a3ac9d4c25689c274b1efb5e35dad9b0c30242e81343916111d2229afa740191f81665fe3c8ee76ecf55191c8c10c68c4caa172dc8ca70872e929fa156de53783ff8f04c2649d27b3622061e32f0e745fd32470aa95b1b4ac6e02f4769a4fc64fbfdc32a158c623fe06860496db660a5b1753a5a478d2f796070ef6960d164a915d24464d8f5d233d02500f06c7cfe1d3d4bd258cc47e690364059d5f2f172163102fc6cc25f5acaae9ea7f5b6b014184596d47ff654768593291e5b9c0ba817084bbdaf3a5f31097ee949e82349d714aabac02a058230ffcb5106279c5d6f0dd4b56a5521097485558ef4240368bf726bdbf58f50d4f85512c9c5b8a9e0ba58bd98a6918a90160d99196897d3843d106a10bacc41dbef539ee244bfe1bd73c89e861eabaa3732fb08d6e485d47ac94534b8b229f39bb6c40adfaa3535a217e79d885cb1abe08e30d629a8ee8a5b7118782be45d27e47bdedb590f012efe251bc59b4da78280c20e8c54c1e5ee95e5f8ecc2b390fb59cd4f468ef0a0f0255b3b330f7093cb98569d2e3ca2834a0db929f23db49f644b58e165660ddb6eb7e1b70f8cccfbde4e59d6c39da4eeb32025710cdf8ce0e91bf89dcffbeaa469e138f29f251fe8f6f68d86959cb0da;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h411613dbb71e34e5d49b5e443e2e0015bb3460153018176109531c3917bbefc1138dc7bae037d4413406c2e69a2bf139a7c3dc3f0d78c543f2f292c6992793a87a097fc87beff8488d193856426f7c23976ff4429a1b7d5f4aefaa948d5d3156c3d680afe417f8f43fe7a37e053aa56d84fb035b35fcd540e8e18488d03d7ded94a5c8e2dffce7f3cae93eaf37ed2acd0f676a8c8ea37afb6f46b1710a92116e7061e20acf98ed198d6e304df2e84cda36b0fc3571b859d28c3e371a5cf875f1afdeabb38ab11715688882c31e275de88ebfc35a665b159f7ce964c825897afbe1c8fc76c10e73dd51a087b056c80a96da04b1da6a505b95a383cae385638ea1d28979497b8cf6ce9cf5f2fc5f75465e28194b5ab69fe4429c59ec9e271aba1772a4a4e370f87c0c38d2342c49e0a89815d8068b79d59e980e8fd68d5e5ea07f3358be5f28dc5b466786b26de1ed0a3f4d48bb93b5381448785688e82a539ce5c1468b9bb93fa08339ea9b3fe48b299e38ce5c250d0426d37e7d51aeb09b972e3110b2e7eb4a203947f1a4b6b16f26dddd77651b86714dd634d1d6338fbd86c8e0933edd8357261b3f5778c1f2278c3dd7069f75f912b688a365416b67c129c07ccf814337de42ea88e0b6c5afc8ec6dbebb46664965a7da772a4c59e026e05b723d1a6c27a0a1b6c034e8daea710f404123ffa5ab120b687105cf1c50d7f2f3bf999344829c7dc7cbab0a0bf5fed2585f479a46d54b96fac667255cf4b4628eb64a2291669dbbd1eaa8764dae929bc712ec7dd9152910212a2fe7d41d94fbdcc1290ac2007a2ac20ff3a190bcbb4c708cb839f77f21ee6b0317e0ee43285f13832b4b0ee2a58d0dc55ae77389397dd7443089267b31f0f5327af39fa26dc631cf9efa8ac04665b50c524b59fb6c1939c771cb1939d1ca4e4a680e4e1d4e573258a91d2836ff7eb5e023683ddaef972594a7191dae50055a1737c2c621580c85f7a0a1cbcb8dc5d74e98c71bb8fcc7889de5bc4ddca90aa6ece46a5dce3f3db066c9bb854c79b49ad10e4d39d085f6651865eb054d72eb8b0662fb4d615e9b170cf4de6c2e39fc991e97bc0c85a56d2b774e21b5259ce0e03d1655e8db9f4b88d69e573e0c9e26fbf5a17ffd36c4db0eb3e6778da70593a3b508820bf6bd9cb782128f776f96f20ab5eda1a96b9447fecbeefb39f7594d601860455e8cbb099ac90cc6d77191b6c2f1e0ccc44d182c025a1b4cb7776d4a0be481bd2d96cac7c2901935e5eef0e9ba1d64e97eaf1b7dd614681d17b2e2b652a433440adb37c3b95be455a7ca3530a96ffcb21afb8560ecca5fb687dba2a765cb3ddda6e8d01a3b54f4815fda9883daaffe924237f331129b96c02584709b9260b635d8a36a0f792e7e13a51f91989b2f356eaf82406777d18780b26e56d6902810f60ae1f4f91afe2c07283e72e9e270820b21d1ec5a88253466896f90a9ea40be85968ff4332340ec2e920151cea8fbe11695d2874a3f52a2144c9ab7ab64ab16e201e40735c0d6ac3d3740bbf1071c09ab694445de9b43cab3016cb8a57aaccfa319f545189f0d7f1ab5aa62ec25055e615d312a59978ceaf22ea47fbe7f3b6508dbeeae7374ecc87d3e257f5a2bc52c92c0c6dd326e20319086c45440267d059d0369f7533fae9b8565e8b49d77f1c0d8ef544f99ad5a52bd1943c1af315a4182bd8b692e6712e661687e0411c2340fc4a43be4356d6654b332b3d16579531ee3dd1c0918f76cf9803a168a1c2534880d811ec6e0d02e18100b2dc3d8146c15832118c61418ff9c9da6c037fd572f6a37247700350232c43664e1060c1b126bd7cf6afd2551ccf30c65b6f3f8d707a2ae2ce8f5d44a2f445b2769f675cb6521764217df12b6d115567973c310f8d363aa00569b3c6d984299ba8f73754c43211fe5ad1e8a3f2b0e932897d8a2d2cbc3068bc96b470aaa505aaba562857a02344f2d106129f7cd644834a5a9fbdb3cb2491754adb8e0d9a9c9bff01d2bb490d79898ffd1123f100916ae187c46ce80e0d6548404c2f84cbf0a3b65217ad6ed7f1215e834454eb877efa6225a6f6a202f11b4ccbc6fea0c3d04f34bc4464fad1c51aafa07618eb2e7938834170e85468413000b642fce9abfc0594c74ca0efb855987cd46d09794092884bb3fb962d3b0bc0374405f38a5fd0a8efb51ad6ce6311dfc6b21e758055611a4ffe575000679c6ec3a09dfc3684a0924b24318f3a0d99c54acf38c887c3e319a31aedd3c91c5bf3329f31b01ef69db3f786769afac7a77403868e8c6c37f2dd8f73afd193c796474eca9e6b38fc032382ea2e71b26c78695dc5df37d11740dc6090ae56f9e4b2631562bee1bde005177413b9b250442b5557e1d028c70bc5023a0cbff10e75ca4682b9cab995679138facffdcabb0f65753b2376742abe544499cee759e63cb9ed176c810b108574b748bc900727a4e127159ff718b47ab04c0839fc7629e668324f2c3223d962b46f020d0ef9c52395da72057bdb86bcfb3c8232f74532d4a5d3f84a639afac64ca65e6b848f6aa69111258944eb398f082c6160dcef17fd1094b6e3e5553d6f870065f257874e15077c52dfd5722fbaf50bc346952e789f913947ca300efffbc666e9b9d3a902f85bf3c792c74436a6f4edc18b7e32ca4a1afc01edf1b9bbb225b1b1bb0d6ac42abf310d829df217d49d9a42abd1445a8df1b2febe71e98c3f50fe7afc7799191fcafc5bb53329e2cef6363d26b047381e9f1370c697934e3a557735d64e6d84a8abfb64490a9a5f8176cbf5a58f3b6d14ae3f62e1517351f370b4ff10a368c2eb9fe923e060e7b4aa010c3c6103042b31e3659afa495a2ee99c480025499c08adc597b7c6874ba43b9b75dc3ef6b38891f4138a40eae5d94be41ad5f9c07fa2f2269db46ded2264618ec30c593bbf9ac5402da735f5707bc9dd9693887d3e0eb0d92323be1c06c119b728c68e6268656a2b5a3ab5275830dedafd7015d1951809ef2a5065bd56473bd2a3bc588e874e741f4b8c7338fbf80568fbf4e42b038640ebd2536e6cc6f032378019d6356f7cf8770e97e9e072919f6e6621ad8b60a55d5a3cc97fcbb0b75df0983aacc84865581cf0fed3548142d81ca9d3223eaaef8a7f76bca11642d6d4cd5d86ed8fe94f528e0e70d3e8c56d1b10f1b635ab865bdfe57869abf417a49b55f4c9b3f04cbdd505e6257b4146e01233b02766da70842c43c34e4baeb8b0ab69cc3b276c7708b51d45b0df7575b1cc242e747d5e9634176f6c8a31e18e202042cb356311648ec9fa94f5073d095d8e9d2a429b9eadde17bc971c857690ec9ba30d52ecc087b5df1a4274f9defa59521be430b111cb6a479176e2a02ec8bbf7880780efb2217bc3c59db801931f565f8f1b43cc3690fc92fc72fb19e32e22b6fc9a4b23ff0c31bab3b8092e14c9adbef4199d1874643d58143fc5f6e121a958df3e443c7adc7c4357ce7a0f9c52d6e9fccc4752762c3c6249a6580b762220b62ab0797782dddd3e10a5a156bda022dd361157ee38d399c37090be61553acd00bdf286ce5aefed9129df06f9413f74e312fe0e7216e56c2fa7006ed57430ea860d9fe724aa63cae2e6090fc31e9f9ceffb46a063f7c3c3d26028f9f85f11af0f1976b6b105b412c7f71564c3dd78af77a0774d1284f577ba8c0ad89787fbc81e9976bbe19c8b0dcfe3ab39d6fbc5edaf403497bf1edd67604494e0b76e85745af36dc916942e4413aa21534e0cc9bee7c81df0c94b2cfec40654b3b6c5b47824a259402d47cdf3c1f6091143f34f841293b9f51fda560d58b6257bb1954744ed7bc208cb692dc63af6b3587e65de26d1fffcfda4ba77caa8840c70359cda1033fa1927b92c692f6d6b824a06541363f6ee397031b6871bceecb269615dfff5a6cd9775f48267380ea3421b29111377f1fedbf949b7a7d80ff74b2d142dcf84a733730cf0f76c1c5fde1c391f77a9413a142ec7e541872e506a5f60a8a9075d99bdd65c1d61d37736195e809695ab6ccb76f0abdaca1aedf02a9bede02995196725f61e8184bb4dfdbd7d10b8b12a146862487884c564a32ec7a7dd9f36d60eb3eae3e7ba7eebe7db079039cb04e5419d84085ee364a7825cadfb163b42f884a2ca377640c174bbd910c81460b3063e3ee08aad073aaf31e23765b611ecca04771409f7cbfe4d6eba6b6118320c55e766ce919cf04d8987f272733aab4e1fe318b7889d6bd5a1838eb403d47b66ac7b2a54ea10d72bb7469a061642d404bb7e3672c9cfafa99cdd657ae469d748a1fae1e31b530393ac95b51de5954d210aebbfa543f7cae439c933b473aa39f125850ca1b97efffd7a921e7899a1e18d920e376ccf8b9ed61045c317ee1e02744c275cfe18c71f665a4ac0e2608bdca9b6ab83570b4fbd7f89e5c0fe1b51893ba9d67c5fbe6be3549c460e9a59d127410899a46de682511f07a0864d1e10a0ed611cb12e9f3f4cd2a987a48532298fd6683dfab2a5b09f6acf9b5524c9518d576f698426c87a02f386da29f509fc10d068dbefc68b5ebc158e3e280c260274229bd84218b90686fbaf8daf95078503dfa9c9963e59868cddaa4598a06fe7b0ab518a11c0bc3b1213c56b2e73d197970990018320896ec59d0142a910006137c1e2848876985a9525a1e4d06e6378972f42e875a89d957887855b128f6b882454e7c2b2b3a6019090cc4c433a49f9c736aaf0b29497290641a31c5fa34251eb1409426ff9f69bfbdcfc5af1eb96f4a49824b9aa159ce2463cc67c48c72929c66bdaee2405431c0190ceec494de2184e2b83cfc254b2260ebcc0bc2e68b811b997f7c107121a8a23eba3553753585d13f020540f1b0c6aaedab2ff188fc17ab6dfb4bffd7abe69f53463c6f9ef16243540af98efc3df4d7da1e20c06fa1a1495451248cec47dde0cc7e6962a903547737855a60f8a96459b91e3ec8d931a46247169e345a88a9a09f32063a0efd373fcc85fd6acb3aff3ca037626ef2553a78c58ffb9a20087d8ab89966995b719cc88d51e9bc04bcc5fbf35237a68aeeceb765e0cb113ca4a39604bd4a1125497b6643775397484de4591c5c6b1558c8f53d25caa052d94503e780c36220a59c7a9c68942c9313da3b4cb48512b59024f03df74158065d191cda051fad284da19b5e7f4e38bb129cec80076b2f977ea6c08a29122a61cc42b7073dc2eb7546952e801ad70a452d3f95d035b4cedb97f6c999aa0b417860392b0514555dcc4d8f293e22b666f9b698a53e6bc28c1e42421eea23553e5b7d688543e4ab7d7da57f389d0c7a4fd426ae83ec23618c9d61e02f2ac5e372e96bb215e89dc375d8fa9fae69d882766ff2a0510f50721062e784c086c7959d61c9e3893858515506141f4e7de364329d4eb2adbe6fdb5e482fe17cdf357c331dbb621f7284ef726983c0fce58e02a011cd162e9945d3812c698aa376fbc20bc9941e7c02cae2ba08d6b7e6e7ccace4e2917468e5800ea8ad0f84ec348c01d0532501d8ddc2c3b197dc1a23f2d652eced76db51e2df2d1ab44bb9ade8f9563338866d6b63a3acff4834f1af5bcb7792f8a6d7555ae450a25c9d80df4a7ac1635955f8e476deeb3faa882214a69bb6a329a1967d9a0316aff8f21ec9a2f12bdb718d232986fc1ef85e93027dc553390fe8b8d3a39d839b7b10f6dd55d6424971189554485aff66b243070ab43939178a7718dfe114818cd043e6cc22ac76306fad0ba83abaa7b7ea61905b5befa0f261;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hdfcf6f2787b116cfd653d2e8615ae7f08945c883f28dee64cb412890b25929a9953dc33f807f0d01b04e221714f0c6ef77f63bf3d3ad7f7507f8105b66f16d1723b02f138c57819b41d0d8f2d6bcc6fda43145b9b0ce440e4cc01f2104e581356a2e49258c9e9f81dc91d5e2214e6ccfba6cee8c5224f669b012f438759cac750bfcfb421452af325a5c2d47ff0347cd8e5d5c865b14505d2e7abae6ea80c1a92e26aa7a0744d2a8095317541f49e290f8cf2621cb2f13687eace8d4fe7a9c4034b3d5f161ae04558f4610c0333aff6f9201eea5ed657289165e4149eae4b6f52e008409b3a4a07f808ec83df53920373075162b46e320f1b17b85d28c1e6cfa7fa0569c79474fd3ca121ba3bcaa00ed6ca3b4fe208b697c3d1ba984938af2c4b473f9120bfdb2e34a95b956bb4c799f44b3d1372640467f35e7d65747102e3e9217b0d38a82fe4d1de0f7aa356bd70a94a2069bd04c1c806bced6f53f5f4ca0e5ce76a0b2221fe827ba549a4705f2660c2a9c6413b85f0c639a9e993de165f9328d419f725b56934c840488a3650248ad34d936d01519a74735045be62c3b311fef48685fcecb3ce12ae6a6c67abed9f8b3450fb08ae45dcfb285f4d7a3171e47f86b2cf7603762855771288042599599d8ae0db69ead75b871946a903e4c9d44b6a4d78ed59b6b20fb2629a0cf8068180e442ebd57a8d391dae9867109db771ed4bdfa64e97ad175995539a606c50e2428dc30c7f2d2daf06d30ba9376264c3ebef8a913cb078fe8f95949f9a2d5f039f7e2a5325bff0aac926ca31aa13c0469e9c3e576b0e69eeee0ee396c2f08793f4a64fc4d0da185f8ef4c4b43434676a9d88abb8fbcc465c1dc383197ab125640d57483a76366858cbdedf8ead0690ef5cbec40cbcf4d7d767d773a75a2b811c8e7e571ef55d380b2549cc8830a7f24074d6e92ba98e2fa8659fcb82bf412b949008db54db33b6dcafcadca0b605fe5443ee79e01726bf39659940930d35c7384d8041fb4b080d991b0e95bffe1250a7d084c4abfc3b1d6ffe931e21ddf80c88df9bb6130bdc481ac4007e5435847656531f62014f3822c7e1a79a629797e539dda60537da52b1a1c55371ccc9ae459e4832f2b633b04073c62b80ed8b1f880e642eb6547842e9f80939f472ced4a7793e946ad4f8873cd80b84a23f89b821f8164b6bf67970fdd457307c5960e51107798affb16f988148b027a85757796e2ee1f6477cb7b2f9047598b897619c19772e170ebca75b89c34165bd90f89073bff1f484153874627811df55d889ae428488a6ff8f753cdb355ee0a7d40fe430b504b87183fd3664ed82767e2eebbe43b3536b3f737f6219ffdc601a115ad3e85f702ccd9bde4e6629fbfbbdc55e482db75b874f1aa0fd01f77715a920b772dbbd904e3ecaa8b5748d5b7f10053c12301acfc25269d4834d6a561515f142fa2ae8eb3b6d4f4632064607ccabee3a3c62133cbed74f9701650da76352960f13498e4e66db9266d30ce1e603b16fa3503b3451592281fdc00e2c9208e253c5a1a94b5d893398823240ef15ef0ae4bcd320d7dda5881e86f96065b900650f9cff0c63a744ef21d126f9e3d4d60570052045c1ce109c874c0658b1b9843b94f158aa5ff9c2c995e138d0bc0689a8dfb60100b290b1eb249f81465e884d9a29c286bfa75990f5f87eb0fe4f226470ba06b889592c510b944c9061f8f4c42f884ec1fe8cc65be04d8413b60fb790d3eff20dd0c40130f898c877d98d5c04b431c213fb1fbb3bad70da2f0103b98016985697a92316d9e356110c6fcfa75df61d1b9cbb59f32669ade33ac9833fee0b52a4bf8d71698a2229f5e1b0080baaf9d4a5090b98b64b5bfa32e9f0a5e3ed41d831b01362473d0c9c0b34df6c7406fa9e43b5e7578330ce854b09764926c7607db6aa016af975c88f8d5cdb181bd07204a3725e8a3fce9e55f17c984de9561e0e9ba3089a61dfa217d963b3a25451cd9ec43c3fbe213cc9ab16b2cc2eab12347b01f2f92c1be0f00e7c804b9bd62b95e445614f09680ee217af5fa28662003502088ccc5976e147f7aab5f45e341f0372c4e57b25e2b865235038cd18e237bd3fccf89454b85c71a74375e57c8ef385f71dc2b2278ae6ac1e84e934a554f127e5ca9c377085d7a5ac898b5890b2cb249f07f24334d6f8c20fc2b9c8a131715c6986acdef3316fd34f63c82e8d3da7b77cf900f92095477b0296e1b2db313a6c039257f0f76546acd383d8ac63fc1aaab598769d9dd1c46255e0a7af6e9033f43f5b455efce6fdb81c3752642fad7461fad3815c4d116150e6de108ce884b4646122b7d8732214108720a5c6590d44398fe93d9f084c70c60ccd425b7fd2e33c59d673bdf2f9945a7c848583219ded371130bd8c2d78646d3bf02a465e15d166ef2d555fa3c50f234b9e9a63743c22174c00944b6d972eae2d7f148ddc38cce78e93ffaad4e3ad94e1525267820661ad66ac1d2b25caccf56a1090bcac88f94131186b8c767850e4728cd23018a18346be8852d4d99ac7e79c8e0473bb70c62e37b9b130201d15239bb44952f7d50dbe336e32b7b99787ed37a6a466202294eed000679f3bb1ecad78a0de863f98a0dac60b26ca28df3e47a3074d41ff37cab2a981abe72e12939eff6f1a45bc574b3b7c88b37502cf046bb49bbf136c69c82073e69608541dea19d9f84133a30d9fd97757073ada113fb45b616a6ca9fa737d177e406715c4fdcbac972debd6538136d46b10830518729cc632fad7a2d92d25dec9c4e10a7e82e8401797edf0e8471e89645c0a46d2265d909bcae2577be68cdb5764352c1468ffde5dcdeb8950b8ce99ac90558dca70eb8f41e143aed1b56f7aee2916d2d066b2cffcaaa5cae9399f9e896088a6088e7f9b3eb8fa61914700d5a55dc73b3571b48dab2130c3f196c29797d16c3304be6ab813491499a44ecf3da0b73470032ace6c1eb830bf3a2436c849bdb63ae349f2109a7c319e86354d744f769fb4455b481ebd0345d31bdb92570b39c12e1a5e26ef099d5d80beede6b5b9f0e08b80c2c4e1ce3d7179ecfb131781b90a522d6a27b37edaf14fa8148e8044fa2b2a8eb2d70bf6df71e85876ce19fbedc962873c0f39fcca9dcc26ff11e1658afac98aaacd9fb65a78c71594646695ff9d97b0dcb8207bb206c01cc2ce1c5dc6ea2147105d8ad715c1fe757a6e57659a316e6ecd27b6daad2bffa89c9b5cedf4982a851af5d198446cd067d789f164c4c2bc1b06d654acddfe06bcf0bb45e5727969fcc30bea85cc3879eeb11459ef48cd17c39e31919aa63ca39abfea0cfddcbc84b06eeadee2d5a156782a8813f45da32e42e05528f6087d532024155132b34aa5851492c600462d9c46540c8a7e8d1decaebd87684e9face8ef6555fd55b02ead544bebd1d29d2b7f663432a4ad81d63287b4201c6a0834b8c105cb6916c820c4118421228f52c25f6265b4334849c8b822c5bb84c86dcff649984c07aa34ca1758cbd295683c45503458eba62c69988bf008b68972031959e55c975b814671f30ea0301fbb7288206e31d49a8c2a1155443df58f1aa0465f60731649f59ede7c02884a556e40f8355b22a2f9bbe20d24f19d1915a809128e22ff40f1fda3666ccda6aa17a9a6bed404320732f8a653ddbfef59f964e6971c89c529f80be849e0bf826c3b3b1aaa7d7d3c82d3da1d459fd956b591255467d5151dcafd78e9f5ecddd45049c2fcd33d7a82d618d9c41bed50bba5fd128dd0c7bc57105d74974ede4faefcf7acb840eb4e00b091890eb816b5fc60bf8c1acb692f1e54c0875db769f79c7ad77cebfe964b367c5f0547a6882bc66ddf1124eb8cc1e84c2762bada2e60d27e9fbc892b1d1260d7b4ca0f3b0e83a7b52422b0838405f39cf860e896c1229e1c01e6565c2d559c5d9239059ccd3f8a0b181db3b70003cecada8177e8ed2ce67d2ddc20d2772157fe534601fe5163312a35eea6a564c1a290f6f43fc17e97eec7bfa096a9a7aa48d6b50765cc306e71a2018d6f43ac5b5de97f1cb3a3dbe40ea368cb703d6abfdfcc82047517e0f09358e75d1ede5ad02dbc0c3251134ad6ff69bec4323d8b21ce42dc2d2d612f1ecb5aef8e608ae979bb4eb500e0651a80f232d5e0f0268cef0fc0f3a4563eca8b9fed1c85a53732c69ae32956a58f6afc57beb60ebaa966b389f60aa3671198cc0ab705b67ee879655b9ef22994efd15315ba6a6d198298eaccaf13e02eacd7c416e82f334b598415849ea66d4fc60652c1321e10fd58787c2e0e2d250df6bcf678f2827dd0eb500984ca3a71519381dbf5b29a4c2919104c43ee29cf4a61f67a86e90a269035cc60e4a074c11a4b55c6551d9186cbc36938f37530d17099348586c3623b1818eed62a6ba8877aaa087f191165e8a47fb73e66d9f92a264d24d8680a8af3d6c29f8d59e69cf3826a05f755d2e7567dde9a6df4db640edfedc2c566c2612de8bcfff61ad147eefa468a800569a84ca9076a313a15fe9b5e9287bd39db87cd700e48eb7dc8f67e123eface4df71d31aa51b0c30ccc9be309c3a8894616ab3f2e6d892d13d1a1bff4f9ce8d9afb41aae45efb8bbbfba99a8b22c9fbd8298734162106ca385c92878769aeb77fd381b664cbf5529c560f9f6901a7a00a32fe39e7c3aab85606236064347b34144f23d9a093eb82c094f69f2b6748a5363e5fc339fce645feebc444c7eac822cd82569baa4f4f6ad0e275fe6e0c7311792072332e405971f48be65d13719f59669505c120bba7a31936db86ab85fa1c541f531215212e95806a5014e2f611239bfdbbae538565728fc6c61b7351ce19189b1fbdb8361cad9318103bec7155f6ba193f81321a00109c3f5909c1f7cfbd515081c3fbfb413df0574f569ee93fb15cbf3d4f36f916d268357b6b9eaca7d58e44546b22152ce35ef2dff34169cd380d778b19382752da97d50bb1ca0346c2a8432c8380e0fddfa57b95ddbfdc3ecdd526623e086e1ab2fd8f1990656aed3a0e33f7cfc10a02fa46607047ff63db58c5eea76ba9e61d90f34913dfa8cedeaf5e3688e8124df7ffabfc6a5291b63913ee4c56f470251879967ee58f43adb691d5b3a7761420d0e67feb3b0548fab02320dde12414b96a12bde9b14684db8fbff765a5ac4d8cc8d1de22cb0e47c6037f615aa4215d598cb68ce6c25cb3d99c644a7ebef49d9b5f1ae6a6e4ed2253dd2bc113fc59ec943eef5e0962adfba805a59a7df764dcd12433035d0d6705ae991b8f401717b7ac4429012e53a0de7aa37bd5e04b9f3313c1447d58508c31138b01dd5f85805603471047ff5b2fef942504c15bca99c4879c53d0f44a2d4e84fdb23e2b8f047c4bbf76212880af74397c4d91ac05e64e196304378c3c3a69fde766434bc9f5ca321628585e1985a0d74e878d4157a676d349326cfb0b301d61a2b627ad1b2056bb5467fe37b2c4eb5dfd4c08b20bfea6b28eb6cbe947efd3102e3d9fb49c838bbab6fc2033a36011cbac88a4c88f382440568c21a65cd43985694bfff16b0040a5eafb60921e4c4e44dfe8d1442a2689c977dc515ef30b107a245cb3b8cbedf7ff1807f11e4d8caae51669aee6652bc5228fa74f141f8c75d1d369bcc0b44ba411dff968f8b774faa6c52a460c3cedd4696583b2851f832493c26c326d05d6f910b34b458900d6a598309e052420e999583bdb4ed81c48a2a156892a19f7390a4491584b5d32861ced329f95006d5479021a2297f51fb8133a3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcc1d7ef4c27dffd51b7fe049b128ee82c6de1bc14931d58c48cb7502c8a352d6706916e808f15fe3a03703027afd46210a6103d1cca509771e75738a1349d00aa72f3b0deffddb899a519b83857031403d8d406a50e1f15eb16a43d8ac376fb65f6efb7020be128aba8589d807cbc6bc0169b966131ffc731d135497eb35ff9fdb72387f27de8a142dbc4f94b2be9e4bf096c43861fce05b3b6f6a5c2f19b5d43a3d8dfb7b923930deb83f18221427273bcb2620724f413b828798a86834caffce9fa0beb529e758ec2ee4c555ce59f17bc108245618bf84dc156142a40daa883d646e24717456feaa2fc1744c961986b9d4b5c5441ab68e7b1d85877d945cf271dd9b378f95ec46864c906d9137c2f7b3400fcc32f59c981ff7d46e53894d11fd623224d30e393181f79c7bd0b4d4ed1e57ef5384cd7037110c176c7ece2c640ed5d6a651f7cffcdc338570ef387f63b5d026eb3e3dbf0033098f7dfa0c18d5f759d5ac60089ca80ffe53b093c00bf4494d82d3b404fc692a44421a2e42089cd9ea20c3b70d8a2d3787a39a328d48a1f774da0af1eadc528b67cefd823d1a1da227c614646ddab8b4454f87211acac42990b82b2fda25f9bf5de0743b657d1b2d76ec29d01090db3f25fc0fd9c5abb9e7dac074280959597e2f0fd7d45fd51682bb4503187aa0876f9f0d4d68ed23d72a4f8ad095e48d3899e22ace5a9f1feaa60de6bc72488efe30c48f4f6f54941830112b7402b8108ce65bd61c2263d72c649fc81354c9af2ebbbfe3d7031fcaeb99017a460e2c5f691646a712eea55883c5d14451df3483f5f1cf7f97a9dc56170a03e70ce4e04ce895c60ac6040332487013e259c53d3a8ecf9ed211563f5acddf4999f524c9b0506cfa8524142d9f042370a1478ccfa9b6a20b826fb30c2d0c68d754a6b7d6bcc7fc3c1dd5da30b9c9ca3a5700003b7c920722857abd75d8e8ade48dda530b85428a72bddc5aaf95fd11bbe01f86bcc379b4eb0e50cfe953581b0135aa94873f9f63cc5ea92857104ae4ca1c302074521a0a1054bfd4077d617fb0fdb356ec28c990af4835a0c46299f87a37009749ade74b5e35b11ca5008a353518d148b13b181588f5915b5f4a762fac65c20c7a51c7591976cba522549f09a413e2b4c46c4592f006d5376345a7f5209dbaa5395a402ebc8bb3662a62486ed7306ed398f72b94ce45f46d1a88e397a397eed83495c1ad02ecf949f12f21fd328ad2f752b0f250df4e62d786d32b8ea147c9fc838e93c5ef1b7f74a3109e8602093d74dac8b91d7e40f3fa0625d7bfd11accedbe73a330718f2b49b383e3f11ac8203f55c87614bca80db14d6ad37a8a31ef9027a794c428d5e2a878b774809217d6c46a17da311081eb4f64d76a72eb4582979f319ece3b03a16764cf3d3c13fdaa5d95c510522430459ffdef8edd9649061101a6af13318efee9331af68bcf1550b5647db517543dddd8d1c2ace90b71a9aa3693778b091f9b019422b396c702608a38321947403674dc10abe4f8d50a7ef95cb420036d9188643f140803957fe1de3b03bfce1092a9ffab0eb25d3f496e40e00821c631e53dd54ea1b828a35e1471b487464c3a35955487631b07b14f563312e596ccf9f085c5f094282fc8da5b6fc785111c0fb2ea8b14dc9860b8d844a6b0e8dad582b6b56d01e2676a9bdb5706dde24f7e1fe2cfd2594b9f67f7354d9991124981aee8200f3b127d113597c3f72b78e91bd3ef06c0a966db0018a7416bbe422c758a94ae6576d972989fa5785f42bed2125f60ed164b119ffa40a0d678a75141ba5cc8dea9a171067025ab41c31dc67b2d9d5eec2889692af744d3f5ef43adbee419953357c555e980c83d7ce1c0079cb7bdb182317af1cfc7bc82c0dff09a0a714817dfd7072bf0946bc377db3cec7b65609f5582a02d289e929b0f7e48ee4a1877b0b609fd94cbe72da145d8924642a997230c07c2e24ed5ca8ccb56ec361e77fbe2bb78427c39b8f9663bf77173c472bd125520428055bb2b5789ce23712cc604474432a9738470c014c5ec4f6baf63c8c5aea572f25f0fbb646d4ef6e30c32903b272ea42409cf8eb05e89ee1e5eb32a30495568c67e60fa7cb9929b9ceaefdda22a0ebcaa0b3241cdee9c3150421a06e57bcfd76bb841da9c438ac82feac10e102152561039e45e17730b3e0cb56f20a08c8a33ee103e72eaa748b27773272b9b3f4ab7d5035e587acbb3feff60dc0cde65a70b2bd4fe1fa870a4748dfa04ba89e68ca1e8b11322b0c5058aa80a5ad673ccdfac9c30e2cd0012d20e0168309ae519c4e5d1c4bbacfc23e3df948cb9488db39b598decbe9f168901e8451a39a1cc20f231d6f148315e0b27781cf2371fe21e88daaba42075d4075f595db625384628ec80b233f5a4ed704d052c0e1a2df86ebda32d1be3c4f73e321c5f03a1925a00dc6da61e26a6544c18201ac5ca3fadcd5c9bd72f25cf8263f9a493ea4be863ad9eac9094ec1a6161a50c2607ae8b6cc66e7833501500116e98a62a13f7a9d731141a24b771f37b8b1a9e721afedaa15fb73b489e2f474d2acbcbe6a3151e423c8e4268034805e26e4c9db4dcbd59ebf1d5a4cbb980943ba9852be5a27706f5f8b5f110e35e103af36a73f162507f901ae5290c66db0d64f5897c0ba454ac047385b14613424a65a20f6ab7aa0856453cc436ce8425571e8d14b481c08cc532e36b727d16ff5af2954b16f695279f0c776b68e6af4726154343e0785e63be64131bb72f45327201d25f764f91a4387b6c0ae51e48b5d6d4fc6461db92cb57d10433ee53be73bc6062e5577c87c139608f0d1b48dade192baa393cec9b9754b0e49090601dbbea2894065ab64ac1dbc5c3e06017ec57b6a064aba87c394515ed7fe84bc153e45fd3da99cab4dec7d8fac9e618f8ad37e173b9b84e86b8ffea01e8d21bec30efd414dab51626204f24369bc8d4420b20a728f20cf06b6d37aaa78afc4bc39f058cd63931e8a2e7928db9378b92f2cc457710c6485e55154c23dc7c5fda6b5a9dbc3c0de1302499584cbf355259498db71e8a94c22a16e036759377470bd2ab7b8654c9b2ac576dcb69dbbd76f4a2745d33e16807d03a8974a28e516caa407d3fe990a552df7c70a9daef83a6565024386ec57545bc35a16d5ee40d6bf19a924d91a825ceacaa1d8dc329d457910c725fc361e7f3c8956ffc2a1afe6b275281b50b3d04ff17d4d06b81cb9683a7c49e534df383fafd1405d8b79fc6f6a1c7feb884f58a0820a2e7d9349b8bccf73b4db5523657d7ff0176a7830b0a1b7e529f7728d8132d42eae34d3e015d051666e7523d4e3b2f4b1a4cd72d2812620e2e4dce199ff128485455fdfd6bbbb1bb08a96f287c7ec6a4d4e99c3ad3d90c43c4d91a8cbe1c652882d94a96dbf5435dce2042ffd179a3dac4a331873190aed5d04e2576cdfbadaf62f315629f516517d32b8fbc70981e1a039ec40edf5b167bf7212e8f2e72fbd15ae23c8b58a8b75b0fce0409bd6da051b4b4760e14d9c180722015ad189b0b65c63259befbeea729e630747b776cf2ad4d72afbb78965867b398387fd4abed383d493d153cb77500c98a296c464020e56c16d7e05e8d21dda582d17f16e3dd14bb32b8cb3488070ddd4efb5206d1d6afb42165ad5cee6b9431fe379553ca0859d86e701ce2c7a13aedfdc10718404276abb3ad2eb50153ed6f6327b64660dd7b74a489afeffd1721e48cbd2aaec15d8086a3c9aa2066fdc1659532c6bcf66d3f66217722bf0b60ac5d85724f64bf4422dee53607fd5e60acdf33424e38c61bf0c0405b95e1820bc418ce29934f49e4f16b87013060bd3c8d5e3723928b938c8bb69445c73929ef2a6f63da176382772c59f7c1452665082d7908d2045f9ecf5e771d3ab2fb72d0ca6416395a76c2d1f9121080b9f02d2dc76fef92406ff837fb226820fd67076dd93236444a0a8d077c57722d6d8ae55e5fa4580142e7c08823ec71dc37f2b8e5eeb8d1de1d2affd1226cc10b20ee3430326f05b782993d2da704bc662e7193e6a7921457a5f5b6f651ac88ac5b629631715e6327a37e62db91ebe273df12b9e5d6066c7ac3ca6a3b50cea19f639215f6691bb462c902f22c5d7d2fe6a4023701f45065e0036cf6444031f4e2ca4eb9f9c3d4f5aa1305e54f18335ce91a3d93e87145afa658c6b82bd56c7e1a14660efcb681d77cb7a74f55fad8586eb1ffbc9ce96f97ca180c47ad3dd30273a6ce94ed53d43ebcc61cf3d52c268501d8c087a7076f74d1af383871e5a7f0fc0d0271b963a1d3f8dea9742a85ffd6ada2ab3a4f8dc4fa336701c0eda6856ab0f9edeb45aed43bd341a6ecb0d61bd07dba3857c07185fd6d77b5a278178b757fbc9d8c1e4781c43290b50a5dd01062ffaba2b1814caaafda207dd8d4dd6f1921f7766b88f0ceb0c7b0507f4dd89d7c8d62a8382e9c0cf42f5669d63d976b2cdc833a9512dc1fce9daed88567192e9b54c3fb1f545ca246b4e6db0ece9125212ce45b0e309b0cc5a7dd95daf134eaae8ceba57b66728a711a883fae6248cf80593fc0cc8ce53361d9ee6642a817616b517c868c5cd251e13ff7b5186722375cd80b9c77413241c2c40492cf29116c62e04c5c1c29849d0635fdc87e53990af0f2aa6bdd3f12d034a39b0e9057349f965beb9a5e46cf624e0f7356195dbd7f4c3d4f46d2274c6f64e522f1f27c36a6172ec73cd4ff21ef28d9548d911881eeda9058696412360dbfdae90c2b4a6855c583caa951f4850592a0a5c420a32aacb8ee2dc6b4c74da01a887b74f6b2a772538a1f50ce7d9cc9b0558547a6b547cfdafb9cbcb78289e4dd21191b18e9102351a32f4cb9e643ad275645a2455a47792fa890f3faa98f964dcab82942d6ad2d03acec887f11b5d8f064b1712c4079c321c40e388a307bd6c2590db4984d91f2a7b114df105fe36eb93b291a81388fd375129507638bea04c4f7259416d4d15d7bfd782c0400da07316eedc2d3655a427c979f171d24933cf65454bebb6e8e98ec5d7a58bdba48f20feceb2c4f56f1bd3fbb1a57cb499380c66ce8d28140238d689e57864722e5479a2125a4b4eb9d762e8f14bb794eaa2cbb8362df9c7fbfd46c2f927cf7e6f84ada22f3771052b42502634d4c97eaa2992d941aa657fc9447202c334092981acf3ffa613bab2939abaf979f6c0dd0211c17af270e0e3217bfb7986f6548cb5248bdf6c9085ca5ba364372eba77553bb5230a2177ae6c498ffd50f2252d1aaac956e4c33d6dc73adafd934c856200599fdee102cc9a9271dfef4cb58278aacbb596387066b41249c5aab17ca8bf3029573b472508525941b6978c3f7219e6a9ce0d3ef849883829b5bc3d1f756a7e0c68a4eeedc33a0d0a1666ebf21024dafcdefe31e4419ffa0e0d4dca1eb73c2104f80e589ee3b2ec964fdf8f9741eb57d2af61ef45e07b9332d6e258b090c55fd4bdc320bf91e1387c156c47fdd39cfe4afb667ebefc06621ac1d3f69c08dbd84cc50d97e9c2e10bd76a83aabda373a085cdb1133dffb8c692c25357e06fd78a20a25ad584f69107f0144c5004234b78e112b0d59986deaf9674ec21375f187d8410265f5bbf8de50ffa43891021827f9ba51e1b44b3ce793a46a7568742b7472a02aba69029cc2702228569e8854da0a64270516236c743f8b4505be4a50cb001ea1815f3b47c75e4d31aad9fdd0e4a1e1e4632264038528b4e779508e77f9bf9270ef063d4d7ca69c00aa8bb11fe643f98890;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha7230475ee308fdb10b82914dd10ccfd616c7849e8940d19574baf9a6b916aa89941693a8a13e797f2939e973a01d5f3b8f4f7f18cb97fffe640c1fff293e8007d6a68e0fb4a0b4653d9240c5637c03a8eca9e865b261dcdf96ee9a3d00b4addad3f8f2b5fba1c29ce96721ccc6ec3c0e67249e4bd93c21df23e1f52330f7700f6746b83d9e13e7ee50b96799525b3e7b0bd3a297556cfaab957b09c26f24d83cbbfa9d9d100ffe9c85e4449fc4aa725d177d3c45673ed96440b60c52c928b0c577eaf93c656a9572aae13c28b05d60fbbf0d7f02c0fea16fd1269f5069440e2ecf4356d80b403c014bc867db24d6b1b2aa7e52099adc24085783ab87d1a55e5a8c112a812b872a2da87443f78b07f4b828a5cc6a37c412e7b5aac8aeeacfb2d6c56d5d14f96acfec38aff0bf50e64ed1fdd17f97bd2390d906faa5f6cc8e34309b193ea9306fc0f57c964182e4d91c6c1058aa52af6f10052e4bdb826ecb0365d4401098abed381c654530bfcb6e2167c1c441e1e38c00b0cedd2e172f17b8365884db4140c16001d6db06141cf48a6033d9ab0272c909fdcf6f2af79cd9d138ac7873004115dfc0587f8573a62e72e9d689dca4ca2b1df5f503d1118c0c3855f065a602e2070ebde9f4aa85c7b11b832424758a1263ed9cab43a9d678fc92e6cd16702060760e610db41cc66be7f778cbf1353e1593b67debd9d15337156dd96123452baa50d1c202aa96a4b38bf6e59ad6fa1829e82d3f7e03c4d07dc01a5b6e62598d52aedd362e8197fad4b66d013af036ccf792c7d1dec5054ee58e106927b3b78b86050645de55a40a47f3b2f45dbcfd1aa9718a6bcbf6d0c611a2722330b4b5e2e22a5eca5fd4b8983883e4ddd31f9920233a91a430a87573f9329e03ab7fcb5d1c0cc96b96a1ccee53de23f9fa0ccd955c8ef2f08bbf129e40dfc08d9b2ef751895fd09845f29c5b27ab7b6ef077b78bb8a8669fbb8e817ddf5227ea69071924bbc7d58a33e8c352e07f04a370f8a3c5734e52ef614af2b9496d5c125f0f6a3d59f4bd2306eab6964418adef2ba54ee9621be6ebe5814ddc92f412593fbd74253195c8e00803fc031e76d85039043253065fd35fbd93e6efad9d304c7a1c4b9074dd6a11970214ab0ed2ada0332a5df3882e4f894ce2e4c677c6b0e7448b9c7e3acfea53b43137e1dc6f552b34620391a26aeba2be2debd6c0f6d9fc4b4a901545bfefa2f2f3b3204e54b48e053926cab895df7444f8cbbebb1c4e97ebb2f1c562d121a82dd22d3448825b732a539c4d20897362fdaed93432e1252963e2bac2cd8feb6884f57713c835206e767fd9824a635d84e567dcaf9ca00f2c2c30b434f9c1510e4fa32ead93039b72327d23449902719bcb8595d258f4553bcc61f8909f70d7dda63d174743c63b52a7f992b6d7a414762d631103f80a8a336d63a324af5900d717f1aaae597c5dbd268829e5e4d4d52806bb7553f1fe43a2783b0b68569ae3eadbc9c6e7b7ea25403b661762461ac93b5aa378fb1faf69f53b15df48fecfd0870066a8489ccc7533b1c565afcdfde440b5b5bbfbcc88fc7a8b5d72953bc54adcb4826960450fbcdd76fa6662b98ce9f8560659a2664cd170e75f9e23b410602937800c61dae3d536c4cf829acdbbce2f4d9b8abf11637ddbff148c9c0feae459d830630964976f6644d8538c7ad71a366cab0cdeb17978fb070aeb61311f6cb3b8e5783e8da41a98ff7c88d670cde5f92a384a5675b66b1a925c7063de36fcc398491f72d95a0907e10d1e724d213c7882724b413075cc2a8a287336e965ca6fab74833ddfb2b3e1213044632058c940ce8cb8d05c0c578d1c94b8c725e6c951f8931a3d3af767bf18d72ba180c0529140d7a47cd46cce97a341e0db1593fb7578a0e262649c07e39e650a62b6d13abcb490e6606289125adeac10abfff14f701209ac1d223f8278d10764e1f9b5a0cf559b2bd9f1637ef6e8f12f2c538d678c9f2f656a2c4057b59c91061c0cdecaf81f92b478cc322b196bd525f6b4b2e61f4369cff846ef41ecfe6ff01126e5d5addf8a62cefe2502285f26abc6e93515aa0d7baa56713ff2710fd85a046865fde872b9a7d7ae0529e723653374b06ea74ae74550c43ea1eee5daae0003f5e156d991548c6641fac75aad6f51a6988082050e17632995af9c1db947c6ef606219083863d148acf607ee1e46ef56f422f6f97613c92bb789eebd44da256bea7ed44eecebc7bf25128d311158ae22803acf2e2894042c8eaa543ed4de292bc46980a2f329f61a53f4eadb63381c528f9be4da8e340aba9901f2aeb9cff220f520b124e7cebf42342b12c8fdc5eb5e34c2946a0de0cec8b1f9b530cc9020d1e631cb874e32eaf5ab1a0abd9ffa18038c58cc2e64eecdc091a78e3075e8e22ff51452cdbc3d589c15c83cfa03d36c3eeb073d7aab32f6709ec716c5e885f6590f194f1cab4fe5ac40693b726040ea8d2c24a5460d8eae4de6240e07d5fe054747b397036599283d7f63dbcfeea6a9e12292c99f34179a0f30b2185f8c2a35678e29e032a4f912e3a5aa1d992f0be99f5ead0567d8d44749b598e22277eb2fa426eb33c89b056e85bf3c30458dc2a352506d3d147984e5095724e29eebfe683c24e4c677546c1c7d73264bd7fbe3eb56c31c44839cf05c9b75c840d9ddcd6d55ebe3c689c7d4acb9ce75451732b21d2fd1a1ad3159929c4c95b48e0ffbfa98b8751bd58279833a1fac1b128f6a1ad02f4017416ac02d49d99c79baf97923fae81b2737f06334f8124c018d29dd32f0cff39aec7b40c67e4853d9533e0408ccf530150911ea47be0a3f439d6a7bb17bf910849f7419606795b4744f932105954c5d93514e760b7094aa797829004bd4c236fd8fb1c6ba218571b86e1211d2d5f18068fe4789f941c30f265ff3a45e2815873b29c9251af09f8ab2bb8ce3c252b0e93b9c5f631ce14dad3b0bce81c9c10913099b14511f317d78030cc4f6a23f7f3ade38f25087673313f657e86a5010cbbb9323af0679032ca5d7a186e7074d14d99d5ec1527589d646f5fe4f5d39d3f41a82b0d5d4740bc9bea820c4b3fb23e06b29f80fa35c01b600a9eb2cecb55e2e314c7811c35954cf332dd2af7bdb542854f8ee15a830223a5e521c30b20e23c416f972d5ffa5311385ed08432e1ef9fb4182ee0bcf2a3cb9fbc2ffed1bcf424be9a1e0f4dbbfe7633134cdebe12a218a0a55516014dc8c8679ed8235c4e518910be8350f29433af7052294b41238816d24cc9b1b6326043ac911ea2946fbf94cfb43303ad8b4085e0807f411fa80abc12640c0ea098308168ae17456d8d373a4d5d55ecc9f2ffb6883175779465361903391a4388df2afee3ed6799ff391ef3735e426ef0d7c67a280575c2c5b2edee51d7dd97a89eb87631c76ab87d2c539056de1db46045b6711487dca9844d89a6bb25217671e3e7fa9f5fbe2beb4150dac13ac5beb4b0c64b81cd5236402e766e698201bbe3c56edb784a04423d6537acc89cc628bb6baef0cf7afdc808faeb81906e738bc2a610f5f93f3145554d2665de9aabb0d73014870655870db7d2c13121360e6e9197ea0496541417dbd462b5b654251a3ac8eaa849abf0e3b1ece382942f6c7a4103912646097ebf3349cfb59d2fd318ea2ff2f6403f05f86e2237e6102bafd0b17187a2c0b7c56d29d217e223507a33045c63d50248e377a456d74744e01b6289549d3ac22a46f0a4a82cdcef58ae6f7ac3c914dad5575630b77c0916eb6bd22f81cf3b017cd6871b0b5dfd90ddce82a3ec3327b01b8566d7e09c5b482d2ffe467e381867169ac4be707c2f9b92033360a337af5d24c2c691a44840c7322725f199b9032f29cd994858696949d39261f8f90d4b33e77812f8b980b57ec906ed0a7d13b28dccdb207c866941a97c770e9b7996fdff0666db5614efb1fff16ff8602dcba807cc2fd2c97b8cb0fd0a423cc1077fe2636b90dcdf078b36779fbf0c573ac2f8d60b67d831f4bbe79f175d8dbd96797adc682baf084a4daf55d80256860c23c11ca40484315909c7278dafae06fa20e85d8b3b9fa3062c0727c29142907def5d7a7541bf1d1fe1972cdc841ca82e967dacb3ea6f0a68d6e6e185093ae2b616ddb757eccee903aaaa8a4e11ecb90648e4bff019a0c9bd2b2e51fa4a8f6c5ecf9fe75941e46161fa108827613ae52d58ac8fd752cbbdfc5bbffeb54fa6038d9734d194545d2349820cb8e62d403e8c3882db856e6453e45ce2a17040500f12839751f2ed27690cd381d90c86cab6234428b1d54edc679052a3f79d34563e1e9f063e861f39633ae71bb4630a066d1b4b484da737ea8caae15813a680d6ba5cdc7d0e797b9dd04e8c0f282ab213a256e0cd28c7367a06953745f493650b5519f449cd2063d7ea15b75f16cb3aabc4e3bdb36bb3b195ca0a5933a40c7de13cba15bf49f8e826d7ff673e9a6f09e5492ccb0a454121bf7ab119e7fdd85460fda9e43e93c812fe7f95010926604fdb801c9c4ae6dd608d90043755127210a788de86ca1401812269d07f871efa8b44f52da812534a6cb97cdf727f5bb1fa43c866acf2b373f31e586277f676b294ad779652b242925a3bf082a286c100bc852a3561e57a9492dfbe03fe1c18ef3475902577b8b1a169ec8c4bdbbbfa0bdb990f139462260f6407582661899a24fcdd7827d033e34c5d7c7f3f5b7af4162ad5bf420e5f973ec874edd279aa216e32f4d98a9f3808409cf0c136c52f31803f84e751be3e37334435c7fa14829a169aa974000843a11a5d909d0045e350accb380bff58f0348e709e1fc8bb39a797c5ee8c14d241ef534234f1c12d044d4b31cc7f218c365f97577b762e92af7bebb32804314ed68377bfc539da85b965169bb9733d7ac8a8677add7e7140d8c921011e628c54fea71d30fe55565ad6b7cc051279f368be3c7947eeba90d70c1c26a9698bc7d6822e6ee022181779d33e5d6aa499890d309237c60f171a6608ddcc8e4404b96622300015f25e345c78582be9d2bc186e98172d9f037fc3803a39d9d84c520dcfd0d692144927cf95364ddea24eec553fc7692a0f809ce9fd8c073003807e08ff9248d6ad19c7cbd88918beaef893d50c7fb0a0a6195dc2866536552fee3281efa633a1601a7d4c28dbbb4f967ba30fa9481706c30ed08bff9e5016f0f5882af8600409f5d63dd91849b655e503942341290650ef0a3012c9533bf461e6f2ae9f76bd51ea5702bb775dc4dd11859825c8100432e91e00ee66c95366bee1a3c165b2f744d77b777fd0af6174b9685bdae3ab481c685c218256971829656e0aef151744356f683d390245e0b947dbe4d53f35f80879a035deb4bb0e4f43756d69476feba1363d43806e4f1db7c5097c6cd9a6735333f2f6e47da7da9147f35d1b65e23dee68e7a96d23ac0e3e80348bc0ea9e133a5909fcefc292a7ca370c8ac81ada02e080b6bc4d0ae08839c03547f76c2f079073f8bf5eb98625407340ed0c7ac8d810402e42c20f96bcef08866745cc8ff32d2f7b56d164ec2af2dae4285c50400f2471f62e091b209e74825ceef2040e87ab408fae05016e8f51aa6f5c0482c7f8e9fa41fbafc1fdc4369202cbd7b727ef8aa2917acee55c2f16f5b12e8a91bae6ae5a7f5e305a4ef64513031fb623c91e74a8d3cbde570adfdbbe8fb06196a079454bbf4434663bcd2e01d316d1fc616b4d79d38b965d51de1623267d362be139db855c99f9ca4efff1f8e0684ab8dbb1a9ff1b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h48b4e207f5975781cb8046c8891b963a0a2a221c30c1cf6156c6fa76c2f36765cfda88de2cb72645d9bef84d4d856cbad71b3072846f51d68dfb053b6e4f3fac957b935b4d259a5f23d12ee958eb2939ab9f625525c472936c40a57c61b6336b456acfc6c3375b17bbae91e415f5e07b5c085428b225c69fcc8176c3ea8949de7eab69c1d27091acbb0f439da3487c1fd912ed1718d29905c343dbb986fcb8bf408b2f42dcf621a21fa459befdccd0e42e5d53fcc7b17b2f713073d51a4c36147c726efec890d891c1c2c4c78bf6178d22ee79645b069960c6f47fef7c9278f4972bc294f3b2fcaeda8212a3fbfe3123db176f2dd2b0936f2152f245868428ce57d9afe292b9aa94ac0a5c7f0cab7c03742a7432c4f6868f4a25057d05a2242634fe4e450481e3c61ff0689387469f3374cb8b3fab388e7503ec087c1db1e9e76b1025e95953b5c079fa0581ec76405b89dc46084f236a9ee0835360fb5ab6ccebc046f652ddb2ee01d28c1a37c67f2be91140dcb64322046ee10db80cb6e1f9e39a994460d8191c3d5727c34dba6b40fb57b616fa1f8b14787d832155105874d65f8bd55d3a70eb69687a1d60863bf6bb5a58719249729518953c56c82fb64e942798bc4e4888eee2a7df3fe11419076b2fe5501d47e1d5149976b3360e1ef5a3417cf0190bf98dba4bab2e704c7e83f8da601978df743731620c7ff5c072840fb6a47af2271ec9cc6c0847de868814fff14c3a935d131206ac8ea48e35c38a0213b9ffad8558e21f48775100730e815b626ada4dc6f20a771879ba2bb7a340a0e4afe051673046d2632ce3a429e67499251a61f6fc37d6eac4468d66665836bce9a0aabcb7971ded00e94f95c1aff6753cb6af0f961dc496a2f03b3b5442e829773a32cbab0425a610b5896cd91689583de6e376e2cb693c635232127b1b67edcaf38644e482d28680f18d2cfd6ed1e4400d56eb3d14b530efe407d1491a156243408cd154beeb7440a5acda5caff84da94c77c870623a548393c9ff82ed7f804a714399a649b8c2b6632aa7fd561fca35fb1133a446caaa3a6a2ad024bec80b34a4c696e998329f9ec3b28032f04dd02ec8d22fbfb60ae42473eca4487c461357078b0df32c65b1b88881266c3508608ac1873a0211426a4485a90efa5538a51e4214c41008833167bc303060511f0538e49ee1f3b4f3307bf706ad99786f31efec6b354a5d89716056d3a789b5100d10918c32157b3238dfe74355bb47bfac9b7313562461a2b9dedf2766f9320af83de3f3ab99223216bcef2305d8ad63a9176f5d55b629226b976106b5f57ea49999fb0b8d1395dfa195d934a67252a07de747f543b8b045072427bd13c6d07fb049ecde46633b6f2bf901a9b8afc2a86a6162e75fdb25bebcd891ef0e21b8afa4de281718499ca16893b315157fee2b718b5c8448d89850fe9bdba0a8348e8dd98f1a238cc04054e7b5f65f23a8d6251b15ba30600d6eb3c7914203f2de1dae742a5e20fa4401a956b7de9c8221cd0c6ba79dbaba99f23b5b4d073faad0cc5019af80d38505f1b3607a4ecf68fb8ecde052151e19d6a96f557f91f348520a58b6fd4f1b1b5b5476dc93d2eff39bc445bc73e9cea0d1ae87119224f8dc6cd86b4973c76a2969c501703dcdef3b8300253648dec3714f48a9cf4fdc8f5d8eeaef0124f4e52a6dec5a0ce743a46878f7fbc4a21ffd35699e200505ab603da22b08dcf562a6872c83b50178904dcfe987aa767a5a37c419b921ffff653c59c58fa69f4d06f81a9dba2675d6f40810b432527d7c604fcdd3a25d563400c62440efcc4410300967fac6fed265c35c779eb456547f006f6f757275997bb5b564d387adcc7033a1c0c891829edca9ff2ccf4e4efa15dc3b338a60bcdc60b9418a859d4e3578992be4b6b173bb65030d48b9d7aa9e0db6f2350219ae3a840ea472c3db229a957054d7bc792d661eee58ac369a1e837d101c8f3975df46d9fb858e6529fac835f8734c4e20bc0668b39071817eff71f340139e659623926f7d77b69c392a4c982db2266cdf71ca277571e19164b64e0b1c56ed7af60d22e693defde450c6e0abaf29f0488cc98014002727cd3c77b040a7143c556aaa5ed8900ecba184d1c8be8bab98119ee7f2e658259428e5d29087577aa049b97f38d89e3288f58e41a91d41591616f5b47ade3fffdedf819574d23a7a44501dbcde1d1300f6201a7ecb16f47d8f246332d90ace4e60b37bd635d4d54105410bb353297405c410e9e63832e8abbed9c5508b2661fe2e6f6770397e6686639308b35cb81a79298dc21f411257da99338f6c1076d4e607336e5918a6188afd5feb33dab530d0d333f722d59b740fa814dddbf6222c1adb3499824dc13c590a1da88ff5879599da11ab4a49dcfe1cbdc815a6c4ff09a77040164a460ec3e8bc70a12f4ea3fc15720fad73931b62e12c413edb9722a6b11ae50842af75cccf4311ed0792a785fe553869a4430fabd6c52422cc8aa896006ca18a3cd6298aef49d1e911ba60f22a1504553a0d5c0e70f8d7630423b91bc8dde845c6ef5f14f541b62a957cb9b36a529a53845e05d2d1cf12f48e0a709bc41ee4ae4e3660f271778bae5fc6f92be0ddbc45f63bd7a921cedb8a955077686ae5cfb32c4d188164e09c91041954ed87326f6ca6e5ee7412a0b77c42490f3c073c30a85dc3dc74cf4ddcd0e913f1c90b07158bf826f10b469ce13c523b2b5febdd4a02dfc9c3b726edd3d3e53e259213eb43fcc0651dc69bf60e2b55b90fe5b69730106f5fb09aea924a1af0fda1ba235fa0f0c248fcc1ede3ae3ec60f67a627913b1ecb02642bd4e88f0f2dad53b4c89f681f438bc64bb1f320e56405419c2d342709b2d191430c926ddf4150c744f0b26bc8896c446d52727d72c3df925090f12183cbbc8d13594f9aad2ab6171a93a79849e291b4202669b72a6acae57c6a708572b2c331a7ca3bd879597b2c4fc3d89aecee48e1c96eff6770e24dd846791c4dec02b8e967651b94a971491045b9d0074af91366b05e937849934e7e1c4721d9503af8290f79af3cbb4c4bec36edb8f2c515a7a984811958084dd4d1ae03523d8a83ce5995c1202751e8481274e9dcf2296b20702d93a567307c8a72306d311e3d29f2707342ae4459ca70d98bdaf2e46c59202a19db769d45873450c69cfe113962577f11738736a12b996153bc7e11510e198c11cd6f12bfbdac79139f5f640283aca551f7244d1237d5b7d8c20ac2829803ab4f5c49ea602e4f624fbf3067a2646736087f45c694367951b836dab83a58d02cc4007f13a7d040846a3dd50671741735848d398dd387a60b3d5448c2e50471763ce8c32b7a5504512541c3fde88d7071ece35f3c576894c11f8df8513157d9bf8e91abbb2b0e668c69f98da94200ab15013aadbe65b9fbe5892eb1e6dd04604a0c8d6c00c9062ace6660a2613a6866be17a84f6c2ec6ede2c24ad92a8064d333505a1e98a6b9e4424b310c724db28b9a37449f5a262ee6ad17583073161af565f84af6fd12afd3a2561dffef9f19b6bd4c249a418d70353b9adbb50d3bc117f094ffde7ab3d03808c115ab738758bb8667552c7ef8cb74a74613c462abe8b0c6320be2630051af575bea1e8b9446a91b66a128119a6f91fd6c02329106184d6db6bb276797d3936f702fb3a1e23e1e4806e06d943d117982b00cbf9bdfcd6049fc08fee23e190879b4d0b7d58b956f7c81b5aa99606b346785c76743198f92692f3b8684243beaac937d1443291ce1310ac4e69dd33e591f93979b03c41951f019b83e8ee6a1d4b78b548ad5ce10645add489b44e897043946a134b784bbb6267eab7d7044992f69482f202ec242816ffd50941214daf3d528671cfab1c4628ab2e57fca936f972ec0fc0730edb215e7007f0bc2d8bf635e7cbb4cad6fe87a2b60d7542038605c2234dddb1faacf5400118c470d63c1984a42abfae535e76c581de80a604445b497d116c9afa8c9b0903352223002d313a310a6d98ccc2c49b910f484bd867dae18bc2a8449b67c8885a2fd61da06491fc2103599f016987fd45ea155676ef42e5ded21620161a4a8bcfc9e7a748d6053b837c35314a971ec116b768901440921d204cdb60a7336bab8b9bc415a07c672f4971016c2ea8e3487f0d809cc378542d6c5d2d807a3e4a65341697ba1f695756ffc440bb1e494c8c6c4b74657ecea6c85132ee424f1f2795bf42a87c643969aa16544e69ba18684c53f7606664d72adbc502b0129a9a608fc0b9036f1a86e76786e54bc61ddab0d31f5935bcc8c3f603bd4899d739511d5f54bc42327f98949e4f7d2b3dc972e6112900c31a03c6e164c79aed0cb0df20302b329ad1e161e6c35dd3948f39f5f90ffe7592f7b1bb0dd36552c3664c5ac750f94736a93994eae0f62ffccce742ebd78b4f20234210821a204949a44990746950b10644beabe11b9dd2bfa194a6c2fe9ad666ea38597e8982fb78ca9d8d612932604879bbc419e0ea8a132fe99d2fbb234939f9cd309906d530aa8f4d274728687beadb9fda1231aae6254b5d0be04502895db9fdfe6722bbd7315baafa418119e47f67d721b65e3c95fcf2606e53a16808f5538de06d2b767f5e8d99716acfabcc9478cf586ad1bcbc2b2ac9346d09186f77b51d4505efabddb9aa1b06fd1626b99fd5b9693d9789330d5f22bb81f57aafc67e92cde6303a6fd9bf5e588a412570adbd68ee9772e157b203ed73683dc00c19e2bf13a1b869a3459872f6f88dcd8ae6fb7a22fd515b5f3c0384d1c6e0dc57cb4f29e461352d5767b4420244bd97bc8f8a36e7ade8ba321502704afd8f4d6d940307d55e364989c0fb1a5549454d0eb6339f5e12a9f22550229e53e2b472afabb5c79ada285949181e931eda769158bf8bd59c2f18bf525fd8ee1138fa1957fc0d7ad78aafa643966b3d71a935fad6eda6ac35139cbc430b206569a8071de78f37ad11954da429c585c825c8c1d195e0e6d1b6b509f297e5c9cf3b4d4c76b4d7d1d26e1d0beaeb1afa2129b8e50f60aea025402cfd7cc534391d11f3adaa15a9714b9fa649ee47845e2295e2d6bdd6ffd4de640fb44e6a0ec1e6c397fec9cea4768bc7947cb23361e77600c444b00f28c8a7ea22d0a78d8f404d9ea7d8e3bb35c91826f02da2010d141837bd081c751106b612df62980b5b5dda28867eddae778484276bc513fcee83e28a75d4caf0bd7bfe5db990a2f9cfc1bc8121c9c1376ae7e5791a65fc74c1d5aa4f455caccb38d34c6d0751ad94ba6da3878268883d4ca1d5868e63cf45d7732ef2ce12561de06c86793d5c8a525ddefc8f82d534968c0f14cf577f6b8d7fb988b29de7b6f423b37d151d04b444347c942c6e24b8e4e9cc74c960eadb708a93a77e198aad6348ad414d5a9ab4236ae011d27a922a2bfd6d15d51bbc12e3059f3d20b7f5c5957ade2789368741428036cac0ccd0a477a224daae42ead69c0a59123b20e0170dde2f5eb73b75a81de93426f573efbb1165bf4b16711ce971be55a816437a5dc19be95145568c4d613298cdea0380f6844d1fe7b542993f9fe52446642fb2f0786bc30176e3b24731dae9f27d78995e13e9e17849c8c27e7e9d2a5ff2717b61d7c6b782dfc969d4a61723147d1faf26316bb9e30f2a9204f5660913ee948b688da0a15e71344e9bbe56d8602bd5e77d9701d078d7965c9f4c0c3e172b9005f89f9ec03a8b19d12df6b2f3c6a71dd532774d87656e6ceb420bf0d0db527;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9c18676ecafe49dc8ab7adc46ff8c12a6d609cc9cb5c1af557264b338af23b3b60e14e06ac7efc2e95c18f1031c7360d1d5051046b215a557b19d8b6248b0f9930e8ed65ea7696b19a91f78300f7a044e88788bc94ec63f49906a2f34603d9381f89c7bb2441cf7acb32c820a9eb9b7cbaf5a549990481360883bae6ce2b7b336a3c0ad42902ff4aa0b5edc560071b2a0e69e9ba84a2afda7376861506d94de2a5d8d66469d3378ea6bd7978678256d1a3e5a62904d1b1a9f55c489ceb84f73324c9fac4476c3bc29a7dd5929f8d59b65720da93fd941400e41ddf73dbced26ee51fed68f774466cb38fa360a9478d43b512f96e79449d2897bc041ed08f3d3bdeb42f51c16ee8eff0a6976886fe2f65affd8f9fcf112ed756eb5eefefce5817451e217a2060adce4081ce609e443a817909c74aa46ffc52f7a32fc2dcef5ba19b11d8758d1e58e875ed870fc99ed3ed71c513b1694f8b06012d4052deda8e03bb70e8d190b108d3e67717ee7aefdb54c4b39ac80b86ba343637ee48ab15e1c6c4d65f8b7b8a890bbf9e1995a887aa23f09e5d6534aad99dcb07fa6a4c4de209f89b989cc2e97ac1baf1781e2d913cfc8b49390d71b1f13bce5a042b0ec264ba4411e4f3669f67479333471b2a28832a24b04d4333d43163c1bdc10de84a2e55c8c291fda968351fcb71f9ef9becee5c197761d9531ce32d1d4fe5682a39faecf730efc1cccf9a0471aca0fcacfa8eadb1be2cad837901a5244cd0af0c198ad629db51b7489b93796c465d425a6a9cc22c0541e7d53b9c380409f7f75d2a4b37fd13574273e2f9a9dac1af6d09695a9fc7d8da0f5e7d4b3be59f3e4da15e22920feb124492737638d2c1cd8bf4aeaab1eb97d145716d7f557000eb22d0d5a218f77aee1555942e9ea97ad8c90ff2bab1339c9f050f886686ab5fad968d2750a04eca53d6296926efcd7800ff6b5f6a0e71b9ecbc5373bb04990274ba0e80e64f1c98b0b4c7fa5f6f7a7ae081c96153d9cfa1d0fb3c89394c29a28a8b4aeecda9ff882d7787d23b80dba760a7aa3d0e4ebeb7b8d33c01415f1042d89c213aeff06d3c554140c73ff13249988aff6189194f9b0afd5f2e4d1fc513e0137e399bcca35701e477c6d382ddd9e84ce7a2bacff99f060e3bf3cb68cfd512c32ed9d229ee6ac20fd21690b7b4c537456bc34113a8e19f43594b48ffdfbb3ec190c058f40491410b0241b711848c99fda6e9dd93f485f063d5a5b7a616eb91c5b1072eed542b3a8021d79fb9785199a3c11233f0bee0e1e76480841fab5a52dd9fcfcefd5393fe84b20f2a1db74f5c8ccce58855db6dfed1162846cd590b3c9d6603c72dc4e27070bb4373ad1b9a2794284d2693a166594649773949257732fd077f4e1362a30acc0e73520c84acc11d3ee9fb96db5549dea22843903478d9825aa7485741775eded6ba28d90f2e561f0cfe1a7eab4920ab96a44d913e3f96e01ae95b040539e92f1df8a357674da5ccb361ef65cdb723304aa70406d9702dd5b747ed39feb625883384820678e4da63087f7457ffbf4beed83e321359afc78270c78732c6e9d01b2389bc8f397a7c3a3b56cdad450f2373028337a12287352c478beac9769b22a752bf106c7d3f9b8d37c554a999f65d3c0f34093e0daee64717022dabc3f8c3d0042a97ffc8043608af7f85a41a7ec49121f5b831d23a60841db04f4127a2c5f1ce2fa43695a8042822938957e40e893b57157123f42b00252b5600516ed0ec549d7bf92b089a3701c58decaf14a4820783dcdca6af717cfe0996027f3272747ac224126a9acfa0750d1ef23b5487fb766a48664a15f9548d350eef617f06bd7ffc824e2feda49956ed180c2d2651c8a823cf1a2cfe126aa171f3bf6feff6cbfe947c25247539f9405f1da7947f97b22d6d55755c986e79c3c54c4d3b1e702c4a7faa78631c7c3e90c2a9fa95b6a874a7a93055a9d00b5e79981631dd4d9228605eb82484e514eeec567c56a9ccadd7e4681469e8937336f214b3075daae265d8d012588997759d53c81733b15bc54fcf9614d924e09281c5b6ec2d6922b7904ea55854fe14ee39d0288159721bb3917d55435146780aa705f595b9552fa5fca13a0bbcbe9bb9ac3fd2e6c4164656db19d9b042ef702bd365e49a7af7cc5c4597250d211ea6940f05679d8b4d2991266631a907c039a4c2ffb6b4c7cefa5d56e6c834829833abfc20a17c99cab66f54cc75410b37b7fa9074befc8e8c46e9ba2fa1879e1da1b08a807bcffba8a9621e61cfe79cce298fe5042b0856e82a494a0db968c6f8cd6d4831c049701af28bf94cdc5808b512f6b3055bb6d81edac0c1353550c9721139ffa07b0d1650295b544efcb4bef57c4026038c9efd1ac87cbb15150da892e99fbdbcee99b683bf4a7c55d352f4c05413646d6be070cdc31412a541a25aa05ccf45802561f5e8583b6b135439dac9351a9b6f444bbcfa7651f94dc3beb8502c88f7473d0cd805a25528877155e508034b6a4c5d88fdcb85ce2d0445583502105bba4abe9115d190517d720453242b1abcd2aa44d36f39a359a540a3c940c764e27327b12c225f24e21be8ceb13024eae0eac1e2895fbcd4f110eaf056c88482ef7fc7b4543638e7288e7352034e6e7f1db872dda97bf69166cdb01579372b8988ba37737c17422a89b7f98162c9a8f821fe58eb779bb53232cc73ddb9db45678b6738a357732032325a4ede990048c1340d37a9fdaa49cdc33c362a1de1306ce1372afb19c16efc3380ab56b4c45bddd2fb1e079040b7fb2881442a93a5a91613972fa83f2c529ad711f1395c0ca6b68c36861d9338ca5cb144cf7a65018fcea7fb055c7e7d1722b1a541161a5cbcef1527823467475010c6dd7067b6072df567d04f2a2ed91ad9db99b964f2d55155e7896484a77294b8dbc65f49102cfc423ff39e863abd8bcfd49118a0d8800481ded6a0ba01ab5cfc95fc5a76c9bb57d878b9ea65d61e5090435c4c5075a11da8610282b2f6035317c19ab310a1a2f5e47e6cd73e753a688e08ac895a19b53943a12b57e8b5c7914bfcff828934f1bf596346a314c0ec558b7b7d1e4c9bb8953bcbeefca234028f8aa0771db2050d233231acf39dde352582a5c36974161cb76ac1c648ca9206893e244da3ccbf3cc5177de4a75a1e5bf1e3a26a3d25740b1d33419862b63cf02bfa3aca2ce190c0b4a3b852872650ad3136d48132be391a1a27136799244d45cf452c23351d8b9d932903874d1032f777ed56495ab2c2f860e9a7a6cd3cac80add1f40d3cae140f3af27d4abc8b49a5d1e97e6167d6b20a77229632b733c1c8b6967a4f42c51cdb4c85e2088769e2cf67a0ef1894b29ea6ea7a600876a5e19c593075ce8338ee9af3488eabdcfd2b21d28ab3a811efbbf76db73c1db0ca86bf9d080bec2021cf9207068835dec6b9028a2e7678e834b0b402f14e5bb313719c048511cd568703734066329c92b914f067d4c467538d95b49ee27d8ebe52184bbfdc056579c2db2588a8bb34904f13b6e9b7ddebf2fd52ef9c1a060f31f388d75510ac81dc41216187441a1340532b7cb1fcf10e857469a200757d78de93d1e44a494078a47c2f58ecff8d51d02b152167d8b3d7e8305ae7c06570c2c19034bd660ec990f181c0920e510c457773bfbc7a5dd7341c35c77713d9d2e52f487d79b9da313beb0bb0ea5f22717c95fa2bcb378b779fe8c7a82da914304d08bb987c39db6e6e95d0cba3500fbc121ea71c8db79ff3ca0d116ab911e2cca3229c27967546aeb51af5c421c1603dff777a618d3bbdeb7a73d94368f0d1f1600fee14c62be191c975bb3bdd4b885f0ca82a61b6890e60607b207070f9366bcc2e31b22fa533d13a1e3ea09d5e51c3319c3982fe655c9c11cff260444a6f6cbd80c2954e29ba543925e2278f829945cdf712a387e2b47d2cacf4cf259cf3711c7fcc228f8cf714da799a602aaf6258e34e1e952ebf806dbf6280f574e5c360d8ef647a6f1d0b7c676ed105b20595162a4dda82f8ce9c9c77d3c02590c4ed8782f84c308d9b2ec3215ee0e207ed4ecaa243a9d62fa6cbb0577fb69c9d7d32b568751270152dac549d887ee46ec2a6ead5c023aed2e1859a4b4f43dd9e69d410509ef04c17da0a4d8cc39f718573f0728b7ebabdbeb2470c7d43c2f5766b2a44990172f43dd8bfc8ebe3beb59401d014ca2f19bebe56545766c9fa986e16b2e028afbf57b6a3cc7b337c967bc16a44bb4754ce9805c0bd9c68513659d6f403115b6bb14869b8547d44dd8960c62e6d5c4525ba828ac8d30f25fa0798ad4f7caa4c063de34ac381d205f48268b39e02426286c572a74f0f3adf050ae81904da284530551c257699473e0153abb79a906d8763fffb9e9d2028a91650d151cadf7f5f44ece93b6acdd265864c4b58e9d1f1e758bea0ddaa087e89359515f97f188ba3e5c36ac12b43bd3ab938a3e436f18d75c509eda32be95b985e1f7d4c52bd4141455122f8da83cb5e305cd1fe77208bf76f3e0cabe21f93f815e774285f0c6f33eb4c4eaf29bc1e69200e02b9dba20bf7707ddea56d39ada7df3d6a940e5f127fe5ad1ddc6e8da37b4ae8aed12aea05f7a422fac7e1d51c2b695bfd0e6189d03c46bd4e14e9cb1df92f091c161bf7baf0e01b0599eb160c59787e275166eec6667b7565d5006c626155ded8cc42534e2654ee9619024255147d5fbce75df2b67ffcac448f51fddf43d04187f3f57c7472605ef0336a6538df2ddf7e9f1bb28da543464922fea0171f513279c18ea9d9b49544e2400e1cd96cf68bcf5b1d3b9b99c4480baa6b31770d53e65e8f39a50d0d7a7b4a33e986e19e89ca56a79bc7fe00cf334b3a8a55e70070645e76ae4296d45d4378685933aff011c8dc709d8a2794bb1a952fc5ccf8c2bb4879a0009fe8370237835226a4c51ffb6d205926f4385dc7d7166d296d37deb587e7bc1fda99a642e6a7e6b6b043fbffda280b3a1cdb2ffc6cd87d25b7c890eeee5a894459b05ac20050a88920affbe814548f8fbdcd2be612fd275ce40569478abb84f8185e354c4561ce941773b2b0425ff6e8ede9d4b6bee3116bd487e5327b197169feba59c39c9b4dc705af9deb498e9d78b9b7d804faf8148d1cf5592593e3fdb504814aaadf29fd21a35614f2f38a78588892ad42ee992de38333336e9013c7f3aa4e33cb8eb87e0a61852e9553bef9a381fe955f0ef5ad44b69af0f6b51a2450db098d915ab7fb809309f2091ce0a14ea058de8e4c2c65b39ea8ffd7d4a8e388e9bf05890ea7079e224c02cb8b38987d9edd8466f4007e94eaef006f461cba6d534f272424a350820f3cb8943b583ff5c9050ce8379d843fe89154ba316e21520311c463a0d430858256f07f5d338a40a29247f3bf82c7981ab249f18456c41b541c3d44888dc96996e658fcf732184e0bcbec6217208bbcbbc3f26d2c0088b7e2b4717a381e74a57315ff61e26f530e5b5c116efc8f54dd030c2308e397a404ab566463af1957c61dcc3a2b657a657cfaba840a0f721388eedb06cf44bcad960b30d701e0517ae47ef2a9553eb521eb2c57935c7f551f3ee3f821f03d60a386ce9a005f34339bfe0692e7a7a0c55b3dec6b6897ef7d387f7f370c5d6b12c460a9e57bd951f42b9c9e005050dcb56589548cd3f8face15fb81fabeaff5b4eb62956ae65cacfb988a21097fb34fee5ec4e9f41d87fc82e3953a43b87eb06f306ae546863966635cd61fa577c40f84819a15277353df0bf1a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd2ea44a79e54528f159da925655b0f3c9be2b51d7122486ce836864ac21c85e4f5f6b9f2d3e41f85e9452fa8ce5461b70ce0e79d0f86e95c0d587b24333ab30104e34f5264485a5690f901f359a786c7e4eb6e7792c6fb7ca1f953012a0ddea0a4cbf62a8c680cbcbe4e126012975c4629d745ae29c9e11210158ca46388c1e729026398938cf71964f254f6fbfdb6f800a3d137bd28a8689308ec899fe3781034dd9535e6138058c31c8c483bcfc8d4a49e36d072c379377915f6814b80f59dd00aa6ad5ccac0300ddf15b4453a80970f9753924850049e1b4c70e582a894288408f0d79d7ad43564d1233de9c065cb0d507e6872d8191d4ce87e25bf90e4ad6de3b378f534d97e1fcb4ef5b29f54f8b9eb8e2be440830f46e999e21fca9597550245334053edc706bf0c0fb8398e182321ba1409ccc0cb99be01df2852662dde3417f7cca070180e2cc9ea7232502117aa2b879624e9825d0e8d9304c921f84da9f58c624cc07f84ea647ef735efeb9f4c6ded0e876cbb57426120f6aba2f0be584feb8e36f28416227d4707a9428ea43bcad54294e57d4ecf599317ef96aa86af4110cd6c6dbb9ecb4990dd7328ceaa8713b1e6b906559d228a0aa67ab0de0b8fe5295d455e2b47274bfc96d4b035a88a7953f1dc966d619774b59fb2d09ec5709b7e5e38ed6b7d132ff645fa1ed48a698fb29ef56eddcb71219f442d12fb3a7382014f7d2e4098d53eda49d08e1dbf59c8a90bf61c25b32e6578249ad5eed0b8e40aceb823785babb9e10a5ecfd50fc678e9dba38f9a7c6e6e51305405965ff47c4d11bc7201e54d83d3ec586fe9f5ff730b2382a55b793beececd376c8f40abf3876321c73a56a0e560b2b4862186733cdcbf9fefd2393ae242b57942ab4a4b482ae9478640b5003e88ba7d4ee4eb4c188b2548e3a8d94d4305c6c551c3bf93996e602e1860721bbd8eba67bd0420bc80c1bfe8d3d63a2970deaeb90524fb1d458cab354a750e5f2f1dd1608ded653844baaed39bb06950143d5a3ce32a51ab2e7ab252914c5d6578033d848c36ea23389b8de41db5e94459e61fc05bf5e9eeb6a28f56e80da20b1250fdfa70b431c00ef2f5205aa7a9862b04663e1043338bd64271025cfb4cf2f2144e0169c94c340e338fb72fac77c8fab0c149aed962649439b168fb56e2698f6a30d5f6bedd02a11cd76abb4b345746c9e835177a5b66c3a0c4104791297a807cc1b6d49c0b0c4f47b00c34d892df65c17fc48b0c0f8e7fffc1781efd7a07bd4ea31971fc8ff09893709a3ccf25342e769f338554e807b9b2f23d254c9e243ebebc2716fd06fd1030cf95d2a406897d58643ad222e9a5c0b677e04dc6b032dca29ec1f7c3322353167fe9526daf5a307a6835984bc38ac0ea81d59e236a454b7a858ca16006246e7a31d49c315830cc357a3ccd17de8fa5089f5e2bb795ca1b8a360c2386939dc6fa1b61075770f542fde986a311069b96b57e52f60846b383890fa8f721c4f251d1190a5de03d1408f12611d1abe4fdc01fd64201dce6b6de5b7d2ed2e47a848319934e5f7c961c03e0ba9cba0c1993f999368578d972558bbd7dec9517c138a598b4d34e8c847ae1c73770d1bbb103274cc066826f7536a84746d94c98785007320386ba31dcead8ebd23a3fbadb6e612da1ef17a66728f5e7cc140a122183c223b1dc5730d9bbe38ec34ddeab7b970285e87bd10ed73509402dfe90410eb19ed7882b0187f25d711de95d92429fb97437b95c92f08ce9b8843388c83e4b67a7f29aa35ca87583b479c6a243aef7fbbd0779dec7387b19201a13dc5d34911fc46147c76cd72e7bf898155d93162a88f9f89002f78cba9eee23ecdd97c3d7eb506003a741c021d8cdc05143a4bfd95fb41be5a7d06435484690e025b7025b267976a5b38be73f9ed903d28f9e12875e72a02b767128da6270dd8ec7e2f094660e36b9c34a9ff45dad3f1c157beea06a88b02783e974627ce316269d9ad1286012f6a417172ac66aa28cacfe456a771f059207ff08a214bb957dc4d4ab28c131a7159a8e1657fd031e652e56966a8c9acb08009f71880d33aa1ce3739d9e70f13d265ddfaebe635d415bffaa9a274f47483a7c570bae50d3a9094716f913e20f7fa122a76484be5f946023986d8119ad9e1a59ec0d3047f10d9dd2b7f404ce8d3fc202a437b4e3d9c686465b2dd3e613ee1d8c578c532b2b4393504c21fbbdd200d96f8180a10730c0fad5d06aa60605d30a6e3fb2c92cd89b196d98e0e541a82ee9e8a4b1ecdfaab45b0f89f95113694135b26940cf10190c5bd7b02e6471f8176f99a845e0cf2d531ef9bbecf6e58fe74daf2ad94f5d9831daa259b4911ba277c4ea978773961d9166d7366e05387e2d9b38121ddd15644c7faba2b26f53c686bc04434d941d4833ea96e73005870eb7febf8ac3d59a9bdfac19b78d603387d3ce16e8595656838feaf0a2d776a2e1d725193fcc38f425371091c5724058c07609858d454e359efa0ce462873075b990a93ce93cbd9bbdee89c35c5a1440ec651de34a25500f729252564546b4508c632e8c85bfa9bb9b0cb92989276f383aff099b126cbd07afb4420880f9d348a9e9d947abb6fd48332eea614338d3c2a5a70027da10720a7193aada53a6a3cab12e475b065890b25af540b74c7842b0af53d941624e55b30a6e56768b26084ce6e6ddc48cf810591b8ff9f73df9eb56a5bbe76e30468f0b5e7d6413d0f4604bed0b8ef742f31eacb56a06dcafa8d15fbbc331b97aeaec3b80c041af14b5624593a36052317ddac96b0587ed88bd6f4f64477f743cb2e8da12e0a078208ec88e6e112bd20976bbcece5ab904926a15d25b44d6f4511b1b118497b317cc03c25bdbc5b2e9878776c4bc7acca9fe7ce096a8f4c60fbd462a0ceebc3fb0e45cad047a22ba97ed070db3384d8fc098f1edd8073e46f23beaffe2aa67e80908529383b5a67717c182c95f35828c40309d3b16fdc51c11a7c33727decb331aedd189fb8627abe48b10e0d325a92269fd0b6daefe53332c0584c5a96e1a29afcefd74135e0c9f1ebda871d849463c6b62a24f60640fd3e76d064a4ad60051209a834a038cfb2aecc7bc88b8a4856a4417856c94b8c51863e1f21c9c42c1790ae390e0a3c6be5b845b5a866a7831401dfe09cf4bbdbcfa3f536a7697261f7031028ab7da8e133b9df8db97061051db80ece76b5e045ac81a8b1ba20bfdfdd216a3641624c8279a8a61ea6a597663b7918f7709c4a8068f93fa2524afada24bfa939a851e599622bd742711d0c14bcc029dbffc1c3246967b407a0b2ed39302c52efef2129766bf721ed754ce2e5d3df3f465016a0f2609f5fc74fa3f1814d3489985bd3de8b7ce75fce0358bfee805726d3f3af21bdad2aa1407ca1d3a6d028797453fc8e1a1fc534957c5f95a4c9997ad5fae526eca31090c11b83ca69dd88b583975c750f0c851effce9e3e59396c987de9eb1673308e5f45da23b6bbbba8714d08b632a1633ca3263c9d77e867dfa1ea57dae7af4227fc4b7ea94b24e97ef49baa53ec00956b5897c12f265dabbf71c6bd554f3346ad9ab4de1e0232458683adc2fd2ccd707f30eb677cf1e4451c637109baa8b57baa4810af3c8c9f123981403337a584f3cbad3465b79a6a24fdbb6aef95f95cc603d134747cc6d8560b2d4fa8e92c0247e92b27da70587efef90945ffb24b6984fdb46267f36cebcbb77428d423aa46e59d885517baf25bb6e6a574d25974c5c8e0db7327d7f4576d440ebcda807c22e0590edf571d190820b01f832d567653837799c527a8763af1e61f3f59c3a8b994a1e848542ce940c7235bf945803603e17e1620c99ec0d67966da8b8254aca1a8b0cded40b0816c40ab0539b5f74f5afef785e138fefec8f6b1a4cb4da13c4fbd1f630b3c398855c5fb2dc35ff994820f122df3176812952b0f14269cb7a4e0a1645232a114c1cb24972f768cc498a9cd5a11297aa24d66c4ff47c436b5ea08fa72111555e5cc25a4ea1e0600871a8c33e74241e647a07df8d02c1aadf464bbb5e2e4269c3c0c732f5bf113d62b7d9c1e1cc70cb576bc58f48916f7744a59746035185a264e6a0cef356a01ec464cc324e17c0466e553732c8db43c541a53225c63e47446c58739346afcc7b60b9a93531c4e1dde05813c7eb7dcc2a34ebb353f9fb684f60bbeef06d13dc87623f1116d14847a6bf13a86e8aa2467cc6ab9e910513b0896cf859b8fb07f65abad0ad53a3891b2a08e63fd8aacaf37cdd9589217c1a6621f5ac0d104ce230f5519f99becc7a727ed7deda468293194ba35d9ec98f310fa0c25c2b9dff1547eb23ecaf878b45840185b4379372650397247aea9c09db2c0d936318c1b1158335bcf2c3af2b1eac49b79d87335ae9299f68d5f5259dc30b4b7b6293afb223b6ad56f800a7c69682e212bac5b475fb4a3905708e812ecf2fed4ac6d7dcf074918b5c7bdb03ab177bb9fa9b777a97e807f391870745a48ffac57323131fdf1d32e9506a78f95b17f99a146fc47b934dedab5835ed2968c88efb83a7960f739448ec173af52df8b9285dbc9afb89df6b30e1f1797ef8a41f6d095285617c0e76a2e5bd77d11d31557488250dba683bda90116b32db5b5a7e0becdaa9a1a599d913c6d204882ec95c54f07e3ff7a2ec7c895a6bc5abe13fe66ff7a3e8ebd92a6cd180a2727af68671f8573b334a280e960b6b12411ff68d9ba21264314eb1e608562e5eb4331fb5c87bc5ef5c38b538207e7ea1b9a898e143c4c6f935872c8831a2f56e3e9f23fdc791750340643105488096ced56f24d3bf32c3d1bb7e8cf79d30e826559df1103689d3f90079258aa991c65d4efaec830aeffa6ee3f07bf75439a35c7a0ba769fe60ede34f8e3442c5820041800260dab4bfb371c228c5363ec67e823850655484760d09ac2b7fd6c2be96b113c96aae741aa171a1015a3f9ff1687cf006f7f531c6457ed61e3d22b61336459f349eca47e3ccc55f996a21ce40e617df01468cbc9b73f1b9930380c102679bdf857f26eb943bc7755142510d506125d5ce3c4d2e5099a97ce6a6686bfc98f5c7a40399dbabf7258d69c9b4b8cc096f2e8af149ab6778d719dda97fa3dbe3422ae2d68c470ed84e38e683ffdabd345915f94717dec90e7d06e42453eb25afb38aaad79ebf0a03fb3b2f7072ada2efdefb6b9c602c9f94076c4c546183cdd15d5c091077b070eb28c90e7bb7c2830ea0ddf801718963c15a256dfbb46116d6d3cc9f10f0de7506fbe200184e8a6e4dc30e96afb45baa58649c6d685825ab70243fe193735634de96ff960aabcb34ae59a84d4ccdb282fede4d63084fb16f32affa4ae3679369738848f29e0669805476d2f2fb28ff616115a9b7ad0f64fc9bd47c8bea8099b5793fbed695c254258f18b84ad0a62460d483f3a640a7dc44dfcd928cf1dbd642429b3cfb787426bdee1f5ed4403b2d3660f9c7b1c1fd9c4c63013f7473ac38ff29996d72fcf0115d3648dd9010414f841cc7c7e23baa423f54933fefbee78638230c5ac03867f36e6d1b623c57d256ee5144b81d019521efb9df91537c8cd46fa5306e96d79962c217a1a705b1a9ef25b0c4035e6d38e53a835b2990e7a9496a23ad73e0e05e2b1cb53764c2ec7002fa726dc52bd5889c86b0db1591efa6d5b0b0584f898c41550b9bd55dfa196f999d8a31f42739dc4eed64648983d14eddd8ee7a93e4ce7b6e1bc540421f83f7c36080ac8d8ee8119d5127a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h910600637340cc3e28d02258c06c55f91b1c2d0c1de015d16b1b1f92f3bb119667446e06ce9a8d48b313c888b87343a34c590d76a2e5c699e093e263a80aef9e580f57c40aafcb1f539879117c30fea5497bfe44ed5469ae7e82594a925e7be18adcb5873fabab045db07b645375d406cc7c74cd8609339972cfc5710ef1663cdd8e73922f64f9ee7bf3fdb828b5ab70beb35c7d7054c29fd85756ab1626fc94ba94fedc51708f29737268daac6fc80308af51e9429bfb7c99bd5e51beec443c143e175cdc06f27b88219e988e6730750055e35dac9e830fdd356d2b8acb002c2afc0eb8738c84f57d51294e64d7c5311a6fc9bf99ced53982e2d37ac07e342ca432f06f49325efb1eba96010556cf855b67cdddc81ea6f23b77f396aecd717cdc3389b544c944cf76102217e1d6d3d8ff220757bd074fa3a48c4e882daaafc2605acc16d8eba25dfc356ce7492035d69fe6b1a437967e395da2245dad90ce9ce8b880d797b9143cd61db8d7978b6e961e927b199f986c79b81728a6315b996476bf4be7272097b12947e25e5039849dddb673b5648ae20d69c0323f50497a5e6f4ed8df100d344e7cfc13cefa617d24bf71add257721746bbb4a94b8f9c9047366234c099260451b26f6c4e767ea50cb652f8eea70c3bad007a51edac9d4a47c34b20e00e7cb1508f30f94ff78c3f36d67c95e31d173fb542a0fba213a21604e1a6ea90197783496e0ae61221e3201601a1f24341d01b83276aa7ad0db033398143d69d0767ffcd06a27a636546d395aa0fc7bd4d3fda6fb70e9606e445a5fdf0e716a496c9e2a77b555365323d53ccc2531ba2fa78bad34287283bd6549f41ed4a4278c4e5dd9b860d20470ce88292cda3c6b4a2a8354e699da5fa319419cf60adc73871df5ee0ee714dbb37d6a6aa265358ce99b1948be8ea7a7dced89c24c3f7bc8d531df9572ef03b63fe515e9d7dd731a3cb5bbcac2ba98f19357db653bcb36711862ee68c399284dd2d9f3c33e7eac79fbcc2de4ec9a64763d013d41b536f4f5d6fb44e5087dcc9f4d9fbd5e1125f014b473f10417ef4ce103cf16888bcf45b429a956d4b644cd82ac8283111d11d1685c13bda26df140cf3aeee3bf9c4be2c09ef9b7b17f9c0f7001c621353c0354e83dba23361530b62e8e69d7facf4427a9eb6d96aa06b9cd64f3ccc9bd945ff20c9459a33595e005f177a5bd265e0db0b1df165058796fce47bd0d5e57c41df4fbfad0bbaceb767fd331be5614d15f540961c33cd66f1b69214c56f259e4afacad1ad7d4dce888727b921cb82b78e529e645d796b772c2ae66e43a24a334011ee2570198290f78b482f5a22e47f8e7896ad166137df3f0f12b4f3c60d39865596fe910be78c38956adb6bf4d70c94d10b78e6cea61fc7fce593d85f4c11b34a6ec2fd48c6c72cdafa5a1207c2b3eec585c648048b138bb5ebe733525a788dd8908772808d3d23a5c2f9e2ec643d30082086ddc87f7d03fc384c70c26cf00ac1f0d07c59cd753be716d746036f0dd9f0aac581fee9a329a5e11d4aafc091731f18612bb6fa2071dbf0aa1ee2509caeba201ecf1a04df18c0b6997bdd7ceaec8031f2bfa54338d4c0e19351c2ed3e669ff7c38f122717d16ae14dacd5dfe103e5667b012f36b92956004112cc03e3ae99616a5065f322df3da23b5162045cd945d9c77ef3c9c7c4e74495d419c2497104fa1a39af3a2d7e413d3dac8f86c4eb7cca8403b9422c956ac3de508292607f3daab204bcbc10b57f3bea13047e84dfd7704ce4d51c2286d0307c67cb4b3240212599209613643c0f3637b4bc3797e8b8afd5d5b9813f566b8c7a55532e557c908e7d8920c921beab71f96dbd24c5a9c852d8c21082d65639de1de85ec0e081268c18bb8e09b75ae26d1643092a31426aa33e76db71235f45df3deb114cf218444dcc70a8643a671175c928f725a6fc3cf54709afaf28de490e41818f07f4f022f006a80ec51882aab20234014f4260e33e420df9023c503e4f336ee887192684dfccf26b766207f095b7aa0ea1aed1e2a9331a460275581022065c68f59de9b0d2da1164e70ea7b04a71088599f9c68a8cbdb34999cc1556894109974ef50bc42041f8b7bc86791eb9a0b0f186ad0d47dc686654436a8eb9d34142ea06124cea95cebf49f844368c7f4f60996a27d4ece1e357fa013d3c53a0277acf9826bbf797c2c2166c659315314c380fec2743a15013ac434e2cea7a33f10b36cce0d19336412436aeb24f1e0867d70cfc4e3ef4ee775c2d9f0bee583760b0c28d8116239db20cec898415205e0d34365927a0574c5d3ad93c2ae37bf375dbd5ca19fc79ac943e4a84bd33efaa7de2dede6aea13929e41ac9133a647ba066f0e4efb562354f7ce41597fec99a544f869b7c1573a398f5ae02028e5833bded6c536ba7f6c751280b57f76eb9b775af81ec8879ef91b577ff94de2284354a5f7a377e4b99c055c9f65731775cf7449b0bb85760d35f4a43a5f7199ef3abae5f7a4ddeb8bc731e1a68062d7a79fd7c1a76326d645e179b5b830ceff46c20a1efd5b3b8b05bef142b4e8543e3097ef8d43aa47df6ecb25b63c75f88bec6ce1ba9134e2009f763a1b2163649b3e7652ecec4affc4ac48041bfd19a6230739bc3bc5714d5fb1116e65b8e241f1251739996362442a3aeab0bca5b037682c2d75446c21c676ace3dfce2ba260ef8e676c9abc1df38e4da2e63ab44a367dbd86d8cee4bf73dad8aca7d10fb2aff571075e3e23d11fbcdad5d57214481e1a492f81b93131e78a61a0137f7b6afd615e4dde4d458db383afdd060878d1c4c211fe88b1dbf1f8e689f176ff701b6c45206672fa4761b5408ef33680bf77bf972d9b2a2b3e7155703094d6c2d91d96f6625839265c52301f8080be922004e60b9b2f62a16281859697f18f85ae8c4c2a1b114169e854d7c137a1b56de71b252c35dd9646e8d07698cc9e5c92514b4025648970ff35f8dd5142597d78084905ebe4c1b4ec5927dfd37315a2e0aa3f5d6929dce23e41c032880b2fc5f510e6b261cd27a9c8c1b991700c614fd628d4e690be333edd077b77778c0b5c4770fb74ea07c3134eb39d70823376c8e7257e299d3d044f0ccf7e30d298ac3109789e20fa8ea55dc901a7dcb30dda02c48045b1f89ddd60b083b6e76a66792a77d27dbfc406ee10360d8ae1c1216b16094b55cc37dafe8ab20701bb8c0e8a7c139eb7a17f8ac3c5f4f8f8e1de7392a48402c3c6271264b2f1a592de7038f17d90a7c78d8d6fba8329b5de1283daf57e5a2790c9af53172d523884bfd8b6c9c0971a9645b0f9d1cb30b5a01540829f071d2cd23b2263b9d39b09ff5ba8efe7976acbc3c24f0f2a70354c26c54f2aefd9f8bd07563d167771acc2a208d6cd02e2571ae25de02e2dd57a27f9e70ba747e0847b687ed684bef10bf6801b5d2887c6ac4f4739cbdaea3624306dfa01a2fdf213087c991ba4a05052e172ffa51eddd7366b76fc033d931b72126006d75da407ea2a758d7493b89e9bdb761d5369cd9dc118380df4146f9d2349a440f09d98edf8513a3b7b884503678ae68b0589b807484b85c2e13c22b6cd2d7c60c0844e87ad4a9ff754e78de0cc43a038bf6b4bb3afa3cbd8ff86ec4e9c23c6838e7be929877b292c71e3bc68005d409783d956659e9ed67615c3b3e3798993bccd8a6a6397091abe755a3b6a86d808bbac1fd7e9e92a3909ff684c50dd32417463fa251e31d514fb1d3033c8e15445e79cc6975f704af593f88cf632c85e181dc63d2f5472ac4109b94deabe888ae041f262d2a416ce4371fc5e32e370009fb5006849ff1b3436f31ae8ac086521d76d3368a80a7643556ff79429a7c31bdf0d8ad40ed0e850c3830bb0b20636a613c1ad9c30416deac31d43062b247d37bc0a864000ecc576bb267e9540fbc0993369ec1b8f32918b8aecb9ece4d5a1a9efd9276206e878634412009bcbbec6c2f3ea141064cbc93b807be7cc331c961bc25c9b6f661c8e08c4f22d7d5d71bd155aa02d83bfb5e0ed14e281b1df76fa61a5121b7085eab7ca51b33bc1d1b20082c5e51097f1e0824824d55626dd911b5b762e827948ec1d646f475d3f6fb4853f05e4a125531fc249e0c28f23e39265c0581c404a72eaf72bab7179a288335cb11c414dc312b023e4f16ae95f7787954d272689f332ce43d21a1b8761b86c62ad7d4f08a4413a6d93c8bd518ae601229dd13d027ea050e6b326647edd6fe06d310d3a4015144762a8a9e8b53d0c3e6c0fae18aa6bb407d2e2326d53a38b17ef471637368d2cf2e633862f4474b871dfaac2ea29b45fb0106b47410c94e23304f0fe51f2c5d1050f8091e546b3e5e68ca1f9b48900ea7c0c96cb4b56d4f777a0b744f8ab4032553f4ee12b3cafb1c473015f48733afde9213a762b553ae50d72aee3cfa78e80ec106cc9626fe9d2b651f184b04860c3a9e63507a615a6d3f86bef8ae286f8fc9e1398b549271f4c8d191298d4d5f15c38cdecf2074e5f1ba110fab332175045e58a9cc68a48beae600ca1ba9fb72cd17a4cca62ffb5d997351e0782a012603a5f15722e2b0eb12f9cae67079e8527ca5d0901e702290374ca57a64c3c676983dfcf3726f77b2d4c5400c6c0025934666479b08250f3e2b1075519f39fe4e10fc5d0ef6bfb2b1b8e228dad6020d647be9d907168f2a0c1917f5b15c648847aab6fb171e59ed8917645dcdfe4930c3dc0438c076db64fcb7b930932ddb923a3d5b5cd90e46910a7a788cd6decef30121762cb52a160afefd0ce2291e24c0f2238fe6423010a6ae004035a1d5193de87f80ca4f04b9864f22425ef91263c91537821ec12de3cab83dffdfbdcd4b5ffe0ef2b358b6b387f2027a9732615f7d469bb7231ca9bf4db4298206ebf5870aad7c1bf36c622ae4b027cc10da2cd7ceec727ab9dfb3fe3987ea6dfd86e8e24de0138984fa8d80c6ed2bc963bebafc8e333caef3cb5310b4d32e92bda508eabbbedb0c7efaac656c75d0e8034a8b2bb600654a06e980ca3bb473bac6863e5de5896e14efedd2db55cc9a67f00b9c1030840e512a59c1b05387c09641e7e380acde832df4661cc3a34aadcfc96b55bd4b88ef21ec30fdcf9d3989c0e4917057c9e4352a68490d7a89d1c6cbff51a0e227936373f9b8b0ce07816919e4da0b37e1c962543e6d9433e6c08bfa5454df20c9a3c12d50a8ea63b1f1467aa3d379c110f85e03a28ec83421a55d58d10f1e16de9f808c75e42f9507a1aa330a9c0d87d2f60866d23409f387c557714541bcc8b2f5333fdec8ee130623187f950ae5ff6f4dcf99c2545f8523f441b6098d6f25f9319976e21de1967c2e98284f8717a0b6478544e9040f33833273e40daf51c66b465e59e381da6c91cd6c41c434a42173c048172c8acdfbb5c290745aeec121a8bd6e571a7b32a0ad601512f22a33bda6d5ed039f67804f32de7b7f3d2f590beb5225be2420531bfc43dbe3482b65e41a399792c309dbe9a46a810fd1df0748580863ff0571ecfc25dfedb45de5e7448342b5a7ffe0fc7f74d745608c72994c0b03b9c12dae9d022dd9bc08795bdc8cf229aa51ab368027dd647bd6220f5a432db5553637c69db9827a98719b1e135a4439c7638657c13dd7a032beb190100ab59faded0f0d1d615a04016760e9e69ee09dc529a2287c4621d4eff8e132bc7eee702c5776f9e4f9f6fa6c2de7d659b45787ca485f882c2768c1e4fd9f768922f4c5593a609e2fec4a08f6493e89fc33cb5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h82e09e4e112bd5e5fe7f9ad2d1f0ad660fa27feb85b922fb65afb4667b7b7d72fedf14c040159f9ac59f0edc52437407061b6b22c0e0663089aa2bae2d6ca42aa93e0fec41fff0e4e7fe688babdec369910b9ea4e4b816b39335232bb0a7174a0321f2ad39b8aa37ae0e6e8acf32245642488107194870d7e4c1aea4ef0a1cb93d9df150fb36b9a4396b52711f173fa025073da6cf13b23785ad38f3dac8052e077641fb1f3215ba2f924c2cd36176e1a70a5712877758ad7b9dc797cf429741b68773557a29a7ddbf093c3a17179246d3223522695a79d0036dd11fe4d3e9357227a833a9d664051ca6f2b0ac6fb274d2c224c7ab59405cb63af2931d490b5d7508c37eecb836d5b86cb6f001fae6260bb31fc91c44e33d52ffbcb6b811dffdc5f8f44517dd8f9ee834f881f011fd20c4d48c07ae97f38664760bb3e5f059dd6411ccc7b64bebe25d7a2015233ac7559c76242f971be5325d3e64822a98e9ccad005f95481e5ea293c2cb9af9429e89d7e9ad4b66af6d7c9f6cbbd00baa511c1dbd47be8db36ce231b72a264cad7dcf5df610a3ef5bac944b3e0ca71cfe0771dd2779b2295bf7ce34c397611bf738d4c794bafdbafa235b4a2e567b3437a6f8c6112350db455e0319e9a82414c1966fc9437284fc99caaa2fb9c1983b489db00c99068965c81251b939eaf34cfb5af5d30100c793724d69999481b7262e4f3f07d357324226bd7ca3170ba95104b804ee7155c8e5c0ded7c562ebe3d76be83d74deb1f7ba8e090124e7ca1027644312d8debd75c69a8e20d729c29ddf45bec8d1765da3a857438eea12233eefc0009edbbe66c0ee346d61edc02cfd7bbf9bef806d47dd01841727c98ad39674dae9378b35fbcfc82a6bf565a443d2ba6800ab6600a4265e3676abb54bbc95c514e336324f55201778ac3cdf54aeff23fd3d1e9544c61929490ab5b8ccf244ed1035919705a810c11ce9b16133797c61f7ebfb5a86655e844caf48c1d79a868e27e41adb2b4fbe3d82f2b8fa8624aeeb5cfcd8e0290826c540e608f82caba6a1c7b2c6319577da6d00b92b3717eeb1ccb910958a2dadff6757ab6c69e488892dbf12985d67d44a26438245a385faed31d26abb9bebc90b78fb9eee078e8f9d9d1714b00ff32a3661d3822386f8eed1f8831c32e23b2dafd7876120c2fda326207d68c41bea80489ce14f9f528996aabc331fc89469af21152a4bb98e379b33bd0403c10d8806c889337fe735bf22103aba2bbad8c7e4298e289566e3c6a9a005809facf1a8f0f5a3da7a1cc49db78935c8ab953d0e6adcf40ad3e17b831fa7771fa1f1dc12526de2971c61d7b4056de81d77d9574c8b7b3d7b4844fbda78f36ed535304c55f412aa540de488fe50d08bf8763d2ddf2f46825a7b53f69508dc1f17f8e6a942351b09edea46406af67447facc1199ec82fc57cb02870d06b9eb0b66ad8ba40f7168c004890255aeb932c56edda1482bdef26e77ee8653f85c4aea31e69b24b43fc428dc6991c2f256f0c77e56f7b8159c5d86daa63cbc294bdb9b128fb7395e106b4384222c2125188662962dea8ed2105beb172988283937c72bbd4dcede3471cc3e9e50c36a06f240e83b2a2b1aaae9f7862abbad40229ebd32f54986ab077247eac166a2a4cb09090736fef32a7b94f651f002055af205762214be70b043658a7cc612522ba90e8efe20b1c2fb716460a7dd4d9c3819c93bcc4376604a82769c2a0948361f74dde73198f5d00066418853dfd31e8d7f37811b5edc24692b34297484fc0d2386b99bf299cef5eb6e331ae29ba476d1b173c33de661a3b2c5a67f19ee3a7862fc6254a7876be495fb8c31e72059969b87fd9014ff7210942e39ed68d2412dd159e83503b2c8d12bde27416dc01f4d35ce6b62b81fe5131a71a80dc7112fb64a1bba144e45fe799c7d0b5728c393d0e0aae11c817d3a8ead0c138b07701254aeb0749141c4ad19bd9bd5d1dfd9ea422a83a012d479bc385c316ec40b095a4d1d7585c6a24206be907695908e88b3587cfa341e01b8cc0260a3242322631cd5f3a8cb97d29d2d6b553e2e832809b57c9ca92d6a0644b1d15e49e7c26669281f010f36b40010ca999b2345fb05dfeb70553ae17417ee4b70d13d20ac7bbeb25156fac892abd913a26055f537ec687b23a672118788f26e55258a8a7aefcfac2a8fd20833bfe987af210d1ac8fdf5bad0a113223436d1ef966d544fd0ff474144e47d75eb744f2e56bea5425c91b14a5569ec65918a849004bf836b2379ffadb91a3df7980de947bcdfde0a956b0225e9566866027cef1aba3d3503733ef2e1662b791dc602ddc66f8515620ed31fabf62b9e80966399304e6c2a66a22746df9398ad9dbb140299a80919784450f8a2b1141b70faceda42c92b4afcc3dbebd6b47698817a95ebbd4bb542e6d38b73d4d0d748074915c867a9b95c309677c64ea42a1689fb3e41ae8f2e552ca222ad2209dab2600fb35fbf7b78236481058f23f41331b42327d9d9b7736b58f36c231bf0fb8a08c15f1e5ea992a48e2fc5786f6348f6c02e2a99dc386d1c144518d0a058a60e16f27fa5d7922dc419224f19f90f8fc90a17087c913be8143838428109bb2e39795d85f0f83a045c7ffc4f7fc62ede414860bfd05ec9b72381f9601c875f0ea6f25f08baba63fa20bad70126f48f79d349fe3a886748dbb3f2b6dbc0dcc365bf5c9eb4dcf4482707b64b410025a2df20cdaa55473d5527f02d11c5fd281b49fe0c99d7beee79217fdb7169cabef1fb969e2bdd68832abf66b444969fd58eab605ce1f9b747d5bd36353b387bcd4e0cda82d05f789e3a72548918e0483bea5832fa4b85ae21797764f4f77cc5277b7543f8d84b2eb18c12211755086f8125273a4d039f7333bd4e4a626f7ebe18e40656a0a649bdb5c375caf0a20eb926b56be6a20722dd4e5396e7feebb40306f5085b92ab427e12afc62474910c01ad82f4aafa6039f5cfc7ff6b832d22d88c9821ebf65aac496bdd3fdf99cba16762e5911ba2f87fdf29f0d9788ad43ffa9ff4f7a7b8e45cbd819c7c723de167b3308512890e70773d2b113efb6c3b579804b493fa86e954ff990ca9fdc73c9d2b3de05024e8465123a99ac994a27eac935a1d4e0654ed2b1ffe9d323f4207cddd5476a9739eedbf7e2de1bc6151d92d5228d6fe944432c5d22f3e20947b3b4428d119359270e782a145ddee91565c98962f490d778233098814b98a6b4a6d9b3ca6e4b6f46320617a13d6ee92848409dd47378c029657832e5ce7ddfc3cdd87bb03dc50acf4127c458c56bedee89fd409ef45bdc128f3de67e284de94c404ef9794d1104efaf298544e2635ba448ae1eaec95507c7aeee8f4c3a4c0828fcc556278724806ed748f8cc975bfee338b7b18ddbd8f6e8e2ce4e27e27b1da8b550ace9c752fe21ecb2644996e7ca959420d2acddb2b04ba0a8b8e92705a88595ee7f4105373dc2f8d5eeb8badc851dbe2299d1ce8b174b05572e92cdc1e210de9e4980f4e3a4f30cb243a54d52a58b7a55dddc18784100cd899b0b1ca6c994ffd1d05f0975997d7790f52041337c24d8ed26231252508a3befeba01fd329ed38df9129a57f6524a4d3fb8029e6262afd654f18d781e1232896e60411777c402f15c920466301fdfecea74ab560f7f16edf9c56695c7ea6b6dee95f9630c79fd19c3be9aa9391cde3406e598b07e7e0596c07a610c983c496bc4abf156f8c1671794c8bcce21394198223d324d49ef643a052a84bd22d14027e7deafd544c83ff121303a277f60d941c28cb9e17c74dfd70e457fb0706df6a002c94eb13dd4de2aa0a3f4ec3d31cc0ca8fb3a9dd159dec0847e225a6c4e1f47baf1d0ad0214da691782452660730df8930470eb3c333b85910b91883aee7ad5cd1f9cd624d53ed62e49bc4f2776cb49fbc6200d81467577eea4af01545b0228353aad17b6a5100ae74ee23c454d23333856bb1dc6e8ea5fc5978005dc111146e9d4463156a89023ebc7667e0a5fb0eaca49cf4510c1a602e52520f9e44d7082fa895391c5984ade0d8b06d6cfa093fa415e32d9bb79abf0d71871b023d0068bc045a2889df7ecb7a254db20d519f9db901bfb6e0333e15ce02c08b8ed2939a272e79617bd19dae471a1650a8f7c5c4d136ea6a56c71d1b7dc4e791bfe807b0aef9d8c2c212b4790a2f9bec3d54dd98710a1fef43bd620edd48190dcfc56671473bd8b399a32cfdd70900be2c12675f9fd7bfe87a37e55a910df50b461e1f5fe77584dad01f05f2613183322343ece729207899c244901930b69f29c8f91b54d2ab070e97481df99f1d21c12971baeed25cff53d7dd215e26fc1d1cec326eaba4f48494902d567f91d1464e3342a375f62a6b935e70231599751d8c23b520a82e314e268da504aee92330997cd6a382267d86b02af877d2ecaf93294872b7fde0b7b912c456c20baf8b5d3fb4ccc464d8b558ff44e757386e04c2617da287f73263f6a15ba196bad2541f21cfdb6526f336307b3a266e0d01b1dddb8c7e54ad5831b9abf5df3789f20998ecff39347a67dcbf48110082e5e6c1deb9b62b1b201cfe72c512ffc45d3e4efc05561750daf81595e028a4be000933ee5d4bac801f7759ad9455c92038946e835ce03777e9b35a927a717ec7655a83e30d31816ef10e20cef7a658b344f78f7dfb56374378c94837b5cb3d99afd93e415bf3c26abdd30ed6f1b0e4fa25fdb2ad3b3f372552d34044ed0c848302f8880040f2b48d4aecfa004360d359b868c5795ccaa5c9208691d1f76e966219adb1cff59837872c2bc8fe5d445496112d489531fc86741a6ea995628ebe9cf02bb99d4e8ed464d42a4dd86f3e9efb18eb7a7321c4b04002c9550001345d77ed04250c2d8e9a3f92d17ed4503e1466e5f2bb9c8b0b35664b95c42237182d198739626d4060cc92b073af53c7bf60f2d5ffd07e1c5f5a4670bb8c49fc44c4300c8c1bfdb3fe95ab7509d092982407b64655f4337af40fa08a56f72c6e62c657a4a12cb39490130726190ed5be0e938b9bede22f880e31271f9c7c3464853e4d26dd086537dbc73ec24db52692054faf0cd1e794489366d91f41204f7a3f7dadc8e7307c20b809058d22ea274e7da46b13cffaca5298d452b5d086fa579f6a0af1bb6c3cfe105577fe7d9b0f655e7777abdf3c6348f72da1822069436ea8192b9aaf18ef895be2cc4ab0001fe1fa4db792fd3fcd3e77c64009a5b0b5600b869871902d5589aa93c65756f8e15fe042257cae1b610f1bb61d81815efe4d5a553c7d859190f4878da5613489505275db488ffb8cf4af269f603fb009d75dcf9522deb0cee0ba5ac4a17913a0bc694611b49fcb252413ae7b659633ef31fe55816ed2a0b25d408fb3bfee60a885da03ae04b57acb6f00864a1c914f0ce4d923e26fd5eadab727ad7cb3d279ca97c637b9a1fe704404898c2b637c0c248fcbe5f216808a4180f3e8dfd4dbe83edfa8a6d5d4e75076e1f0251e665b55e9d7c66a2bf9fd3a67d00cf23eb7df966d6a519755453cd93c62632156b03a370889e05107c9ae52b777a5f42c03efdec4eddcc40a8ed02065ca5fd0393cd831082ee891ef87b7d0e6dd507d8bd0cdef385be91fa0aaa7e1805688fca2d8c748212376d3b4d49fbb9cbc1a1cb198a0933e1a75ce0bd95bbc2751d94664648cc9a8f41a0bee2b7e9436e7c0cf943281c9009a133e74eb96fc08c48ff935709a5d1e8a4969f67fe3ac57a654311474e73b458254;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8899f5bc3a7a74ff7e2f1262f22fcf26755e03998b6ad8bc4fde34651846ee6b2a433b18aa2486e81a05b0e63b7c4e3443b9adeba3003d8f2d5765a17a76cbe5e6ad355b4e4d9abbfb65cb0b93b100aaddf8854b4d7d0f8d88e403152464d0a18b8e5c940cfc52b3ee6fc995da838dfe2552123deb1ff127ec64e9e25145b42536894e3f11e2d6021a0edf0312fa04e5a74125ef42ea4b85723eb8fc173c2dabcba68ab4edd15346095e0a0692b6674fefcfc9712c955241c8dec74fb040d6e8f230a425135f20bae0119a1e4afe91b95014837b58e6a8cdfaca45d239452b101a0b778aa60d450d8d3dd1f320d305066b24fdbcbe194bf1fade9702f43c2717f5637a73a7e30ca2a8437855027a8176f5c0d14e752ced6c65e8a8c362151185e62353637215292c2bab0b570901d7ab5effa7093b9bb6021b049fae1d8b58a57cebe7deed9a074a830033e55c43f5f1fe1b0265d77ccbc9d41d7e88edccbf477dfe633bc2fc369595079a3f2c6f12e096a2284737525c770873b0d114e2124c4f1558d0923bebf9a2245319f23a39937fcee635fe0f96d8fd07da62f316bdf6eea89f1862a7240b637f60f7c627766be1cadf50268f54333363e875e01e752764a543c61a98c67d03013427a90d38b3447ac919f9aae41e4a08634a8053fd0204ac0ab3783299eeceebb3a8e3026c42dd023bfa0dae7d21a00b8ef0c17a591601258f23bb8bce7c48a2a114720a91710b8de46ff18c60e8d65bb5a0d0969a717499801b6e766574677d2835b627f07f9e6c4a9d62747d2f7ae729cc366366e2a00384f1bf862ccb0cb4044f31aa0a083d3dec11c734a1f839a998c11979cc6054bee6691194e557050c14b0ddc1bc253f74917a95e1b63ee5ea8e28e312833fd40a67ea2abc6beefd0d21300807a73ccf6ac3db81b7f621d6aadd162e891f7f283e7327694916826457dd347d228ea3772556c47fe03890ee0c5c5ed3b6698913910ad59bf8e0617ed05ad7fb38146d1cb7a1d3a2350750e18f6087a89b74b177f63aacdb0e5a4b0f8a205ba6089546eb981f5e94d30886c2b7c50b67cd6e80e0e7726c5274ed2159d491cc98e3cdbfe0d13941e245f831233539c5dfbd3405974e10eb3487493f13c0c5af1cb5e8d42b4b79f5c190845924ca46ca80cfe51dac1a05894e311772fce1e0f111c4034fd6e52c2c9bb419b227e1f043b467dc0dd571706f7afa80a6eb58ff35a81d0538ae6117e904ec44e875f75fd6f475651f539c5851e8db219a4b76b4fff4b29f5f85b7f803e4bb9288f2ab3a2ea09054b7621fe58b7a3c6be2ba40cc80e9d9708350a2a633a8288c77326557084c8fdec575523f532176f899685086233575bf36c2bb9845bcf453b783c1d4e6d0e7a56bcb1b264cc454a6ac25de9b77b40a6038c078eea1b5a71cc64926e227cb3a4afa9807d6d07db5c0c74a36121ffc01c4bceacab457fe72988bdae3b5afc359ae21b4f12576b53560f8bbd1535ecd3f13845a762210ea6e7b6fcf5e9e9aa657f90db2dc433f19dbda0b653c1b234628f030467ac110f94426f1cdd49bba8b29a2f915667532f1fd25a27649a5dd6b4c90ba5e1a79266c83f4567cc05c9680ffae3c80de471940075c0c9c8534da4f98177da748f006d1563b7d9458456062ebf7ef4727639dd0d16ab1d93e6ffdad25bbc5be3c9cf69cdbb80ecc063c7daa0e85534b0ed10163420859ba815f629ec4096643f307c6cd16cdb5af6bb9951d0b3985f4cfe919ec85f91e527773e13aeaf4f6683928d3bbb8ee96029a85ab7c2f3962565f6fa6cc8cf0585dedab97edb3c3577fdef1f7b1b29f46484ca157c347e45926367b5ee8eac3acc749829e15423e26bac68d301fa08fc8b1d11af822449fb23ee0a9ece5186eed15eed3c3d197a45c8a654d293b88a5be6cf3b1145ca128b7d43a8d66b62f0aa298be2b41e398d348d8a4936641e8f14daad5e8afbc1fbf5ba9760a44e2f416961d75725cdf505f78b83e7d2a42e3345f0102ecca12b045c2015a00f1ce1dfa4d7972780a2fe47cdc645f9e0bb182fd005ddd237a36e5877b9a3817e5e92d77465b37823c3d44b5ca38f73468100ab1256eb9ee954674b7623d97a9250faa934c60c06bdb90f1030d2dc393d6f57e472de2e57f37728ad9317e4c2de7bbef4491623f02145aaaf71455081664e47f8c2900d8e9f71e78219a2180fbec1ee343ba66ce938de5d903934bcb690f69a17a7a668c6ede9b5f743616474d79e673da73dd79605fbec834f9f473b35e27d2e89b7b0c9e5eda8f3ed08c6ffeb53cd944612ae6f6429f331b27bac69aa96653ef9e6eda791b50fb6f671f2c61905ea1eeeab2fd7471d27abfb98fd17036299d420debd2ba60be24899c4c4a094d06fa8406d051ceb696b36802bb50f42cfb5dd24f9548516b50509af013a8f49526545997b664fa37a9e6548515b551e887b21ac29ef14b8bb7a10d6abafd52863a02a005db534bdea3931044904ebd186d717e83bcc45ea9cc6cd782bb59ce1d9e46e959753f36d9afcacc2de1ea10e737ec61c0fe1861c7559116983e48322b461cb8ef0bc836e7bcfd4491e64292d494b1f9a0fa0da2408594f61e40100cf844052e5cc15eb10d35a6d723cde72bf0bf147f8555cec91072359f831ba99d6615b581b5fb89f20f422db4085408b870e2e121d50ed1783774cde53d5ec1c5edc410bbeac816504a986fa2ea607d94b584934d2d0a6f68cf867c0b35296e654817be6dc203ed3bf006fcd323210fbfad383c4aeecf0e0633a9eb35741131ae6adae780acb1ad9454d05cc4dc71b7f10cfec34ada6334b6eaaaed9306471447ee75bbd565dfadc48b1804450fcbd88a133e5ecf6a5e93b3ca9ab3c6285e8276642720c535fcb302b906c390d464f2da718df6f3358e50068b377d2bc2ffa181ed2704aab4eba47bbfad13c79dd5a6c400b2053fe32ac12da6fbf12a5866795db6585f7461d5bd83a04f7fa574ec3d383608408698ff3358b006d4c16cb673a7c91891b86b199281bbd826746a878234be839ea2cecc3efd85d9367fcb98cf6bc212d1c8c441e0336c6c9f365a89b06447eab79f84b957e88d4f4b9c094c411e8dd57201cb589f4ab2b9dd089fa36ad6622a7c102a9227a2824a50cc39da0ccd47fc335fe66c52fc971799833b61020c9c46ff25ecd8102aa707806b4a460ca4c9221520e3fbc9e7c5d77d9b13934dff5e4e549f5084053924d7304ee531745355a549006189bd7e567c2b87a95891899d6cdb5779b6f46a9989849f4796d6077c98ff594f9f66a403e5b7286c2c7e6d0dceec06418578d3ac9b91cd8a0f72a9c719af4c5b055515d49868344d43a34501879e846da7d985fb8b6b050d60b77a61a01e1127967cb4559558dd4a483f86810584f75a14c313b0d5e9b3fac6c02de4b79b2fb2655bb35965846e7a236403b1f84e65f22afd752191cce2eb891c4215d3cec9d7f97bf29b85eca9beee25084d9a6850c61c6e894c6bfe982db3c282fd5874f21175a15e3aed87454956f071e95a1ac8f9eda5262fd93f5a27c4f114dbd0540e21248b264409ce80b53c7b4a9d254705316d9242fa90bc210a3e4e0f94a22f62ba90e1d498fc6bf9460680491003d57cdfe7df75948303ec49f0df9151970183032e1aade6349b718f3a90c9476c81b391fec59c7d4316a215eb2dfbe679f993c2bb2f60d2129a8a251751312d48d260ab857723537b31bd61f523dc254217c1dc1e8c92eeb24e7226c7eab4a3e9bae9e5f22e3e311f3505f8beada5ec6862b67f20a816b843459458362ce827b165b3b10d03335c316f1b99f6d7707b3ad19c33f56230f17173df2230a5b088949b56565f57048196b6124cd78a256c8b55121c6fdc21d8ce2fbdcf2c629f6c4fbc9684840432e4c7ef26357ba0a0dad06508133a8da80c77b4412179bfa9b1b9cfdf3e80479e08bad931d0d2b0700134898788b7d905b944303744c8fd3d54953186adf6acd0a90231049c419b691a6d48e7df2fbdc0829738f043808f8695d59c648ad163fb68d8737a40957894b0ec7310e9a0e2fe997ddf6cf8cfd86ff51ae96dc314109afa09369e57eef2c5686ec3f3a0f825d547fb1b3cd7c1ef07723e2208163d4ac3f025c02d4eebf6ec386d991f105326deeb5838222dd3eb8bd1479adda50620baeae3bca990e5d055af75011d196cb7ae9c1a8abe7db426422e0e334b3ee961a858d29d392b1962393dac595fa0a41b71667cbad178db13c50e50807f595a9b84a29d7088fe03e382126976325a52bcdfcb9a27298066f78a9d11a8889a4b13e6538673045bd00cbd7cef6afd43ed8b0451df569d97a615d7fd859ea4fc467450a5f41966690b2902f144e7aca9dd7496f883bca687d98e25958fb4c20fa5cc6821acc47c0f926d60c7f645aa1bfa413c7b784650890dbdeb7d541e95e928be377b3612c39f370b298b7c4be4f5fa7b61b2a60f91c9906a7b1a3ee935de545ee05c684f29f4da8afe18908a072909f00f13883e15878f473437252e1d2d238724392373e6bb1d26457aeb75a2bbedda0db7cbb58dbdbe95b2e5f28fa678ac884dd9e3deab811392490b6c15d7a328272cbd108f2ae34636bc601e4cbde08512f846db2f367547b9ce22592b6d5662ebef3a4226cb1c879188f2d666f0ec34b1cb3f5ccd274748212a6c5e01bd4edfc668e3912ac5e548d0f679a93bdd21f5233ff5d0d5bf8198eebb9c8dd8381d9dd3da293fa035aa70a42d8b311294107013083f90a6f8e86135ac3c37f9004da8d483c3d9b872d8e78aedcf2af0de77131574dae474d5cb489264e4a03dae249a48dbeda6afe0f94c9167a78c4f41195caa3652f9a264e194385f064fa81b9664b9ae2de9fc0cb5ca7a9d81d3861f7d45a1f2056676931db91610526fa3e4b3ce1e67f56e6904eb39ff3b1a481c67867f96d09230f4c4fc0b80a461bdb0ed5a9281eff11cc784af068ef23912c5e8c5cf51802c9659423add3c7bea5583cf64561fe7e24f8847e43e7a6929bc99228500b191711a20981d4c430a3b8bd8ce7b6a07ff29b13b2e3bd13aa2d915fe0476f65d6b2242749757fbd02797ea0c79e7a9ff96622e4737d980458f75525bd12027abfc473ae6cbbf48af4caba8359e6b4b07b25b3b64db58a2f48075298c6c76dace8aa6e4166e8dc970e6979976637cf804a8260c6315a261a2dd5bac98fbb32be8a345fbed5ebb4b09e6b1dde9976f4bc7c935b499e161c3c99b2aeb7701ce36e80418a84bcf80a99b6525c83729a7928e8f2fba0760a5e7804860cfad3b833646feea67d8ffef8c8a1a91da6444131a897b774f23e86d674157be3dab53cc53cafedb4d0c00b496bd62e0713055ad5d7394a67bb3af26fd7838172a82c4ed60bb3a7ddb4e7ec1e1e64d970c2acecffba2de4e35277eef62f955001a242b060c0e05c1716df2001c463d4a065b29c051729b598e889e7db283eb5ff7d5422625261390f072947b00a9f10e58954daab320fbd82e64378c8e3005514fb5ce985d0a4139152fe71483ffa74fb1c740bbf2af6484de1dfe70881e2ff1d6ab134292b7dbaa26cc774a0febb1a069ac831c437caff3166ebc9fb5f1682bfd325fe87853a26dca61b5b2822200d8042ab9b9928476424d420d1c4a5afc5bede66a4cc89a751e544a74ccb9838df69cbcdf5a795c6185c69300d86b83d0a91ab84ee5eb40cdc0b824119b3caa2227e23ba2cb0d49d8b71ad55febdaaa520607d6b504e23e28688d03edd3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1396034acda20f9b8b5fabc6c6d24fa793ce5185062418807e3211521bc98e609ef1ebde9e6034fbd04c249f7755e89ce7a29f22d26cdc2c4a83c18bebc60b7555869118f6b74f23508bebbdde343d3b75dcc55c5ba9c0db00bcaebfc8e7c25d342ef4ab28091fbc64e839e9b93b0e84790053078d66ef4444e5df5cbdac9c0f319a894c24900ff73e44461a13d83d19cf9755cca877be35fcc77bd550f809e4dcebc38f630b0fd28ff71b97a52cada143fc264c8b55515747e2105472449705c3d66b3f3fbee5eda65c1228573db10c23a6d727fa8b91d59d07ecae089b834c2712bcf92109d6847a6b28dd2a8f3af18f0a344d10b029126a060bebefaff008e0a3a656e47053102a18b95c3edad1f571731218b3e14b6b0e6402c3d5d0c328bc52a63d5da5f109d1a33b2d032d6bac1754d6272247f7ea9f01fa9d58a01d0e09f4c6e933663b5948f2e84e7970a563c58e5dc56374c42ebefebc07ae19c5056fe39cd9f17f8b69458a01ea1d9228f93b7e324c3dd2570b198c3d7af61651f8b03d2a96971d3921b4a7024aa5a50b72c87e609be49d2fb87e2e5974ffeab35aae7a6a2e000b569a31e17b580201c2627313054e4c16ee52da200e814e152623cf51aa2b6fe23a06ccb515f5f4e64f52a871f5400685c18c7a1337de8954655a31de59e7810fc6b68347e221c809ba81f9af4c4ba83f2007b9a864483c73e4d7e274a0061f2e1e3b2350e86fe838b57931828b3ec7e1898787490372144a3964b38d2404f04a6a95e949dc4e9e9c134de9f7d0d318ac4da9c2b31f0b6ab1551d744a1c6bd0c6ddd37e6a5d3e1dc812badfc8a46bb536697e8fb632576f76be77c134b27a1c845e487dde607248ec11d9595a6f8517e3cf2871184e1cc9ebe4e0f09cf0d50efd1e20456021d203a1ca8aa06b697da11747b98a34fc34c30a23bd8b0ed4bdb1800b308c3b551912af39e600b23a1af08c446491ed2b6a3778ba0c38cf96185c32db9f37bd78a4c82245f2cfdac9b0b9c10903bdb95317c95cf9d212f65e795ee097870c09a322c77783eafc9a82a424f8b58081b99d685051e1e77aca1cd5004b997a1bfb10273bd6c29ae82f989ed8c6a12b604fcb9eb71febac664d62bfe7278c6490ca81a77069f639b08b2f570dc1296deb9c178fd4e6faeafc6100f5465402e48252f8d9b5f63aa152248e038df85dd4c10a208377eb6728c79a06a3c3cc85f9a8dfe1104769edfa910470e083f2142fb9b6ef49a93c06cd6e7b6173b594c96905f1fc56e013ef776a0df7f10a8648500def407036113cc2e7370f9461d078fecfe0770f4aaf4873a8c0c58968afed0437500f55c08a8d47fcaf70a736fa4dd0beb14bce30b576f2224b9a0e32f80aac8d76dff6ca3628d53d185d0ebd9556481864d840870f4c0ca6ef937411eb5840cb8fd50c54b93bf821e329fa4d0c28f8fec2835ffdecb9393a8518559d50e5468df064e22fb13398f9ef259d2c8cf0dbefcfb759b0e3473558500c4c76a4549fd389f7e74a9f1ba82787fc0a239b2d62e8d96cdaf6e84c0c61124e8b95da1f822e7d29b360eacabfdd1955f7bc2664b0650f4ff927d37d67c679906c25b50535fbc755787efbc9007a3cb03d3f83317eb298111ebeeecbfbf9975c9ed02d250a07371e4eafcdedd284a2310d2641a2dc164ed3a2a6fbc570afc3e38ac34d7eb6147d1323c207591e49492ba096055b871cf3270743a2d0e29c9ad0001b8d1964c64f4ccaf344d8591a14820e4b9ecd5e4af8fb09cb6d64acda11bf4d5449891fd4aaadc05ca12467c3cadcfcc5816b04b7a46698dcd20053db6096448ba12889402ee668d588c5466f242fcc412e4702059c2998ef6f8ddcb23d335bf74cc1938894d5eed73790fa8273571f6e590f87e9e3b920ba3bac9b45754318c0383865c3be0e09d500341a627c99e48de6155664200e1d50c32209df8984a0e5e975edc248acdf413373754d963de5380df748244a6fff894742fc0f614e1a1d6a92663882d781f7f2ef650333bb181cd502d21ed8d722a6765ca4201c5242d76a25929c9bed33047fd486293b277ba34ec6241555a78f3f356539ecb9bb11ac282135f8a86ecabc6d0e40238ce5df216bfa281142b37b780bc748b7e2a87ac97db452287cf3137a9743ba9c6ad64532ee6d9bbabc882be367a3bc62cb2d60efdfc389c37a94baabb12b536bc0d314c9fa1eb429e3e2bf8da923b45020774c9099fad89382c6738b40908a729781830ec7561e6664f1f893673707cf623856c5c1688673d7bf6c3ad750080706db84defef120eb69d46f06d442db1e52ff239f224efaec5d9812ed1fc2ecdbab2acd7381cf56dd511d2bf41e6bca92bf580d8d37e41685a374db8c1745ab4ddcf9d612c762ffcb9320b18e92aef9e3de7fc1dc9c3c587d1b1391a3eebeca89c55135f8616b191f597fd18254c257ea9e46df1cc4ddd53ad7271e289f38ea1a017a2748bb6a7df0c5bf5d59c08ed388b7dfbf12f90087017057fe7b0a4289193f795c215d638eb2d8ccc091bacde8c8b2947c498cac3f3179c12ee443494cb26118334552325ace03101d7ce420eb997e83d2866759511542e73af16c045d92804969be72b780fd3fba41ab804f6c402826005fb8281f1d7994c0e08cddfd5ebbe50e3750f5385e2ae8f53fb1ff393b28ffc6719ee1bf83a14b0aae937697048eb10ce2dc1e8ef8f8522bb42ef2e525ee13ca69ea4e02c69cc2b03d903d204c69c1205e4e45d8f899c4acb75b6664a22800a2506e8aa5fb1889f0d1b7df331bff3179438664129cb2dfec4a42525ad9edd1f4aa5a221111c836f0dbd713b727caa941c990f2e01701d92e149f4eb289dbc225fdfebfdc9fdd7213ab9afc66b79c083da72e056398ae4000a39961c66b02e73971cff291239225aa34c42f5df7125095ed48fdc4b0b77483063ca9814cfe0074e0a3a58a8c506dffb1000ee9e200068020fa2ae942d5d19fba762160b1aac6b714052b93776771e135afbc5525ef81474fdcdfb23deb8816ca7a9d661ceedf0e5f36db8a8c09ebc40103ba21d8dbc94ede26b9b77367d0ad47c1777773d1721c8016bacd7e65f3bc10b46164bdd87e37dafc092284ea2fe6a6843b97b5c848768ba4342a96eefe5722c67f05df53939380c48a496b4eb07c0b19570c533e440a26bbd79a2d5cbf07defab4181ab601a441fb45a3e95f7c3899f78a03310e017cd55d2b7bb1f1996fd628ef793fa294cda7ad691e2b8dec0267a354efabde60a243500ae7a86f8f8dd74a259532f65927fff8fd6a482acbf29b0c5b2afb9ff5f3ccfc5744a869c8125977537e73ffd4f376224b81b2f963afe50ffcc0cb4dd0f89fec4cdd9e509c9aa3c0ccd3c33930fefadca11e567f22c7204ddc08a58cbbda1c9eb312545ec072941bbe136274c5cbeb02cac478d612253897f61c69c6978c242bf214195211b8a92b554fd206f755639603f404bb1a7a0ce914050b9ab2e99f2f684f34406a5090075d38d09f962562e37f7885b520cf6cfaa35e4fa57edb3bb082c5653003955d00e3a6186b252f5371f81bdd6310c873696397159a938209c486e8f6b874629ce61b668e2c92bcfbeca773de3d42b53c577872265c9b76e33ccda6e609bf6a14c9c6ecdd8efb135759e6960bed2db1f8258b385106b7ede35e6af9afa15c6c940728c2c2b8b361cc425eb0c8a43fcb10c4610ae6dc8fb9971820ed697f483e26beed4d5b492751493dcbe441679794ed099f2999daa036433d130d2c73c96dca101e7c8556725d2082c1b65bec133645f5a379a094123bc2f601832f2d74eacbcd1b2e70c4d2d86642f6aeb5b9a2cb889472d5b355a3cd482ebde34cc52406a453847b3b4c6cbc52326929becb6cb37f4a0d8a1c5739eb588e339d6380b13abfb487a2ed011ee6212bc91979ed5cdedf0baa187a22f90877b7805b454ade68f9a6add4321c4c59a31b92add239dac3e8cb00ef443bba6c8e443a93e2d606dddef8a480e7663fa62e53131fc187ad0e8451853e8632db7d75014528830c665a0f07f9afa27649fbd96a7edf505fc466df3ab19d774cc2668502b0ad33f0fc511ccddb5d4e97aaaf06fc14ed4082d3f3dab176577fdbda5e659a59d79060d0f7972d9b8d4967ad3cb1ec429c48388295ecf585b06be0ca541e99abdec7f68b48cd71be1d80cab85c2e2c97d746d8f2ab8753f9f5289da82456a79afa96651dd56215dae91ed89dd2cdc2dbfff03243a03f36e7c200cd4ff7d88ebbadd0b46c7bdfdc16ca6bbac16a6533a5653ce5894684f6ec53ed7fa622eefbe91e14c4577535f5b0f5f3b5d5c5035a8ae04a98b0f611dec0e04a7ca8139220488a420f571323a2471267e0a83dd4ccacb19e1f38da2a45e89bab5b355aba25516efad0c4883dc7d0cd10909d3f9c6f46728f679ec675a8445b3a875a91d2c8404702482cf1d8cc1860c3f3cb46150e5e8252f6129393b95c364d345b1d41fd7c1093eea89d59c1701bec292c30ee005b7b299a22b3e44668f4edf9f312b44ad94c43e9098975fde7b955ff0f7ca815aa21650609a4e69218f6d54b6de120546575cc19041eca0552c64264729ff23c7e980d008b6a29bb39993f29ac2ef4a7152ecca4c2c70e1b1ee5395df0e073c7aba4fa8103483b280751f23334acd6162c57ca0b8dab0ea11277b58b196331474391ca13def8bb62de4566c9f73a55b735db5f635ea4d9838bac734d76f0fd07bb7dc001e5851f12fc10567d210c9e8c684afd9d568f271dc4115e10cbbdbc5fb8e8f5068a470720728763e4be4dde8a7629410d0d67b97836c91e6c6d86c3b4f312cfa9f08e2624fee40eeab7652c7e4436239493b2252e5dcad737da167e80bb0791ce54e2b3b8806a2af151599b3d8ed347df783804483e3bccab82685ba33378cf23f58176d12acdebd810cfbae57f155ae7b3ad9a54d1df585d3d108b0483fc04043aab435ee9b791d94f35bba854406d1f64bb21df9bcc41596777c6b56617e38a5806251a8a59a5d26495568eeb5c3802c50c8e6fe8d919d46a70716b289f4410a76cea66d4833154984982f74ded815cd781b33c5e87a132f60a428c46039f49f5ae49b08e094820c30c50563b57f1bc2f56ff6d62ff416616849206bb26bb50d55a3893ff9857added92d2f28e0833f1650d6d3eee2272a99d7e7bfdedab4a7c86319d2e34017dd672effe43d2fafb228959284c3bf5b7207f83b243a1ac35a3920d732a1fc4f1f0730a0ec319172d958ece1d9fe83e61fdd8ccdb8888eb64d21f1ec58f446d9c4019bcb0ccf6b26802fc50fdb1f65b688cc3bfdf9a58d777de95b9b8a9f5bf9b2a82c5a1c1ce9de4a51f0785182e03d30a25700bf27c55fe8a7ada461facb8a1b729bad66a33f3f0debe05038991d378a544a0a5fb3ddf32a91c1a9cdea341cbd1879eed33550b56a12b1b055940cedb05dcd21d1c094617b340a3eb2edce6ed1065132830d5131c2bcd3783fb91297c9594f19f946d1213c5aab25c2b3fb982b0546d883d25939c79a215f0041284913fca293e326a7e15cc426ec2704d650cc8729688c59899df6f97e5b0b752f9fe985d0d0983ccd14323feb3f2dbce0b8ecb1254ed627b52d45c7445387a63d0597e8619e41583e3a30bd53f9641077aa8c4794265770965e4c3e0cc15f2309b8f9ae84ed837947d5a325fbb052eaba2d7bb519199aea1ee18a6635787e9bba92155c0f802fad8d3b1f3869fb2590a1d86437e108a2b81cc897ad5412ac0c27;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'habc773d362acaaad6b684c0ed2311d90de6866ad86f8144537c9745da0174ce9c84fc63cdbf8f90cc3f2217b2c9ef99cc442c8337bae9b55d5a155bb283f7bab78a56aa15b61a4ab9832ad4976d30cc9a4fdd6fdaa7023231159b3eb9b27629ed68957489cd349bbb99b3cb0114d4441d513d1e0f4633b6c0e310f313e0a86422966f3982b57f336cb79bd088de39b83ab1e82c89783b9fcb27ef585891757cb63cc3db471c32a8f6b95cca191c48ee71247e90ea79b07da223d6ff319c8f0cf639e4b2a440d1ccaa32c24ca702254caf9523fb6e52404ec6887fb785545009f765c8fb7c65c5b888e4a05ee1a3ebfb6d473e63513e7e8b0ca36b50650dddea40b68a34d94fbe2f364e0bb506c70c1f1e74c92ab9b519eab6c0c9890507c7b66b6d708b4c648477d88a5f8dbd1aec4537ed512963bb20144d697c8f76ba90deb73ab5627eeec68cb6f4e8db7bacff4062277b403aca1d0d98de63bc2d91aa02708f13d07e451703e6492e21ea002cfc9c9e0c40f05aea87aa9ea876e45657abb5cb620cf1ef094df97525c9fcb79f0bf66224eb406724d8a9292347875c8b50aaef798aab692e9387ce78af64438f64193803d2ca2a37cd7113025958ec70ddc89f9108c07dbb5bc6bf938eddc6856655b3bc979e994f6bb693292cac12a22ccab080addd60610f78dbd39efc1f47ec414794cd463641a3d5b3945544332fe6193968e14bf8d46e5c17e3d11c5322216a53fd6a553170e87734e98f2896b8501f577945dd243141b8cc656738be2ee5b41fe2c3aa9fe279ffac66869b88521ad1a26a2213b7241231dd878a15795b57271ad51eafa5c6d8681d191ef51502a6e711aeaedb7429dc9ee80b5c3acfa76d2ea568460f22ea65925c77ac30c27edb1d334b5671fe86e4c7dcee85f599aacab871f53c589461fdb9ef2c6e523e849706b99bfcf854a0dc8b148c854bd0d0202b1d1d9f40d59b854f71006eac768b28d7193df9edf1d71613151455ae0a88940c067b150d1f3dcd420bf43420b3fd8cb2395fe20a6e137649efc5cad7eb959f9050eca7cac0d7995c0ee346d35ec7ad3ac4f7cb4747d259ca6fd8089d03a2060c4a8820b4d54bd835aa3643b2a7dd0daf0b574b70d296bea5bd6486b3f55820de0ac27a0e27933eb5d2564ca74981e246974df2e857c0629d48e00132812fe9e0e4707a652350b3984d61c20a3a516e4b6b74fa1f185e3bed7481decba7bc4abafec1cf6d6b04ee6cfe5d49c6b1cfc1960dab535570825437de8ad4bcc09291adb984704ac77aa2786766007e20598b6328baf83394c541299a7a867d769c22de4d47a54efe0bddcb7b3a1246b8f0fb3c2468d0624d6b24315249dc321b659371c45284126164c9e29476566b0a2ad0af32e50643c353b8f8d79790752964953bbe7cd97ccbed99af707da47c160f19ee516c39c476233da67b0cfc5a40c399929f1b353da5116ead82687e819691623153cb8e04a2ce9e98cf400bc867a5b5a9e3247d95b2a45505ba16115850ba7c168e645737cd02cbadad6d360515d9dd9564bb684f50167e437af935826086053d852c70e6a544fd82b1b5497e7ece12fcdf06ba2edbf3909ad7764d35d0d3102a87e9d8fbe0b0ab5fdb7f133cff862a73aa811d98ebea042660b2028f21d666322b473da3d94a2cda828dc5abad5fd5405a05c022af80e17992edc7c88be9ce96aa8a077d50c46c1960db06d84b8e1f5b42086d443fb57c7003dda0f87cce6c86e05dd30106b83a377556e8ea841b5d6051bf7235aed24c6426a9b9af1e7e3589f0c09df26b8c964cf6f75d3ef2e54f52fb38b072f1ea592b49c393c288efde72721a664bfff4dd5a631447dbca43796760ee3eca1c133011586fcab44325f8abd867333557a19b5f0a7e0a47d2de2eb87d04a0c8e012dc4803029f7242ea33604f9895a5c1d4cfb0dcadf03f3b9555622fda3209fdd581b62f7720c5df7f6a6bc9f94c04a046ab490c29a01a244592f0e196b33d18c568aa752c6cdac713db77b483578316af8e100480b7e72b6e12199ed3e6f5fd4f0e11f4c504b0cc5f61ba5ba8968a722087dd64df778a786a0ff1b5078c58286c51be2356e8bde228ea8f2ab981b966021be7dd8fc7e1eeace481afc3bb7e761a64b510d6e0b5af5f841e36bced36e5d2d8c7b719e466ca537f90d45fe704723beee8c6a472e0ab878bd022e262b0fa8960668c13d3f8e2e31bcd0e02112dcdba7dc0ce363830a03616e64a66d94aca8a9bf02b18474d5e3d5cd1d21ceeb0540a6e5194eb8e622a46b8bb46c57803d49e30133256432c539b8637aa0cd5904ea710a097a115d7d33d0c2d3031e8e2a92a9468318551f342c158a43b47a80b7771cd791e2a6a3c396fddc16d85e3ac8f1b50e843e30b290ada3fcb303978578e2220c4bfab2cd9c4fb9a1ca033bd6b0d43f73811a7531759f4e42febae72c442753ebc016ccb776555b9f45364407f45502dde7542371e331b9154bd382d4d781fff1e36c15d3caf2d58d53e97d591c2233e696f2b62a647756f85f2922bcdb3ed06dbd8863b0a0703f1a91a5acd44f1b6541cb5b4eab039b9e1e37f38c029a7aa1ca8ccf482d6ed590ec02ab48359355c23c2eabebabf8e1f27f9efed2daad20f76b53e4867eebd587ab1c31e330056442c7522720b4096587b72367f817b89fd89e7e417153d3c1313c89316fe8c21ff04e78ba65e1ee11d3a20c125a474d90207e54fe38f0252388708120662b5b54b3079a9f8ccbc8abc02d5e79e0b9db2b1e1d1e7dcab8abd75ba432f5cc004e4d651860da8857f97168ae9df5544fbec349d2c42efd26bfdb9d73ed9ce14c3f896e3340d4571b7370208beed8d1cb239e09bac1d2340d86cb18c2a912771418d370c8d9f67b37e6bcd9ac7551df3f5ccc629550406f75ceda6fb9f8edeafcedee883a8b8f1075dc4983034e14b3e22b732b7269a234a4dc355cc6ef7cd08581610eade5120afd836fd8df66e991761326379f2ef4082dfb6ce4891925c6c766f2c0d8fce5138baaebcf2c5dcfbeca72836241bd3998193776d72c6cd6d82d268d1b213f8542f54061414468ccb5d37c9a8d72d0a53f0ca7021d995bcdede693039ca266c402f0542ddca8d515fd2996c366ef7830afa3333eaf0fb75e91581e58b71c8850a0879df720f936cd41cb7919f5de76bac505df45ff497cdb8caceb455c8a7112519e71533cf1ebee9f75e4862a5f19802545d8fc1cf0895e3b810c5dbb99cf8d7682347cc7b36c791363c0d6f2489f971c11d236215c9983ff6d7695101615255098fb7da6e270431bde61daa3f0fe616a33ff6ee6b56d9bd60f6037b85b9bedd44a4d1ce882d22f2974e85a7662a6dc92e9a5ecc368c062f6246adeb34dcc6f4707962d8865fbf68292e8783def5fdc60f3f09b02e39814e31054122a43de89ad2f5e93619c3ae010bc0f38995f1b8a67eb5b118031c0ebd371e9ba2a9de22d48254c521ddbefcd26b77e0a917c3bc096c66a75c5fab4794a57f2657945ca0b029d471c90d412fdf30b7993d0ab1e4330d5d2a7888b55787c6bcbe33e3fc6ac3e4d958a6d160f6cda08732f8a817659e5cad2b7ce1a5d68ed8e55e4b0d60e52b581793d601db4c8f7121ff0d9103f015acf3bb10bc7cc1a2ad712f917f904f1de148a900a6013a4b7a034ab08470f4bb6137f8c754649105bdc4e39e4dea3c420445ccd155e092b11bef83f616df9bb7ae250eaa8bd2fa80c3f87c2935fcc516243a4f4e70588c8b2deeb2b023d3030425d19e212eda7d04c593169e3827038227ed3a1349df980ff0d36641623dfc5d8dc65607c31a3e80cf9c3906251fec282cd0e62e25be2bed61d0df09d965a5c568c5a1f3d9a88f929c3faab1fb3f455381a5b680e7076c793206e8afc5502c2f8f1c2313dcd813076c7b6d6291076ce82ad5fd072acd026ccf04023dda8f48753ffe2253ea5cd42099a8ea75813df93641c7e96c9efb79b74752b4d3656581285e2eb9d021d35c8db7ebeda1daa4acfe132facb5d0dfd9db87d5bde174bf36e8d8e139b0ecc91da8b66cd24e4e74166a5be5125ad3820c975c7ace83c572c8cea22e17ca41c18da00d0f1b0f8039bf81af49c7ec38b7f71c514254502a78e4645c3e0aff48f564118758ea1cb94542727120a1063903c375febd411e97134b080503fa0bfa6e67f4dcc2c4fcad8652e595b59bdd7ccc905c347a0c4546f5f5b4dfd163b7891e6aa09cc8ee5bc65b13717cb586d05992f82803051666f6df446b5ed548a343a0c450a3c9dd032cb7074f2f9d6b94c70f918e49947d775bdb8a034749ec1ad4e912aad176c96a5ec594289e0c8fbfa7ccc7c1f4cbe3c1e6764579171835887649b4ece63e2d2eb5416caea7b907d6e1e0a6080af3dbcadbc676d848cf9ee7d9c9bcd1cdde763e05e9dde8096d08eb5012969751d3a50d6fe3de6c3f25f05637c5d24d4290a4e034b2a6108fec44814ddd982f10d2068237f8b9f45ea89a9cc66cc4acf8aec89ddd570f13b108f290c9d35bd9a88be875b5ce32c45a7bd70380d7dbc4f263d8958357e82e50857594ea7a4200039386a92e08178d5bc3e67d0479d9c683abdfe44951bd2790cbeb3a88f00d4d3133e51c5d6b39b4397aee97c2044c5d7fb8b464d8543f420aa3a4bb5611326a38fd052b49e99371835a18156cc27b90687d3936a53d2f36f7e324f527b40bf1c41c09a6c1d82ad236b0ffd95d4fd76db22e1ca34be7d104b2d7cc6e45a3b3e429c1be6c9fcef43fa5365de5d2912847c4ff27a86b811ff00f89f13691f7c816c3d6f858fc841e7e26cfc7f7ebe8de1af87a7a461dc25c55922b14f8423f6aaf84e8b3c570cfc0a67b30a7e31be19d60953de27f449e69e840e7c7f3182921aa6dbd7ae4538110696edb9c05ee13c4aac18a9b9932f8c1ef4ec977b4a9ac4fbee1c036de6d72d59f64428273765ea400d939df75e1b37a7c5d14c06f0ae751a48fd5fc5ef05fdbab957728148e3e33ee145855b06e9a6a925ed5e3d56152d8aedbe24ca795f93b4eb29c0629b6825463029441e467aa87082db42a2208eb7f52762832bbc8f4642376e92cd77a8317d42be20b5dda7d4a5a57356487cce19ebe984da7a36fb4f584ec02e42b7b63c7afa349f3ccbad395c622fc8a8cc53d41bd2c097155b135c56b57057bde9a248da42a8fefd6a4375a02da08ede6f74a018e7f3ce9958a338d3efca5ea5a808ff02e0ceeb98ac85b117615269e673e4bacc714f60de7eff5158a9d6643efc411b6c5adbe8a69bdcaca708990ffeca569f704784138db5e7c405a46ba7be97eeb725ba8ed8f3c684971b15e36155c3b0fab2d42c2e70c9fc1061dc12831504c87250698a0e2997c52bbe2bdc95bab5304145a52c9decf57a7ef675841447032f4b0be3f76d6f87e3db339448b45b0bd632588eb81579190d2f28c4964df5037ef326d1bf9903335e53ee9840d55367f42d8b9e84ae6c57f6c79fc293619f52e2d331ffce90f7f73775b8c3faa12ab203e96fad12cf463f17750182a71689710df1e32b13300b87d6510de78c4f09eb360d22aeb2847a67100d2d74efe079af8bfa600c0c74a51b171263430bcac87ba5e2aafda6e6485df88f8381198082e99ea18191f22be9ba08531b9bab53a539608cb814a346a410b7feab455b3b31bfae43d4db4a9c4c9805cf61927966c81e1aebef2832f006968f5af63a4655b1cd2009c7bba0aa77087fa91dbf4596a778b26af3d67b9a1dec5a18d0d0579ca805e4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h558d99bed51851df2811a4dd996e55b1fe6c7890e686072b5fdb8c5db53773b0a3ae159a02a5a002f736045a829f6ae6e780feae4a8ded1a9790c255d4fde3db729f974823e795f75a8f5b8e19c00056e307caf6113667874ada9453e179d46832ad2359b8cf22a8c3a3dbd52ce541d37ad2c289b8cea8e144bda372957b71e80b2ad5871ec9ee712330750de68e8744d02c73e06c70974e6b39a77fd73102f8110de911f9474d05ef3706bfbf698674436167822fa7558d0f0ab24624ac688f481b820775f74f4b6010a574d99c842f35cb0df7525e2c6c5e9c53f349ee5283183bf9b2cc24a4e116df6d7ad020ec06285b66d30ea051649c866c902bbd2ff56b0045f9863f496348a76580d934f54b13a78c467c9f3d85441022fe207ffe8863b0302b0162aab9a9d48a9960d93e820ce0ea3bb88d309f7886876486c08d5797a82fcf0d03c6b0a8920feeb205d24aaea9855488cfe0789f0b225c4423a7a2198e7fc032ed1222cbe0bbe70c3b5fab679518abebb8e837bed66704995ae2dd20008f4727220fff9890c83c5e6ea84dccf8ff0994aaee20ae1bf644a6c73324788ed90e1ae8fba4625dbf242f70fc9fc66c56b8d206667ab528ec98ab13bfe6dbc431a7ee70265199cf5bc1bac80abbdeff3c65996a6153a5e93fdee1276c30a7f1c7cb7a04dc28f03e380ab8b6b8d6a8f4213eaa7f9b442ba24b9cfd69faf85e64f3c266a3f2bbee242d0564a7f3ba3e60e4ed0a063efe97920c9e7cf7d63827de3499f3a7331f39f8c1da2f2c16788fb71bd06396ed1046bf0c6bc4f1a8ab4b8bab2b2b7bad5f80481d00b34280926b3e0a619666019539312a26e03f88317ef5534e271a77d282926e730f7080657f210aaf2cd35ff31edd7b6397b7963af0023115d5f4775231fe81d7e79cae5a950198ef29713c9b1cc386bf0307f9c1da528ef46b235e15d0d27435e5fca2defca2bf7a27eeef293ec4f380e9d35f4ffbc2f2eef3c9a26031f3b5533c9f51dfb7c03c00bc067f26768ceb96a980b49ffaa2bd05154a5deb6fdcb0ef60361f0d107acd3187ae09ec6a525a1dc90975b3f281c3c24b54ef950c7f930aa0c0da6f7e84dc66b7a3ca7dced3e7e6f15583108b879532ff4874f9a12846d33ff40a0f0d88b67d3bac8a859c3fac8c0fa501ac93b38ddf5025c51788c2aa2c611d4536a71276abf2ad776d90749c1a4af3d2163264faa3a7e60fdbc50497717c7ccb45bbdda9d44a95e278453b04e5afac52ed4e344c42b9eed8154af66330ff8b493357c76e451b4b98538c3c227e00ce29e4031e20aed12fa53d3462c48b10c0527c2d34c894aeaecc6b72d82b25c61c77db68a31c24fce985d8ed059824a087580cecbcae56b935e27e1b86d0fb6b4280d1f4da18164ab45ea3652846e2c5a8531d47225889a6ad4657645d8cd2bd6f8a54b415aa96adba739e9a25e9c3af965d2994907b04d2962bea8570de143ee20ffb0ea69039335b080f4c13039ac195f3cf754c03253102a8a27cf961e33c964d59df291a2ffb2991fe3f752d61cf3b4ae48da4e16b77664cc7fb27a1e75610a655c7012053336833ab5d536313126b35033bdfaf93f3d176af6886f38f5f2e9311d745c076d7749ddf90cb4732a8d0fda9e2e3dc9a31698d25ede64f4f2a023c5467591531458f24537db0c6a1b8e5b75f4740df0327859dcb63c500543477468135553929e5dc6b89f3745849c58a8fa5ec7e21ccee057b3065372cb25b7a28259863087c48cc46841cba804a8334a9ac0ca1d2b22a923eb7215649403421e7b365d4601ea3f26c93de82ffba4f4d2081d46bf518b4ae23d2b1e987cda01ffc45454ad5362cb940047fb321480621bf63b90d5dcd0339eef8dcd0a18cbe3c8afa1e4056bfb7c735c48f77e7ff150b6cd2290bd3fd5c26169ba149d27d7fb233e2ab360b81ca4dfb78495393f7e1ac112e663cff57fd65c29e3b64fd77b1de3c531f50dad5be9af7b3b814d281f92978625b6e33e9902ee24d0c2363449931c4172d30f4c3e6aae1f3e2803372b84e47c7752e6708526be54cebe60a65d2c3281bd40bbacb7e7be46c5ead4af103b6f3f7580a1601a6af6181bda8a0b990ecd62f1ca091e9d8665e2cb1e7104d11c22ea05e40709f27965fea4195d7c44a382453176c513439fbc6430323e5148cbc166723328a2e5e32acb076ca880bd9d4518a273711e1e17fa36a02990488aa4ec1e811a0adf7135f8712a28754f555c984cc719b87fec9fb7ec5c39266f94ea58796d700ae03ba1a578a7da6fdb272901f93dde27b7e80716c011f48be47721955598936f0372564598611fcf4aa9a0bfcb4297be6add03847ea1403f667dce5976c61cedd7c904e5f9ceaf1d1bd8230b898367735790f282911cd69a286de6815534a887ff5c9dd81bb2669773758dfe451f83f4b29d26f1fe49383263afd4acd7e6bc1d5c743fa2e309c8f155daf2133527ce6818e039c42a7390c48665305c04a1b7fd18cc4d98dc718f90f6d95a097cee116128c2f642b62a2a317afa52309063d2e47b3bc9c2095f8a6fa75233e85b9be96e20b19d3f25de21764ba29ae438000a5dc2dc92f5aceacb3b80814a80b7230fabfe0ea77934c8f540d86a7c4d3837d7c2fc907e92a6f400dafbfe557fb1f9fdfcc14ea25a8106d8ad693db53b85cb356d600ef22b1a20ee7bdfd0aea141c52e0322f6b15c6287a344e6f623f48cdef3efe94791bc9af871c2783773b254bbb75d21024f9d295c22166f4ead617fd98c1eb3ab0e5b4339208d21efcde4c10a2de8bb51aadda18c7cca721a570dda96c21409def4cf0851fd2a8de93d265414ec0f9272eba83e50a5b74f30486f05759e82e2a10df0c205cfa493181f16483da01b3dc924abf477f304078f4dd7ad7d970e535224e7e7f4b5dfa5ffebb4ce68ade41bcdd3f50ced498974273d16eaaa416fd4feab13e007bb8ecff31fc519a700da757199ab14e78386dd66e853e0a82cf70ea3dac3f33a4f7ef262c8c408097c680b76bec15f74234105e327fba1bcf8c4100abd52c0fd326086e62250749b7fdd33a61e0d6a3d08014520f17507caa0ef3cd7352d4ef050c7a8604dbf8b793a1e8e1ca89a8943ee2d35098facb8e89a771ff6bb620b660851b37f61d3c11bffcb6908444794e84be4d4fb34e629672f40499a6ffe15e503f87c5fcf73d8239a57a52520e9a89c4c07dd406a6794db1728dd4cba6a5edb5b481a1f6c59727e9023f859107382eb8fdd34d7c4fa02776b422cc74d1bf4ec0b1ec3698362a6efa779654fb52d97bd1c79b8fddc022e837e13d41dc7d3612e58f1dc087bfb8e7b51007637abf91327e9de34de2115625644b8176cf7fd9bfcba3f4fc502afd4f5db606c047ed26a963ec565cbb5fb2a1b4525e8c4343c253b94c1db36debd2bd40dd9d8fe1bf98e200424a1178a3210ac02b5fba3541608526152c788c2631c4ad3cec435e9dce0ee3260f774ade9031e170d785192276ec9962e8d34471ed047691e96c7c882713bbedb3de997c2366f401005495830ac9b6460a5eacc72758fde7e80fc6103db8381f4431c48c4214fcbdfd450a246b2f41e399e8714329d4d0c3b44c666b01a6b0d1b44c181f87f90c65075f2303f697d2ddc98b4dce897939673c7f64895121e6bb2c71b5bf8e18d266f79ad3f3c8a64ea1dc50c72e105b0ea26cfcacd5073a48d5d9f91133400f96bad82a040e78c0d53ed01bc55894279cc7bc66653bba6e7410237063d850ba7d1b9ad6b742a0311c59fa3543ef69ad61b708052d70da9363a74336547040a7a98210318baf16333f805d1fda650b521e8ee2bb0d89b7dc8f3ce08f2ef22391f771980a36a09add79a6885deb06e81b8044901f2eab3487dbd168152156ecb05f388a44c574f64839e40acd01ac213aa5d5b0836c33d3935eccfa9155d14bcbfd77c94f1d7bab28205c08637d94f733327d11d94bc423072092cd5f9080e6b8e00428cdf84235c3c30c995fc647129437e8736ede8d453a83deab16276ecc227dbbfa0ad952f5e801d36bc483c8bacb27f057045c6ad4cb088acbe0aaf98847a4da5d6b7dfab9bdde5cce7407db53e88ecfae1240088208eebe83d873f3cad1dcdce01ebfea9c275488b7225f1f6bd92cb1f1493c51b4c68145be1daf19d77d221c058c066417958f5431f388bddecb7084a542ce62610fc7102aefe796acab0074032856e1c67a922f17552269bffd30f852ee8dac2b6d7a87509ec8fc0ae282da34c431342e9912cab10f6e3a08fa9c419e69c1103e214699836ad5ceeedef6f192d776efe3d73271cc87b8f8e8980462af8e72a6ced91734536e1cdb78c309212e5320d32899241c780010c86b740d6aaa6c9a04cf311225f7aaa0ebb65d5ad55df6f0f53c6e74a23a3ea990835f6ba6b160034b9ee9240b6e1900fbe41f1f76310b20d1e4d298a095e6b75173705b318e486aec3e208db4fe15292da2013e77dc1a1051ef816c173c5a190e17808aa19a19f5a67dbd7ec5c47631626ad699fbdcae7e7020df6cea3fee3775eb39397b58590ad3b63adb21886247c9cd52b018367c2c288451e363c3f4a74e24bda08a93bcf6ea139d0a3c6a33c0fad498f19a101636a89aabfa2719291f32546ae1f80c868a3f49256984375ecd6644ab3c0ba5927c2ac5e19f755ef0a1cb665f2f109e9645b0cd5a9c29110731a2f203e5b4011dd0630317419275e8c995259520d31bd6b0cd3ba212245488cb4e58d96207bc286bca6053d5ca38f1477d8cce5c409b2fb13e6bb019e76a6391950be197c34b3cbcf79d8d94da26e698127781aea5a05edca96706d958b795d94acf438ba290552b197442f57e66c08442c0ffaadc2d4c3f6e8d286566f4686950073207b09ecde9d0b0f3773321be18c89a71c06f062c6f1372c144491af58eb19c7108047b56b86bf759b5e8cc329c36ba3d94833576f7194c12a1cf22f1eef2d77719b543e849135b1023ab7c871cc9a2825a50b5a0330aeef99bfb1d005f277ff9e91bb695cb971cb8a7bf2ab3c314f177b6e5e5fbcc1d0ad3ba70e10e9398731aeb4627d07609b15b73644423a848e94ab773e18da99be1d579f330c2dbb7e6db9ed059282836157a5b84a92e3e74cb81cf014d84b8f58e779e49abab034c2714fa5f8a7f79976918077198bc3f0fa82361bac389d9200e18c6ff77425a2b0267a2cd6f5cdd07615b8b4971498c7253b24403545d6fe87a6233314667bbe4fc195321ac2609e3678d8a0315c306deb3e58cb43f04a076d2b3d9039fccdef4929bfacd799ee2c08e3fe638868e3943ea66c9cacaa23320ad0b32108e2b3e251c1d214f7db3ec873ab175f4a6a8f7e7dd42ba60a7e006d0734a7d567e3d0e4cffa326d55d1432bff261b1952f4f61464c8549b6834ff431041893178af0311ed954da09974219dd2caf173d4d080f6c180a966b75ce3b7c009128b9083c0d4fb2dc92add6afd323aacb9e21afa521391e3794399b67ebd07d08ee333de86a5099b758afa3a7e625554f1968bc912ca42f95e5e708b97d8332cdd7b33f90a72a47cefbc09b017f57e0d71e5d061544bed8ec77124869909f7053aca728261dd4f4ea40a0a0a74d2b6348dbe77c1ee72c1f24e2f426e74c589eea4b1c10a7286f9f8b70b2fbd0e02cde5360dc390e7485e0a85919505c28eef0bbec3548f52b40e29d76cfb6c0f3fab4de2dc30960856add9cdfc1553b6fbb1b68209bd0549bd3ede9bf2448d3d98a5f297f357e69ea5b26d4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h18e4979620f1b9cba3d6a74fc17327d07b2ef4263e31ca8045a0c2abb49063e782752ef4f444468584983d08d9f16360b19ed5214cf07a619b6621277c04dc321df1a3725b05fc2d60d90eda2e3a102023a8c957a5bb7bb609413e4ec730190fa5116be548101a5511cf6432ae7e4ee2141622b2d66831888d1b54b595e288f150f030f9251c2b66ca83e43eb96fc1569d8145637a53ba15c78ef513fa9292d6c108cd07980e4961290bf50609d092e8f734f7e2100e4bf5455ad7f38c107de6a2a3849c6bc9369b95b467f3e8f2fdcb59f0687c9f3234abbf1d731b309dba4791414a1f558bb726abf4dd152ddbaba314f87a4ec37e41bbd406cc673d053ac0db79985f25d64aa639b96fe16f660fe0059b72fb025eb03dc686099d34d27c5a689c6f34d5e9439a83cd98878fdc82c1ddc880278217be1d8966e3ae12407d68192e0e6d3bd717d421f03ab0b5ce0b26496e8fb57ec523e466aea9c5a1f8de2a841967062679e61b12bd85d65444947f8e108cd68f92e0caae8f533c50ef52660d3d1d5b2b74e754d4b4fb1b155ac0f553b89fa47517c454ecaa19608f17d70a6513353af9f1c290c1673987e13a674c49f757d70b8d25657153c444cb82ff1928bd1b829c14d6d5c48ed8dae1fc336911ca48548df9f45835d669d50368ef3caea72e43a4e57c82935adcb5bea0fde1c7050f9a46cb8b54c9e3df156913017f6dbbcac71bd772ca64e63fef10e123c0f7b99888f1c9885611f7e2d00ef0d0089d3c19c89e12b3e4711f9d1c13a87ea3c69bb8c3e651818b3d3cf77d1574c24925469f43709a0bb2ff9ce5292266334dfd40b1f9271421d1bf8dc0732b0aa59ea01e29fb3a4583723216355bf0b48d0947bf54003d842e981b43048b40fc9bee89b461f8c8601324b6c2f94436f6b8af3e2f5d3ffa0b76a67bd4d01c86effe1c08b23521dff85115d09c06e04a64f08eecf6e6b2a64a07bef33b4ca61102b9852bdf0c8e11dc64e0c5d26d856132263d707d61b4dd2492c141f9dc1d57a3b9fe48b08a601ca5d7260830fc707223343ea59ae28b0011fdcc2ca078273c5592de7aed1a7dedd497daf7fb5dfc6960ea271b5e9f2ee1566222042d700f12563b77a592342a24d3ff94763cd1d2d97bb78286c41ef7ebaa5551f8e42e72683f5e63160142757c3875c039ade0dbe81e131dfc372244a70095a4d304f3064494ffd83d92175ad2ec09e56ca9c1b9391dce616db965c13a9ec851a6ee170f1af0b74814e8920686b73fbc4424a77e24d68d722cd08e8d3d42fc7dcbfb1ef04c5fa6fd2b5290eee1c02ba488470765055ec1a3fb8422a71bee2cc8128d665313b4bf6cee5b89df251634da90256888e175b8a62a9a4c4ad5b7ba556a4720620129693d1e1cbbbec9e9d2dda683b525d3844240194f1f733df98753e48601f92344552ee1e9e50c00526f4caf44c1538727ed0dcab984bf03f236ed83f97837cd2b92bf0d6c7d8cf47dfbecedf0638cc9e558ea0c04adcda3ae733d3182e2309e6ae53691ae7601d8cb6395e8b4d16bb591e1ff87d88946cfd01bd82d36715595912ed5c943554237f381a773d1287a5ea1fe43db45294b48172ad547b69d2125452c9d93fea62bd8bf0a6f168bd34949f3949088a315f6df59044bad63876a8e0fd8a543323c34bae278faa97c0384d71c33520048ad648bb11a51af191ed5afd7d9b5ddec12bd89b5a6b2d6a78727786dd2e924b20ab2de4323d070653c08b83e519dcbcb2b879213982bb839f23adca12a2e0a1c08c6bd485468bb4117f031801106ec7d7a89edc1a27f33a75a14bb325a0fba8a54d328ab0d1f7505ea7c1a347de01002389a97b257a3fe0e7869002944f809f041f71b66a5f2a469eb4a49ce545ef8788c3e4f532c157e8681d4c2b5b200f4d730d145134c5baccef6764041dd8f957fd4b7f7d5ef45745effbd4058e5b7ec27ab10394bfbbb8769d6c7040932e171c09ff9c0cc41539eb36cc533ffb1d09a203859eb42327901bfff25e63de98424ba64858551172019b122bcdcf88ea9fd3a04aec6f8cb8618fec436531a30f7b269598b652e85d93f11255f80a6996f8c17bc579acc9eaff7ae14c1a5073dd7e12ee0e3469fa143a346e5cf0ce2aa27ccf9e688a2c64fb18853cdd99b82a6affac9379dcf88b44991cf7d4b3915d0e8e089aad22c233b5e28a899d1e504c8ea82820dd0dc03a3322ef4295182d56aff74d8565f6b5fd0879a6427f1cdc241ac5eb5c371ee73eeedd5b5a168e75dcdc244c7facf6e06b35e9542657896afab3508622d27e052005b0ec87e61cb31a1ecf4c341dc4b15e8f567b7332b6fe92e12deb3ec22242a601047ae303088e36eb77a7db12f99357a411fab52d37d10ddea718a7775ce62b5337d0824f159411b753ce5c59f01ba5e9ad41d062ebefc4d0c88725736c682f493d90403cb6f81a61ba7839e79fe29130fb06ad63ca10e15e2dd712c1925059f8d0ed4cfd14a7401f71fe65514c8ea4c4c4d3ad1574c27e470ec3f030fc5a3fab7e3a7b69326bac39285e3c6622afed9a6f5cc1409d97452993610bccf00bc723206657a86b26e194fa3a944294a29c50c1c13b5e6b108008f6ffd26d6554ccf514163b850b4d2a4b792899559169bae5d417cf43c4e44f8c8b859ec0bf0fd32b2c35989733d7dcfb44da440f76240794407fc72da1aa40d87e3f065562d6ce938ded30ce7ebe1054dd26c84c8751d886de549a0c2117014972593d704e5925ff9f207c3bc79aaa6b2474470d60cc5e7da00bb5c9217f00960e4339c99f285ee3425553f9991aecb3e8981e6d625a11280cc9fd20751eb97f24bf54ffb6603fcf4acf2d95975ee1e7ecf02e923ea7ca09176e0ccbedba91aaf87692bb2a59095ccec46f62abe665cd16a18227d5d2f8f3d7d26c2b788bbead532bb49d9c99fcc5d2c1e48b79141ddcd41420b9a9d9ed4472621f2042e9a685126002ed622359b6fed7df975ba46dcce60dc39ff6aa185a9124bccd7292f4958e5ecaa413bedf7c7d70b7409aa93a05c6a9a5cb9ecc09f0e33dcf8da9d848e00d52e311fabbfd4b1864ab27bc4fd8066701c32f458370df8deac459590c648504315be56a5917035741fd987ab3232731322da723fb291f8f31c3f3e6c7069c2211d2463534b821137c04d75b6a1c03584b7d2ab7ed2bf2b054483df7a7618a008077029689d8c1f5c579f2833ccea7bd4c8dacebdc2b456c266820243623f1cc56173c95a08ea4bfd4c9c7546be51f9e5d8bd320c9f68dd0b3b1ecad15ae4d7e86c58ddcddad7ca0635aa2c674d8bdf62f4f3ab9553e3cbdaaa896748b2c18ac25647740d4a3135f54bd3f552d47337feec7e1d348571f484f48cea8b56f77df5e992992892b9be47f49da7cd6bb9830f0fae1a5812cdca36125c9f0a96fa981add96d91dfcc52ba9c098e8fe86d30ab0688a9d643f753ac4a255b06a0e7f62965a3668a3a8146706a04c8a78fa56c6f5bf4c5cc95b44571c3c98f988cb82f12a782883a6dec399ca95a43398741b133c77e0e3ab13396bf90cdaac8b8fa6d9deb62a88c8a3a401c8c0b5e8edc6fdff5aa0d393a050bdd69ee2e94effac078042fc2b2d1adde51f47168afe2b9af2617e0cc0d31f3ee4ae731136485af91d2cf7c98d825811ae5d09c3fba85a3fc90c7ae4afe30cfb7afa128601364c0f4201e8f8414db04de68c03becc74eae02cc65cda9289a524ae4ff5e3567ce53aa77063fc5231f96de5fe267b5f15592e044d5fbfd7c4a3210cccbdca87a8856da897f1eb6cc8ff1d3b319ac4557ca976f0bed7062c2b0eb8c2b3c320bc07ddd598bc6640dbbeca38f7edbf958dc4106609615396209693758c10fa94f162c30fea0a0d1262dfdc8281045ce5ec2f16e72f4e99282ffd7be2b8042b8c8a890c3266005fa651579c256f9bb64fa4d9a34d506b812e6fe422beaa7e2b6a8d25ab8373c904440f6f961ee09f0a124e0c408dacdb46df1865e0ae60a9b4557ac62e32bf80bfaf2463af591cd144252b144d11472c80d39dc568bd490fb437cfdf465bf4aad5e5e289381a7c1314d0fa08ecab78644e81d3372cb02a26b983e9ab8cff19349eb5ba63bbf30a16be0624b728076d9db1eda5b6d602c8313444228844013700c6549aee7d0d948fc3142c70227c517f5ed1f3babf73537d6cc32a3a29a642ec58645ccfb028bd9ff20145bae6109a753288d57ccb9783ff5652e73055592dc86b80253cd4f292c2f1af3f0ffdf03ca6b4cef6bf1f81ffd39da7a9a107dd1f562275d71c97db53a28ccd13b3242703202d9cf868d0f73eeff621ed96edb435c5b1ee9c650bd21550709ec3db40519f6a5eee2dd06c87b6dabdeaa97ffaec6fef37e86cd1dc5d33b840e1a7f9d57f1e1f6ce89817e024a0fa1b1ca987d41b37f78818ee0cf5f55639b25408475ef9ca0152268e21d797b840846a739f6c282284b366f55ce992bbd86918442a039f8dc082cf25d2f09e8c8740f9e0ada139a4966dabe4b8c2249147945800253d15582f29a84f17f0989f6d8b57c05faaa937e0f33b060883e503f30f68773a4be40ce094322b80ef23fd70e27433ae0e805ab3677be772e4b64b31ef1650db37e90b47377f6c0c8a82856c1828dfa8a19f80a2a94a505ef376531dae7d3ff4cc139a7cd33010ee4872a3ff90f34662eec8a6bd611612f84199250c2ee59540731eb5969d47c892b4cc04a436db3216e7cc7fda15e2e91e49333a07a4d096cb80c8820cdb3539211271054aaa84df3cd057ed06f5f027f8fcce9f6ee69dda5c0f025b2917f6e3b0ceff7f0bba06a1f97953ab88d0d33a09f9584a202ca8fd87a8f640aaf88b6905fbf1bd99b0d561b5c12c8ddf449c0a7d88f0f5dba12a797ae14952b9b9ef76228ef952d0574405e73ab42509d7d08995d4947d15e2e4b330b56f60548472ea010c5b8de1960640d9bf44cac5550043c4433d248c7888e40bd7e9a2cf23d44a85f1a210c0a6505c85a6b04da1afa0f792b836ae28c5b195a09bc932d35d2a4b5e951d7e5f611b9007551cb7abd01587a6ec4570ccd1b6541b235a66a63430cd580563570107e722d0b55b156b0a0d7461d27fe91ecf3e2b943e26333768c0c7c17adb7decbc52ee68a95d51eec93363a81f27e0e0d9a892cf7ec5407a28ee0d6ed753fa5690a6a497fd3374861b181557d60bfbf539240ee9737180dec7f865a9340a52f3bc8d46e4d72ae0eb3875d7b2531127c971ca261cbe51c49df155482049cd09a88575e7fc52ca593a868407d21f6b9e5c1ce21d7d0da6063acb51c51b8650b67b60a86d276808d38fce64c7f3799fefe567e46d034a6b4d283cb89d71a9e67db269ff0c249e63ad400f852b8ada901c4b8ab0273bb1f09f57b03db9117f65c66d9a048350288defcb56a82d37fb75ca9b4d97d3301229292b53799aa3ef8d378bfddd75a15e2259485ff54676e3e320728981f507c7d4745c40da65545765b1624d4b73d84b23cef7dc4dfd5b2b1d3b73bc67c64fba1681b767a22636ead8ff5a357e508ab5ee92a775baa638703b1390affe7d4bced4c2ab89620378bc07a55c02a10784f71f68730bc1889882d5a5bb98c77d81e82b366cc8d0664be49edf5430bbf537254a5cb065b89a95200b96b149268152848312a44aeaf5f4a8a6689af7c1684def5c134dfdfc552713af84e28a9fe7cde2eb47199769a91811272824dfa1477b363f2d0d9d6a0f4bf0619fd1cc2c43e196495847e3a321727ef0e823a272c99a49f113d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbd5b86ee43a57d15e7feb3ce7297936608dd3ccb3c73999b4442bd652366f27e70fe60df563abb376bcff8841e9c12497138a62f8a6dacb0a4dbac69bcbacea748c999b853862c998bd33f9477195bd7dea4d656146c71a27ae2872037056f09967763aba140a33f017946a57a9342d71121a7ef6a6dca027983ada30352e3d102c417d990b59ecc4db0e23323a9399b51a67ee0c76bd0ee2cf6c88d86b4f5e894c1fd05e84e49cc0b0e4a1cb3c0dd03dfb3ce9ebd8ba9cb650b34040e7acc809e71e18ca9da99361d3ac5f2dbfeeafc4442eb24018784d6c2453ebb2cb95cf919badfc534d2db012ea6f03234d919c6597de1768a6e8118a1e36a491717bb19b2649ddecc2db3e1f278c0006e887ebd1c1d9b9d4ef33827c9a37a724c795a15401368935e5a5d159f119519ea3aaf060a98fd0eed6999f0f1a6078060be963129a3c46b3658309f1c8cc2c7ade697972e7ca0088985a6a92c5497f3408d12153fc386005ebb1292b5203ee7cec5d2c05963f2fad8e620d53bfd676c5b9343f7dfbee69005a0aa5e4f36ea6b2e5e1c1f172e85648740e78162b3cca86e0ad11ec05d6d559251a18b31cbcc8174564af4ef6260140fc48da4dc26e2a21721fb31db062787c8fbda8e0d140d96748d9f346f10161e00bd22415f89e01cd9c523911ea0acbac17039cea2574de0b729fe5f8421190b770721942aaafafc42f62e52b9845c41d666ca15fa668fd096fe67cb8e22580dec88a88a3721e3e6277b50b4e51f28a23e69772b3a680d62d28ac1aa0d9c92822a4bfc5ec53df574467f2d13197825dbf31b8d2c103086f108cf8ef45e9bb029e49094859338dfcf4a83fbd3378b6246669f1c040f4dd722358e877aeaf1d9aeb57c0a49794e34bfd3edf3fd83a685dd641c6d147d8a12f7ee0c906a824b99d63cfffaffd7d883291721faf8b5d8b74c5c08577ed02088e7b739eb4da7940855617b99eb033f4a08b484de849d8a4af91d3b9c35c038135c0609f3e326fc51dfd762c68978b987fb44aeb167334d823488b12cca395213aa822fb460e9a0df5be739501d776f5203f80dbf38633da03a10e16e546a70559254b29292b1b1546c4d0cfc46e8d903c741f9ca4e1e5751a0b4b64a46824a922ad6ce0ea627054e4aa4f69c74c554540f7ba075378910cdb4931a5911e2a0e05060679c8a412290724b59b90ac95ad462432167ec6fdb3518e9ae8308a3bc4ec21b6cf0c3531774dad00773e9c44b509d9333083fcd661fa44a7fd526f61cb4fef012d2f4e954169ce9d1fb315b254410caeb6650efc39fa18879b93c476af1572ee3cc7dc3a1e3e434fdbfed6cf2ed181d43b7d456811cfcf1db1ddc922f065cac0f7901807497b9e20156a589be4429a3914047303e632d4baaaea657403b1fea253e4305a7ffb0a4f7823470e6cd6a5b3f6c4d27dacf7e2342b0c74972d300c016c741ee5d3b23b78619a38d305943774fe2fd1740e54372a0c88d52052801e1cd3e09a48325f88898e620db49a322ec7bf3c8861e9bb8c0f54fbe5c80ec57b11f77635314a72f8b4f8467f9337b9fdb46fecc7a706fe06d0fcd034444ea9a883b1f18e7e324ee297462cc90db81e6b01c506a17b789804ff15c306af104542c3b03e1252170c7cae62d669f3d4bd9495ff64e5c2a158007d3d7bdc9ceca3a1305c4a146079b4c2d1e89bc9c34458e663ac5826baff26d00ebd051719f0126e0456431ec89d0621c023f2f6f9bbcbfc95cb471ac74b3cd5c30dbd401f6c7549685ba6012bfed3e36a4d4a12152f06e5e30e605af85d0d06db0ecc283774d8e11f5000ed1ea4f05c80bd09656e74d8c1b0915102da1316b0e0c21f427f6421df675f7bfb532035192e53e3f6948f26398a403164baafbacd02403ec1a62bd5679885a3dad8f4992c68a32d93f1ae1e680ba8e3d74ff79d77e47f97c0517406d5232599126b169550295e2b96c60b68ce378125dfc9771e5762d7653a77f6287597d38c8f345403eece9d04dc98ec1a5f52bee0c8069179bd8aa1b1cbc65973900f85694844b67e1db28845743409f7e88768b937b8c8f129f66cfc9a7804eed6ac5b93a6cee2f7a777a99fdb6813e194127a98a51a78a6a301a5864bb1a8326c7f8c258ce2902f6d24909c8159bef6774811c5c12407c63e7198e26382983ec3e02264525667f7b649b7bcebddc71572769571f4a9d435ab46e777208acaac3981bfcba7d9f5e83a71be3ee1ee3b7de723f8a3751eeb54f2be14e4ba0edc7f2099fb46ca62241683398037ef881c4128526aad1860dc09e6168ac0830028dcf2fe43cda0b795a7d33e15587f6b2a54d640bba697d0dd64617126772d845bdc0e62695c0df73bfb94f41cffff4e51e9a81207fc93ebfbd6c706a56dc4505781720895912a2ce953dc5120e74029802fcf97e5a572f87c510716f050c05798b95d51096f3c4e9312fb7a9c78c74945162d2f5d3a1b596332133f156099e7d39e643848616ce3e6e784e822217c1e983eae34be8758db5cf105cf68f07cec6f0e1c7353f04f3345826277f73ee36f7832ae472a8419d36a28c3b5b896301c3f1ccbe72b3c788bf386f8e4d0126432a1ccc0d8a31f73b4e7ebf03546f6520b5ee455a6fd4f4c18581622fd90c613d1bba7c51938cba0ad3066541d52aca00d361371b75c88160370b402aec996cd0dfa397bdaeaccf851632548e57c22d4e7a97b10cc84e4c682c7ace8b8fb6b7f84ed4c894e103960a78a8ceef0b276b44be41ce560abcb4b7af5baf29ed092bfa78ca221fc06135b092c42f797de5cb7abf0fcc29e2a22baab367d0e71ab9182eba94f3a103a98f434d38e6f9d4c3301414d24795a5030b114f3a771cddaff7787a3a1f3ea359f0f024f0d30762cc7e1d286a8960469e283f37299c098ae86e2946ae23aabb9820f48ba7c2d443973a737a5eaee430cdcf1198d8d0defb99f0a07f51a2483ca8a361d28e01ff04676df3d9db20aa1a2a1c73c71667d264c27aff757f590f50e08db9a3c1ceee20ecb36d2f27263b7f7abee45e001f52ef12c7146809ac1c6efa55b06e82183dec0e2810416852f10987653bc14fa5ec4aadc8c5f3010612e1f86d5090684e374eafffce7b4fba3a6736bc159ec232a3ceb5729c15210f7fd66d812019edb597e8ef1bb779bc0ec341f201177321e24fc20740e35f620a00a119ad59bf4e3e721c283e1bea75841da9c905c2a7e3ff6d781894d0905ba2dff669fc2d59bbf317e9c0e52425eb6e8730677cd20d2be29bd708b09853b7ff1534e5446fb9dea75288bdc11c7f39251dd99d8eb3b434d036ca7295a5175357bd7d17b312645e7d544dbac8d6fcf38cfd75f56f1a0ef574d77b5c63a08c2c383cf37d0357e7fbffd813465ad485a20493c1e84ecde57e4b52c4c2089ad37161fcbdb107adaff780ee755f14c9fdd25c15d606ab5756e151c13136ebd2351c9c5aa6d1208232c2d9ec53b2c1cc9b83688dc693d0717f96dca3f8325a21529d3c916d81593c955fddb54ecbbbc42f913fad0eed6f7c52a8b8ca37ecb153e1693e6d3caf97bc658660ac03c8598ba32f7c55766116d4a8ab56a0b510465182abcf13c13f61415ab4fd0b44255b31ec9fd57380354bd77a196988b4b9850a5c19181a0f18e99df87e12028c4ad53f485681ccad2061ccea8e997075b827561beba6077e8a942361ad729212542c532cf837f745359f008420eeaacf770b2c64f88013741050e9cb24ee27522a75bb430644bda0eca127eb81c575db9aef75fbffbf6c6e726012c2afe48192e0741e6c87a96843b4516be2d97d4b3cab08f2c33c8920abf8d1caa1076f1e5c4811fa257cc9576420c3d77fe391725b1d7f751a0ebced74831e025e704ebfcd28712851f294bd36ddca6ab5ba1de137d76ab54d0d56bd684ea7bea5e535d82c74471ba763ffbb93aabf25c0b52802b955aa508de91ccc1fb441cecc35323040df143e380b6142f47adf7eaa3f1bfd61c6b6e22d29342c489670100697c92c8bbded8db0dafafe8bdd66636f9a615da4f181035f53c5a59f8bfeda095f91b638296bfc0dfa6ae583e61bc9b59848253e75ba9da55d91feb2127fc8a566ac946a03624abede1cde9dda52477a4cf8b39cc1685a402f7f1b8435d3aa69ff18f783ed227fd8741975a913f8ab654647b41e9ca0c3ec516b7a283a87899b782289eaa63ac3664d5a3515cbd70580f5cbc9518f4859e4ce17d5c3dc8ca8d5cff31d40892ccd34813af2f12e3ab28caee27eece29893b4cf6a8f4466ce41954df2bad6ceed5c01235f568dede7cc91274df20ccf545a99c3b743d279fb199645a187def6cac5d77589afc73cfb16bba3f909a3bf2fc143c965d4566c02666148b43bf7f6abc7f18adf3d38c20074acc36025a73b71bd6f3988f39d54054293c6d575ca3a881deec67b60f1d6bf0c2df27184ec2944c8f5269e9b8425eda6d5d196fc27f215e1b7d7b4329809244e3d309e731f13bd3fda5faff39c78d4eecdc785226a9b0eba658ead3db9501f3d3500c617e33e6464aa59ad6e63a8107d14724e96e2ad3b6b976be2b2f99b1df35baf7a62c028ed07299d0df989cc887dc952e19904c2100d07d2fac8d67cb63b2077446b232c34b6cb29ff1bdfeaee9261f052681eea855bb5cc603e144b0243de5f873d8e7ef8f693ef0ddd210f5453274e5ef06cc3276e5039aeabc8c6be28109aa6c814699472b374840343e9e2a54570f825263cfcf0023f10b66297fb3f95494e083ca37699fab9aa3d967b0dfa524923331cc1c569df5a2b68ce9289867d4b84fce5fde1b780565fbf4c55c7ac6828cd9ff4f81f55e6a26dbd4c96f3f5de611885bae155afe46ea0fa1f1b60fcc654f15f2f7e58acb6becf034347b61dd4229d25e9aa9ba233f85e56b92dd39c689b0be18639c3eeab777ead5d4bbe56ef7d8b4d8c19b53923da939b77c3b045df725218b2a43ced8d784e7ab52b0bc0eb1e1e84404e5c4149044dacb3faf4ef48fd8223b4a7ccc159175b937a696534bcdcb4ccabec709f19a52d41a45cb1cb854f8de9c8e420f0742e7d3b39a81694665a89fb1abef9c9c9b45e6b07cd6fdc56e44f49bc7f7894a7e795358ed1ff5b5b95c1a1408abc07d1eb3ae8f27e15e960f0623f83062803b4234559b5016fb2019dfe16b5a1d5b9e38baaa87a6c9f88184c7958fc393152193e3cc7c6b0336c25db873b79b212771fd3e12847c2a85622bae00322161ee074a1d428d9e0175a9bb0b41944849596099a9521e3e01a8ea9180a4f54236cf349e93c2f687964f4993b2349366a8c0ade11b310bdf5911c591161e570a4dc76a4fc3a66aadf6cefda9f981c48093345355fb2228e2eefbc43c75458b55bef5889a67247e723b9b5ea0103356098f843e671341f9320583297138186dc66d9c7f88efa48cbf7c9ae64b74c2a66c5b8c2ce007a7b1f48c9ea9d0943946b214c8c4d1e368b41c4b26b4486a3fbece4ed65fb68b67ef91ccc720fafe2b90f1eebb0c2495a3012b45a299a6c1a8c3bd4d6f266fdf3ffc99c000186e1f6fb6e50c628b6eb5d2b966d5ada251ffacb5de0afb30ba92a3bc799649d52731b2c45c5e35f50abe7acc7be5fa02d3e52fe71f8c0ec95e77b105098efe0ee5a1a89000d73f206e4f5f70d13ea592de4293595987597b05f41f7d0622f6f799e84bc469b01bd7efcf7ccc818f6ec786077342cb0f2700fca15ad2cd2e0709a3460c8851e389f310bf6b2246456655dfc76a3a76c67b4afaba159b8c05e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he3f3ed3c11fc58b584bc547ff31bbb27605226fad699a4b24b14bd4b6c38f9f8e55b591368bd9972eb42b92e94553be62bb6b33dd9a0fb2fd05613b3fb29ca0dc6d7eeeea888fc809927407a61d56785089c1f68c21dbd97d9dd3e9b97a705bb2a8fc19d6d8e860a6bd7fe76bc65c95a08e0c0edbbd95aac92570a99a6103e7c48991af55beb947e2e991ad18e967b9c4e7a6b214895f2292de08a741d57759ccf07d46d35d46c5815b3f6fe503bc28021e39c7fcc49902c15029984e250b87503b30da4f583c2e1dab1e85a7dab55e890daa656ba6a88b54a8289aa9308a58dc219a7ec7ce744757ae090793fa1e32cf2dec32ae1feec95355c4dfa0da40a5eb89fcc36ff97fb0008d061f6767dcfdece745c5c5735b8c731d3270db7bb165e23c02108d13f71f9847d0e694bd7c365a83465a609318f0db1bc5e761ca25aedc0591e253eaedd38d16ee49bb779deac8c5b2785535b2b864a96dd641faadf257764002f08060a2d2e8cfc15f812f3a1ffe28f753052d92162082251bf6e92eb9012500c2865330f60ec0fe1d0ad61ccc2422b0521d40fcdf835e2e228e1f5bea2529e87cd781d27d94850686fd43bd5654885562ee7bb61a501200a230029c80ccbc4df02ff7483f2bf0bca7a76c22f31649b8e667234b6081058c1e926dd9f5ad18ea011d9cbe655fe7066fbb9dd9787a7b0f9f5a82dcd42251dfb4fc89a728b200c14a015ac8aabbeec0e1e26942e9d7ba78a6da2ce1f5dd891c22ef60e43915362398f5101d532c216a69753169d16d9138901b5ac5e5bd0bda834fd60bbcb77c7e0f2de787cd9bbc32b51de54923536348e649aad32c05fca5de9a6fe287f778bcc349864f4b80424c74ba1c372e122bbbff6fc55da3a357d7498b530c738ec498df7dc15a0cdb1f8baab295a7eeb496fd505e1335b556cecaa2a3598d093655a91a06a952c486ff0a7ab910c80152d83d865d9bb8738f0d14bba03d675341e0b5366430e4f327ba0e10ca6b69a95311bb46bd35c19f96965ea448217ee235999a344e5e714bf9f1919aa56517a6c59eeb4c49abdbf16f0407751d71a75f3de6dd9e3d7269269c839fa58b3f3742dcd881b7fc693aff07e64e12c9eb2622f3a5811a4f51dc3c4ba2d3ea0ab3b03d1338654a557fafd686676a48c165a6bf81f9fd30257ec28f067b2c03fae1e6e6a38bc9eaf633045615a72452df5b81d0f8d3111eed05f6ccadcbaf7ffd08256387a00299a41e137a606abde4b62c3ee7e56b66bfb830cc8b0fe20051946c4e3c6fa510f77bedce28361897be8aa10e109b6275cdc4a39a8741c24ecd05f03eeab888348cc97d6d64d6c322046de6ef1404a962e1c4e49aaaf7573131235d850bd5c99d4f2c8eeb7ba1aff3b1e4b9cb8e4a7574500b4be2134005a019794ae1f0186b0c3ffee864091f6e443353923ba2d506221de33a8056efcf7cf163c705118b3ee9f7bd653b312fb25a83a6ce00cdf9ed6d3a160f84d323db83867d714459cde62689080182133c49336c888544f6345a1ad772af2088dc5de5e926f2a67332ea55fc997f3dc3af41b0e8643c8aa3b599fd10b1c8daecfd51747c0b182c4bb4a647c19b434aae7f07a27e95cb3b92f4f887717999d2a86b08acac72f5ccc48e85c91b60e97b1efa70e84a952d8920486241257d05970bbb54b375243f68f19e70d637818ee851661b4e9cdc80c563fc5d333515523ff1c413033af13bd5685fe5d9315ce3c3678723ab81f1428d6b08c562e750b68566de422f0a1c7c5bebaa430fbc8673e241551c1160c8b891096f3ad24707f494644606778cdcb099f6a7f572abbcb97f366e7162217e474c4095abf90ec31d254ca66965d8a59907ae9daaaebdd492b4e03d8cdf1ddb80db831444d1c48796ad4f04d4938d4e18d376a59341ab2f363898dfd04909801ed78689bed403bf5db82ab6da8b5c48158c23204f4a00dd26b181a392aadb06b8ee4edae0a09db02b51d44a84f80a9c3fdf6f222a140743dbfd04e204eb8280d4a6ac330ce8261138efdff27d55f886827e8368c43e6fbf5da115deda01124101dce7c92f424494c588bd827bc3c9c1e18a90f33411c3700ba16b3b59bc00cb33a6ca6a1cd8181fd51c495239e15d6c9980f21cd539c218d6f31c4e30de68a0dbb91b66dbc8e1839811acbfe00e4d2fb1f3d173c2079fd82a492d1e1a9b58da912a7953884a583dc8e88398a81d4eeeba67b352fc91d770021b0b2cbf4955c27757a7918f115f22a901040310ff10a20e64c2971c226d161334c9bdc14daed75d387fa79fc92b56a343f2b8490676f0d4405d29c7d50861f85e830573309fcac90ac8bb378497a7bf370d306c98c63d593352da2ff4344fd53a83625a2c614fc3002b527a90f3c02a9e130ff7675d5a9a34443f50992813ab6cac93cc0acf56e3e53302c817a48423823489ecc7a5910f0c13c58781b14d26df399b8299739125e1661e1f8e6c719aa7ac8eac225bba2c501b3577fdaabf5e6a7bd7eafb19227e07ee2dda6697c7318d16b39e3496481f733d7f1656eea7503c254591f81ef0731e55075e7fc5f490d652e6cc81668baaa4456d296cf70f9f4da856bf16e29524bd689097586bc500f9ac7a5aef10797fa0c748e04f96591cd2956473137fc534edb30de936c0ac3b3bad23de0aa15331780b2b8b0c2af59732408ffc7e11ded838358ef3254e3e69f96a1f8cb1550463f912584fdbb91f1c0bf8010cc981eb6335dd625ba5eff2e4219a0d37303308d059c1bc7ba2c9b230365e83385f9d05aca9840e89d6365166f2bbcecd4f14e642acef53339f26c118e9ac3d1ccbdf8dc7383137f70f8b53d9f2b86f4bc1dc2b6ff36f12b6b6d9608869a8b6d0b555df19f640ecbb3f91f39aeb1676c869f6ec265d1c1b0e7603d5d032515d5ff600cf32cade217857c353efd35c424c3967ad22fe06b177d0aa3c216e7f4c1101ff0707a4b2dc1de2075ef97ad072ffad268f467e33fc4d8b9aae35b4330cfc19ead2874103b8132c7a1a7e13ac480c08953ec39929eaebf622ffda64dee7bbc0abf5bc2a1bde536eba1f95b0bd378b4655057e4837a559972bfea25234cfaca9001645108f9d714edaa43439b02303d16e13aa92f5df75de794d25da9561a969d640db9b32779f3f4ca00c94978f34728248ef1e702bb3b6c6dc632deddeeacd38043f6e44a0fa0243d5a33516382d7a7e1b3a05178c1d96fdb3d4b8571ea083d09bfac93b293a019547d2e5c4d626037862ee0663b9886bad9d5e4eb76fd1dadbf99d8e8ebe663d1a5e5fc2743f55c96c12ca1a3d267aee1cc487dbe2c50fa293e745ec01511becad823472c1aa216771289c6992d77f4abcbef834e9af3a94f07137d00e266e912760b7b3b2ba48b2e52e377e22f9c428baedf62c698eb130354a77b3505fd7f0dc138933df1f7ffdbb64dee8ea3283293a06f64e76f6dc5724a48552cefc3a6301035bdec3d7ced44f9237a5b43363989eac7ef80cbc49aaeeb8b05155f51f7b016edb4804f820d644b649b12414cba8b0a9d70cfcad51d8fb6a759c2ae7f6ee320124d1ecf1ac4d6b37050e37c0a72f4ffce764c6001c99360969d29cdbf313e4bf9489256778086602bf5c0cfbeee856ba797a8b30f727691c106ebd5ea25ec3d2a8d3a3869d87216577c56593fe483848e20bbc1e54f6966a26a3363b51c907bed740be8d30079fe253bd9a54a13a3cb6b6a7affdfc90b557aba755b854f978646ce250e853b20c21eddc1e5fd2ce8ff32dbc007e75376c5b88687fade039d5fc6e26fdd6a38b9890caef71bb9232cdcaafcec3e533d6e6476d098f9ff9ca87dcf65fe7e09da3d661565f12768ed463efc3d6ef07eca2fd2c05b8fe6a1673407fd421fb93aab841d7cddc3e24cf273edee8d008346f6846d628c04550f4308cb1ffcacb5cc8db17c46f58ef02a9c0c4154a8b26de42c34e8356a4f914b832d27b1dbe6660164ad6f09af50a8c11a99e4cb1d98c9efb276fc5c0576fc4e696efb69c24d7cf30ce172cb31df582de7426c332d8a7c5dd936b436d1c71d65ae0c9e4242b47098d0dee160450842847dcf95491eae5f4ce3d67a6b0f779f86d9bb1c87b2ffb158368a3097930006b7f3870a80612178eb76eecd854db62b0c0f22b8e88e1b3abb21954000825ea828b500a526ef2e6fae689be7c3281c78f923ce582b9e72ccec941d9201ca4fb4ec2fb19a85107e878ba5b65bb9bedbde4ba50fbd8bbe8c8b6ccfe6ee618363117f883e02fdcab686db97e7304ff3bfd09eacaf62f27cda52ebbf7d44f506c49cc81a54c9ae1270d1e6a90828a6ef1cbf00b8f657b483cbbfff08eef7883fe475ea04008f7226ace095bd8fab40f1097546c02b5c765cb432b196244d692402bee4cecb7056ff5d27955295bdda469d4fa30a397381ffbbb9690da8a4fa2a2bfa18b205548d53ad37533e907746b0d0115df5052d601d52efb467f958313f4df763670e2d08859854aab029ba0d7b2282f1be77218bb5b4e518cf69c768dc8da326231891c6f05a644569813bc8c387f26efa3ceb910ec6b484d7c7d22a2141851bb53e9610b75cde0f1898deae0be5179799fc1e733db1160961bf2997b74e38ce0603c1a434c5d8ea5837fc14a6f4eaf4701e67a6ff531fb66debf72c2cf817c9825327020e5dc0e7cd5f272d35fb85b8c59cef11edf8746459e13f94c2f360000e155479dd4026a074d718764c382d0f547fca18a0b2b5641f40bf4c194089b4691ef0fda59a6f067ba33076ea4613da7b82c615d95c53bf25a5f81afa2c340de3c8a8963f9f2658fa889574b779331235d47f5536cb2e66ee100bd9faa6de8fe04c6e4f0aeb802ed9253eb9c6172ab124f836e874af7dbc778a8de086720fc1a0dee9a7ab95f13629d2134c5d12e8781ede9a244aee3bc2b23902ec328e1907ede9a63355bc8dbec0c3f6fcc9d4177b63ea7c3f5e7a37fc1ee9f62a259e5a90e19528be7326c8ec9ae950d9ce201cd17536cfc46857c97997d4835e6566921a7d2521ee913ad1f84f2392cd8f64ab0f843b4b18f225978df189bf66a40bceabc29617927ad8570466748296051c4c21e9155d16d1832e4c3c4caf927f1a6954f4df9eb352e44d2a941e3a18d71f6bb1267ff24801a99c4478268a58dae208f846a8fd5245e83c30d63f2199a0bb1987f8e48132de5761f6d50e38513e9da31430e2f6be69e1f0070dfaaff812d597e6652e2dfb3d5c647614e29629b374fa8856e7991d8ea9e4945d42fc94f16c54f39786760eed67fe863017d4a811f270397f43984098ec92dd5bb63e76f500e7ec4594e30b9b22e2c13db78332f9041a425b30dd7c6a7f006eba555f666d9704ef843eede15a4ba8743af3cce5997055e08886e8da9d2b8a53440395795fcdb7c8a3e2ece561a33c1b085bea19b276227802a91202dbd11d3bd7a2fd5d59733a380a4ffed5e1fd55c5aca9445986bf5580eed1a23b05dc4124c1f944fffb21c513445511ef2c1340ce4c087df36b62035584bafd85453c705165036f5e661a662c41096a020b665bcbb46c2f0f4e61649ec5620460a4163df096d79ad8cfc05aba356073a0eb695a37afb686644db1c4c347187f3d2c66f68d4fad21b49698e8c77b0dc3729f164005a109d9222eae74b00fed1c98726f0bb4070412fbcb3c29ebf961618486afe6b09a6a9ec4eb20a4c417d427370a861ff972529b5f152740b8c64b96aff0373e34feb18da9f528e7e791d1e2c7911b371be4baa2271e2b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcfb7c0d3de97c82d8a7e772803bbac1f1b246840b96574f67e7f3351a75c32b5dbf62cd3a6f26400823725b3d9eae37d06dda8dd886b923d41682a6e067422576541775a691082151e1ed7a2793657142cbf830400c3da1f3a67f4a808596d4fbd4be275be2571c905b1b7f4efc8b89f61923382b6c4419541ee2a0c94f64a34e340050e7b48e35de44290591380a1d28a7ee6826b190d2bbabddab64cea07e57d99af89ec6d4a1bf2ee09ac07329d7762a4041de737c543b9837fb5af8eb3a39d45779aac703fd4d6ad8629fc49efdf09cdf800b735cd120d4aacb90200bb9a3664ffaccbc51703ac6f4023cb2a7a9d574dc0da938fcea4c455bd6223be2ed88a4527e2aac05ee2c27c956e229d441a70545c72b1c27342fad7bca687e19757a11094159b2dbde07fd7e15aa53768c7f4bf70f7719088b0303c547d3244cea9c48e0542357b68fba155c8fd6a8b0c79fe945a7ad459433b313eb688c119fb9147df7c22fb8e5d281188b08be0e0071c6c6b37f4f8bbedb5ea699df3248ee809c0a20400e3033002fc88f02fff2d49abe2b2fe2758e2a4c190db1dbc1312c9a31f796a9c93af3623a54211b0760ed5a55e27e2ec714ee19bf4652a217e7f2c7fcac10a9b04075cb9aa19142934901e7937fd9affa9b9b2c620aa8f315643814965afa0f43583b86c4a0e1053c8e5e93211a55707994d45cce63a67376764e0c37128c72d68ee0c9d1ec8fcb5bc7dd1b8a0efe56ee628502eef7edddb959c705b6f70bb51a9c52fa18c28ec52c986430b7e3c7244d40242aa61db6d7b5373875ccc8b9decbd8e16735ddb05c71f71f17f49c90c064fec6740f09d0ef83ad1ce9ee092829b68565ffb113a2ee764c426f865327d0e85e4f0b719df766aedc8c84169d8a72b3e794a54b60bb96a3c97b41d8bb5db567a5975eeb9a364d6eb93d6dd6b93c9746318dab93d43fcba4290bf680f47e7c2d985f61dae43464518470a99dba44faafdd31503b16e757592abdeaaae15c8f9d13c6f1e108d79e74de5ea609c1caeadd7c9455f9b77dbbe47416e5dc91e7b5f8bc65ca57b6ff9062e99c7aebba7cc2edd88ee8ba6aa7b131804467cfdf01c802aa8d717a12f850b1241ef14799801dcd412172bb26c6c2cb59d96292532d3ab7d078d38847facc89901b55e7a0dd9d5f696df42b848fbc73395749d8dc9fd1810a10ee9b4eaa11afe978d175f49ae718398a98651d674fbebd8854f3856fc07ced7b6a4d25af6813982ab9af7a9624e60eb94f0fa059323a67b11245fe58541959136c6554a5ec8e4e5c3831afa728cdde3f6af23bbdcbcdd5ab57e2a90f4cf9d725c4fe314d00b28c9476a4bb52552f94c53daf87828566d5ef9201cf2bf208d5770fcfceaf81f76e2f38b5f894fa65fb87a73fb6ff0191ac2851dabf1baf26fc51d37ab59a465def93968bf4043a1e79544b4f2214aca7af043d65af7e163d7a552ffb6543b32d462f3e4d88bbfccea50d184d0773a107a4f3a6382995f1af8758dd8c55fd70d6b8083fed97f900507e009d940152ef57664b913d72bbaa51836d833ab9e745bf1f4d54db56351c0f76f86aef4918c78333449e742c814dc390904da26fae94062718edf7f187fd7efa3ffd96611065814624cc6a536f4f226f55177e52f13dfc339bc519615156947c1ffadb714b8467d6c23042dfdcfb2eb125a87b5a3f6e0149c0bbb12f68ddc6e5c97c9dba5e04d1e9d0c72f344fd90347a2295c2da3020d19ad6f3db36630e017b9228d0beeacc7bfd45105bfd28a3b52c359f084831fd4966cdb59863d2689a3b217bb544ff91d427fbd1f07fe7caeef6615350c915fce32294b2b7996660db20587cb099b3757bf7a37b140838c12e61d2b3e7efdaef94863deb5cda24e10cc06d5f2ec87ac9ae01d35bf2c97ac4deeee2afd1566c24b3f1035607a9c8ba53e8e5120e03bcbbb43fa2ac787d68b252caca60ab723c001d21b8ffad88dc494a1c7a9056e6ee486387585a57321f6eb228a9f7f171381f5a1c829267aee7537aad960414b4b173ee789fca6e9f5053662f2adbf8ceae6e9be0e720736692e64e12b67d2b1e51114bbb90c9cbe82c916d1ea23d557a522e26f5366e91af108ac9701e30b8d2faba7c95817be1171d4712905464ddcf41194cd4c754d4ee3046f79d44a8378b33432abdfe293c0f5f9af03b12255dd54aec9e5b807ffb27e4610cfdd95c1dd243c5e2e89ce3409f064cc51ef5f1a909c2eb659f784d41fe525dd786d926047a7461eaea8a5e4f4399902217388dca45eed24a35e5ad2961e93bbf361f85c01335216efe398c22d97414fbe68eb1d13e21e0200a63a3693249834250188f2b6344632ca8e38b0083b9b792ec38b1be2073cf948e63717ea4837742f8d9b8ac09f7deeede25ea1f0f5efdab0dc994d9c5eacbcc6e6cda0b815454cff5dbc514bb821f1a817b886302274f6b51f695a52c1546865e13fcab88634f7fbaf09c4389d80ea809c1c22d8353e4aa5d75cedf4396eb8938e4bfa937895e81050cbb979b0829c6045ab7ce885418967c62bd5c61a80dcb54c6e3e4231c5455db08d1f8a4623cd64701d3879cce8368586b7a81cd471980871aa37ec671a16690358258debe0e835ee34ae35a151279ee48e67dee7081a8b1ee469abf2e2e8633ca8dfa4a2f353bc33507f2af61e780deb08109ccaacd251fb610c4d8b21b2b8d2af4df1279a54fde9d7c35f90d85ec8094034241127379cd6e0006bd189425359844cc42defabbb52de01ec17358ff9d497ddc7e2c31e0051913c97dc51fcab79919fe2ddb47414ae58f8013d2d57702910115ad7ca7b729293bbe36439110385a02165ae1b5a2102ac8fd8f44a0b38133b9e31484b6927053a0053c951a97d4883e95cd36da11e8ee878c3ad145d33d45c5f8b1092ba80d10a005036dab518250ba50d0bb8901ad2926f2aedade1c93d4295f0e419716310583bc8285d2c06cb9f579a36b7dadd53a9c95fc1d6df7b9ecd8c0e2675a1b6e591f52ba986d65a61b2c7fdd085672d0ad6d5f9f1f7afe112aa1298017a2f61df15b9275b57f6ba70b5fba9d85bfed5651ae8a0701301b7f3edc24c9589e53f004c04c5d0f0307cc07b4df47a80874cdd2af13aee58ef4ee58cb81505f21b60ff7d3a03ff96b61623b590f86fbca77d4db269dfddb574aa0f68b597737f53b8e0f7d9e8b16535ee291961b1dbba5f649d976403f27a42d97b2036605ea317a10c5e7bf43dcd7755f5c14fea82896677273530fa08978190eb13ba334bd7f6b5103b17583e7d62fa6acf0aa2f27e75fb9d04b34592aeb81886715f7d89413ddd07f2b92c06779ac4f94ccb948b8d44676e0614d83e13c3826a316817584c2941bbf9ead569a79873e523e86bc40f5a89db67558c7994a2290e677d99730de57bfd53426ea16512c78b2fd90a6f016ebcf53db00601f98f61b4dd5e2d9116ee5a2479b205a030e52fd5fd634a0562baab6f4f0ccde8747b96df95ff59169f21b2e72d02667806b58ed6802cd5916018df2db09ee967f9fa7816ad202dbae5734bc5cb1a1771c72c5326416cdf3627cd94fcc3761a58fd86437ec642bc980e5d350b6bca19fc26f4f68ffd1a1e14c80b992fad5ffacb32e3400e9cae37403f88b1835d2aa449f9fe93063e34f78d2e37df2651cddc8e6594657de4b1720fc5efbb72c17a8feef9dade20f5475196b6c125f034690f39b3af0028b12e3cfbcc5f090ec8817b0a0945586a9d61fcdf0225da4d52e8ad0471ca1c66b189ef4b9ce2d0041d1e8824d7d781e7d7fec2bd6e802478604553beec020a7d8064b6044545bac80475566ce61660b19507f5d6704cf36ffd8fbda1b497c59ae89bb175500b5869d3b3db656a43da94e1cc58c54b0a5742b3f056367f75b4684ccec6136539ff72de190111a5a72d3c9ed3a8c5bb4ebf19f67f4ff5446ac2ec840808a911ae3f59486411bb90fca6e6cce8b6ac7c1fbf0197bd807f84fc38d33921e4a1dfa632e4e3edc709fb32ba1eb92de6d069f549e92b14afd557a20d9d10e50ba99fa787b1bfe539c425b398c25b680b265f1afd08f97a8ae40c68d1bd429760689683d4d6edbe7138fc11cb98f39a7a04d0d390e9d0e920440ac014f426fa557d4f1a9c15b903492f0b8c1f6bf99e977e716d3c08cb7a68b11c0df85ca14df45e1871908523a9f8ae2b308cfb83747b9d94039f18e4f96cfbcdba536ee114a2d1fcfd413da3d65fc21f6c4eab7ce42ce6668c051a18795a27043afbbbe2a0b73a218a2c87800a847f54ac590a2e6013371228a4fe9b5f69ebc9e2e64396252c9d61e2ad83ae5ab669f2f6125045e86f5111bd19a54a93c3fb6a8c9fb5f0b75429418b50d661351be3d367b0f6002d48485e62c3fc84911c39e16fbd67e51786674afa614e1b2f99da453336459cd4ac69de01a3d8bb9de6ae72956216db321ffd16f0bf9c77f724ba4ba6fc22d483e1103dc3539bebd3a1e332877990dc2a2d8a858c1a8e3b6ae93d84b0890f268fe2ab08dd25844af40895246b0895ca82b95ca9de9ce17528f0dd34f0f0f5186869cd7e3fc7320fc46b5320918ae78b42a905f50865c575b908ffdcccb4a9cb4ffb55e0b152107864dca72b4e93fd3d06cf82d8e8b5e4219e79a5ec47944da8212843bc857485e0c69c5da6ab449ee5e42ae93f55a3718f0b371fe8d7902fde9e40123f9f66c070bd7a9b8a03d65f86f41a5ddc69de503acad776895eba016c79dc7fb66df8d5e36c6f67fb985e0f6303104ceb9177cfe7a5be7b019158350e175af3935eb087d5fb25ebb6bd80d406a189e036a346afdfa34ff004a17ad75169f09af465150971492fe8d38ef515a04af8b00a1a946838750a05d338fecf3d0050e70cbdcb0bdc03bdc9026dad64e7ccdd23f4f4326e42ecdce03d1c036fc64ef199d72ddc3d3d1f0463fd4496a8c010314b2aba4b4754b77152f03e27408cdecaa8d386ebd3d74d498607c6e2eddc4373249614f5806823edcabd568919b199258812a9e2230d4c8c4ba3b58ca676fd99b7cd1a6b88da0f2605aea318fd980d322af57a7fcc7d0f5337b08bbbbfc9d867dcb2b51355af6fc346ff3ca628c81d60a7d233052b8b0e1442f5902d82bdc8a63c34c3bbdf3b65dff6298892e2de7ee4e9fa039a8bb413958c795eb70ac4027a06d2d1bb0142f49c22a20930423dd036a5fcc90380c188ba1860b7d7bba0069c2e4e3295bb3c747de52fd3fc9f1c52c6881f56cd1273e471a7cc4c9cd074749fbc8167610aca32ea0366d954d705e499554ad010606d34a1651fa08329f3f94255ff2d81663818cab48b1d2c5a2377189528a46248c48075c76a229256f4864385dc98ba330dc312e217b30bab97b5bdde01142f9cc985f95af68c03c423616f1a5ff48de9b2cde5eb30ad8d94407bfd80d827771191f0f2fab804ce37407a585c4700743892ac1297f4d8b4794f973d277d2c6f1a020d4b63f062280bc9e615a21d24b46ea0ba62c8c9619bff56ef0187c86e8545e1a9b4bf1573b9112d1951c8d27236580f03e386039fc72135d1d734e2d6af7557954c58e91ed64e65df65ac92adf968b6334e68373bed98b24d113a2a63796141027c24b5c1acb0d2277adca6bf5875f864f8dc6cdc0289db0f6d56d7fef4eca72073e34186a10ef85b30d156c13016e796bf7ff70e4813556a3c3c84c9b7010894874ebfaee04e6e0a17a581882013bf8cee07c9efe084a7ab6bae4a2b4e5faca61b6c2643d7ad1ec37e31f11695cde6b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6f757caf2d5f3f49be9fe4268e51031a9fbfd71bfbf5fcc94ee027220c010b7783e9bc7e3fc5bab6b6f8d4e4eebb9663a1298234162578d0f8f59bf1676659ab7b51bd078ac6b1600a651dc9e2ef6b665a874f0421930b59f79ad46ac4a698a2941bee9b66d5fc9fd3990d418b3fd35383a84faab5a17e42a427b71c85516746b5a5dbee332b76a71974cbdd6a6d10641f5649b100766e69a78c042deccfb1fd8d2b75fdd785c60ea6d5c3d864f9d8a72d8165bb892e10c90b3fb14801f5ffd6ee1e442911e3e77a6bb3778cfc90838adda496cc5f9a2d00bc82a9ecd913d0bd84773dc13c8fbd8e1f8e055ab5f77ad80fb53d2204f010fbd1a88d0a8836773b2239a9abd856276979093de119c71d65d6f9216001d0d67795aff82f652b83638ec45ec44347cb0765ee72d5448935dc3ee9649bba26dbd030d7613906279fb20bb2a3372c7ec4e5a83840d66f92322e2675a422bd18c416b943522efccfbe5d0188bf8e409471cb1a0c210a12ae0551e24db484f8c353a3d22c775aa717d2d668503447902e13421f3712c6134f27b9b58b2b3f2206d7ae002f17b9e2f7d22d0d9acd5567202977d5c6ef4f26e40e973dc2cdabd49fdbb6b592bcf11c338b8a587b7a0ed9bb6cc630b125077dd2685d22c004954ad5a547da2f2210c861f10aa76dc26ccb890cbdb2b8a0e202ea3b955b47f67f4556f8163b7776fd5474feb5d2ce23f53754b8302fde846aad253d25d6d3dd09ecf72a769a8af25881cb0fa0b3ad5acb72c344752a156245c590af0e4cf780a0018856527eb8cd9d4d0d69f5fb61a5693a00eef87069b6fca3b702b7223f27b71674376f068b98547b92787faf7d5cb3f42c0d40b30ce43a1be645029fcd4d3131c4810beb57bd1b7f05dc83c1f640c391ed7f300b34d7a8c8756295f09e17c874a1bdfade9e09164ff27cb5964755f04b591a07fad57e72696065f2c0324bb17d921e2dc245f23fc8fb57da41dc6b8f7c6671b8983dcec9010a4740d8bf7be95fd525d8f7bcda7c4e5c7561d16545fee2a7b10fc24455b1d69bd3bdf057f5b2c065c8e3528bd4ff5f4ff22508e36801c9c49c00dc6df57491ee8227ab230ba2d94d9f282356d4e89004debddd3c58577363c2c8809af083c730efb210994f44c64ab1692a739f9a6a41d77abebfd5022d5f56d7ae465b3fa5cf070cf48760eeff8366a5f24e46bc37f1b22af191d3641d7d66ed9deffe5bd80ad520944e308aeda0009e871c14942c8a9b086fcd1f6c76c3c11f90e2343c8441d3486bcfe0eb7854c076fe4188a682c0ebbd323e7a342d2b14456c51e561c4b30b677fbceee90ed9ddf3b49c16993bb05d62e08348c14608d4eb16bad6eed045092dd8438b7f03d56d1b66a3edac565ce6fa79772c7547829dbfa79ad4b8e4d787bf84719583451608639fd3e3c951157f14a5b8409fbc811ca3ab1be39dad7c49aba96e320d5c8043d90bc11f15930a721dee2f26d9c9a20db9af5e289fe1933ce5fa53600fd41ecbc2a9b917b996e24f806e0d18beb8558eb5379157f743273e777bea6c12902d6be63f1ed3f12b6ab3b08b3eead15df3f56e3a78b76575249fd5585550c7b166eb05b0db6390b1c9f811dbfb1f2f77c17e5ebf83c311eebdf1d1fdb1a4d5c7b1b8e04e190ca41352995ec026a0b80c87e6e639d6dfdb5d830501d564d6934496f6a84966379b2aaaf8eb5ffa05537b4382a9b282362e8edd91441119073037ba304ca469a780891ffa1a2d5ba75b98792c9fdcaaf3dbdb9c9a0349886282282c12a0f08d469f3d07157c79da557a4a9080529defe7659d09a61527983125b1d56a214d02e77b482c37ad4b5a5fa03ab19939020fff7c399f596d1b2ca7ad5e64a6bc77c8a4ad50f6cd520683b78c6650ea4ac960aed74b916e293f372cf2beea70387b1c75be3bf7012ec9b7a62ea2cfd60d0fcbcd35bcee5bac66c843db73e2e44f8e44c6ab4aeb4ff6bc500d8bcafced7aa370b7c1c3bf8aad31fc5c84ea80f548006bfb0296edf4223e25fb1d248a6c557bd2306258ea8440751ee4922b6706a0a1f1b8b4703cff6e880b6e1447167140325dbcd26b96c42345ad970fee7de638cfe8a23690d9ac2e225daf452a940278d18d77063a4f21176c95b897600efdf2d4067e4b3e55939302d3a58a8d0eeaa97052be91d4e4aeb69d50674185730233d627d993fa84ec050b82c0b6e4114687ec23399ec138c4839a5a3a176bc5307b9f5202c7bd0f418a9727a374030dedd05debde47e2e90b9b3c48db0c0c54f9632d2b02fa14ba92c282d48e1f34a9a303d144d64787b93ebbf957d065dc450c62855ac89d2830db1066695358bd0c2e04fc880e72143e96c350bb5962b140279aa1ead663939d043f90467a537146b016fbf3ad7673b3c598cb3ceb07ea3a93b5d26661e03d730ca651b87f80bea8c1c5abdb205406ce0570b16d0a5ef8289a311301ce4cf8f606950894d47e1b008f6cb8742911e376851b8b4e2126e4767a250ed1c7ac682cb19c611d54b5366e3b0db670ccd9cac034eb1bb8100bc7eb097ce1a66f6fe0768b71eb1bf4f63f1f83d92312c0eb6b3594d9433c26868d9343ce183138adaf2e832c8ecf307e420c1e0c45b64571a00cdd4086cbb8aedeac7b8af25c56bb88be996f9e0fe580d1f1ba37b29e92547f9ee13006be53defb150948c03f26e675882ac998811cc3c64b579c087f00d92ffc82d81bed65d06ec84f7b0618d22f1b3ba8e1ba25ca844bbd321aeb045585a08fe424cab7bf316577fe118100880ae19d2f2a3036bcc221c01a1849a9365ccacaec4c96e31f3db248e23a808e796601f8b405fead5483d0e7c92fe383ba6f6ed77d1068078923106cd8a1e5e0e566f7b84f3598e71d7cc539e162303f018a4af0fbc12d5788ddcdb5f73ded8704650fb9bd3cb9ba2e338c68729c10ee76e8ef12d1a683126d51a06ef30430a4800f07700b238a3f09f8a23dca2964e63150b500e45455ed9cefa9df16cb2a2f23d232f1c29704a85b713f4b51a5301484759eda01e8108878106fd1d7399c4a7c054c1de69197a16993bc05f36b4c39b45cb8df81a350909fd269efdd92792163112f5bce3a0fa29c5fe86a9bbeea67f37b6348e6a1bf5988099d30ad8a1c1cecd68a2270f549ee7b235b0ae2a06f45175c577d5909ca9dd0dc15000c66d3874895d8a9cac2aad8e413076789221a9415e5b20f1e287c434757310f67f42c102df3ff64a9bf9999756abec2a18b4f8f3842470b24c8c951b2f75f5055096aa0dfeb3a042af0a8a0f5f35fb901a662220d871bfd19f081cbb430aae0fe707c3156a13536107440beffa0f82526421b0fea33cb3da02010b25566c8b9a8216a99409078526be2e5814161a6140187d48ab5966f4bc5048205d8cb62110159aca05fecfc555662031470ffa75cd7fc848642003e4ca64a47ce0be2aa85a6b573aa192e6f86eb2498815ca854b95b840b94b32d38c52c19f959a514534ef986f96289c09e3c1cf1365a60a691051eb4a8cfb55af7197a257a278ea80a114dbd15a7296fd205083b56f0dd319b0ab8e00054adcc31e276bc12a9a7da1c186e5283e187ae36869875d19ea023fc8d2a43e1572feb6d7a0edb1ac4b49ef5cedfff70c354a841a4d36ed3969ea907acb9ccb349d6a2de73a7a6758041eb5dcc944939dfd8e9dbd8ee1569a32614c0cc3acfc420fe117a6e66d935a3ba14d9213b44fc9f9502b41b3960768c7f599c465773d2be3d1de326d10a199ee436d4b53365566326e4e37a02e4e7f4ba3167fa94e3cb91abd16267503e5890f2fe1a2d5f284aec959457ac217f49ae3bb9e144e2a9ec15c31d71221026f5565d7dc858479695d767cd5c3ba099a474c5beb4e8615c60d3a05044169bb204338d52d0dfcd25ce34ec9240bb67232c721a05e6de49e6e7b0039a5fef053fcd63bd8011776f9610a63553fbfbf0ab1900575604289fe2e48bd6b44e77504c63b8b77fe1e914ad0272e294e1291e43047f631ed3286298040aff9ceeb73ff6328f60b3d35cfe8e298acd5a91894b53b2d4428052cc2212d497839a25a676982ab03e055a6d47eb2fa1f0199f1ed4963ca305afd47702063a3f42641ff9b1a984a8d96f07c0057614941c076a5beb3eafaf71eb5f10929520dee889f8c649db101e825ec2eccce2ada199e0236f9e8c299bc33a066fe15a755fb9691bc7a411b4bcdbb916b42a6a32e555dc96ef77ac486df11664d721c721f822914d60b839f2199e0f51f08e534675531ab9c076d3fe811cb1827da8c6161981e3403b89f3e95dd73b67c035bb554770bbafc2d11b9113386ccc2f5d80c67ed6bb79de091bb1465f37d91afc1d79d6a59585ffc18ffc9968c2e04a6a016424f863b1f309e990253c95a6eb64cf835b926e0e325cc02f4d9c4ab5fdf0466425f8330c0908a85e80d2ae6c72297a11137edd4e5d7ad0484baab7176b1159c580f40c72168e785fc3200bdc319866bed5d7295caede997fbf9a87553b402d26e264da25102420bd8a1e7f64bd436c9c9106ff851e8cad4a2e85b7783643970f05c470cf2eb2ab7b46b39878773514b9199e2cd55af6b25d956911c085725bac3362a7f4e0777e4f3dc5b0617b798cfe8bd5dcc209c5694c344caf14f3172bf8a7e826da22869d55a4934ce3ec571c1d4038e3b28a30694aec2daeaa602280953654bbd98514bcd918814d96588298f7c9d44f250a64d5f862328d4601cc83a59e97045dcc636dc24bafaf5817e0b970d316e8c1ec0cd2a388854caedbf2adefb7107d702547ca21e781ff4194862ec7c31fa021bc513ced62e9df8677fd04e6d02143c088ebfef9971c46624a4aedddf4517516ba66fad4d68ce6f3412a06f3083bc42fa81e87195b399b71df99cdea31c886fc07afc5e65465d356dd501ef28cf5464d9d250e659d6fded06ef9517761a7d6153065d6554c2d36ff54a5cab1b7e7e54d86079597a4b409fab9948592ed3ebefc793498f46dd18258656f28f1eee5f7b42d5786472bb4ead26162d657efb8c7ed05c0c8fb442286815a393f99b8319eabe83fcf3d848ef115e79609063c96471f059b9e83c2f29b6629930ece71bfa47a9efeb770310d06e539bf636a33f87eb6f104e5b44b854a03c7f9af606b3bd0fe416c793f26fc58210fbd10f24ccb1d02ea2517212d88e671a68838f172b9fe2f4c61a8c4f510ca70d232f2cdf2273d9766d3870ffbc83894e3607e6a4f85c50b96c84309c8358867a198294a4063ef66336c12137b688d4e92f3c2cf75d5122605b36212d73d1ab49cf8950f25283e64f2f124b64c978551eeeb92ed5ecb4ea99d41111777e72a6458aa2f669a81274324b6c3e4e6209691127e2461c1f9c300658702fc070edd6fd340a210f23ecf6a5b9769893b6916c8263155bb855f8a9cc8b9a26132ab3f264437b22a042bbcf4d158e0ab82e63a87a3d313e3def4223e24a6b9d462a34562040e88751a69ad2978fd635674c34c3b89b56e69005d6d0c021325931d459e6dd0e8f54c667b0bd7723aef51af8e185311415fb336cb687bc1ce10106d42cca762b0cea8a12501ca8df7512e8ba032f1c1e0eb96c6ed6185359e7b3558a6146b035877e179f03ca514e2640ceaf217afda668929d074ebed3a5ff135b26efbe8a201db9cff8843b5e5e585025d664cad2e666ec7e4b45776161d177d0e4c89a3e624be0203e64fdee00757595317c23b15514e8df835d2bd14e1907492224ed77293367e6054c63443269;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4b69f2975b33a7f7b49a55d87779bf9b6324fed634daf61c46432b2a32b4263fb2ccd4dec41be6c01850f0adfb3d22d19a6b808992b4d2261672eba1b117909c81ba22adb3c35ea2586e9dc9a4975bd185f0d700ffa63a3112abe26b30bd69920bd3cecd16c8118cf49f6686421caee7c6622f5f4554ca17f5209186ef0e1652fa60cd9730dd76a43d27ba60f2359caaa2e7e390014a16df9306c14399a87e10b42046e6bcff80c4a9f85c4861d6e4a7597f75dd768639a4d1d7ca819e85a512953f46917582c6cf2c9020bc6387084d854b34d89be9efc34f1dd215230bbdf056619f7cbe18a5e501589074697b197eb8913f811ed67a63b77faa23315b27b881c9f6c4e7a487ec52b0d0b52f7219027fd6b33017c8df27d20015e37ab881c37d1430075c26a7ac5e24cfdffe3d88a0eba2b12661804c85eeb3340207b6b6f44bbf2538e788c6bc304c811e9a93dfec168c65323ec7563be51c80236be883938cb754b15b42c86efcf5fbff636ef584815b97c5a0d938b4a48c48b8f12987be7e66e0d7de78a35c1f9cfc87e0e53748655ed0333e57b6cf596cc46fc3c79d3ba3317a9c81db27d37ccd42998114172cd6993cb4679fa4bbf33aa0afb76c451dce63434dc61ec38c2ec31a8fc70f1c3191a2f03ae1c4c73b890551e816b957e697058a38e9f791005dda765a08d66a424cc31f2261ebd178e5285af04f076f8897d51cba3e647827691699681933dfb008ce35189cb8bb7afafba6910a2b328ff869531dbe693479fcdfa52a80b3d32af7bca88449387db476f106e7fb0fe3150b5034bc3075f77e5995307df4aa83ff9b9f639ad441106adac0374c8cec08467cb283b89ce470c9df8f915f40d242898e3c441a9085a19b318fdf4ee932c1ea564f1272462d3bde81984aeb92a7d70efc63021ac157dbd35d0940216bc6201a72df52ad3ce490ef4827ceba7a06a9862a63fdfbf4bb4436c9efc0c6cc365c779b673dcb12fbe1c0f2cc89a960c3a805c9eba71cf3c374e5e9af47e225ea889719949a1be4b64d431dc55cc36c66a2a617aa075dcf2ffb73541c9a9cf430b89f89d351a3e722486b71ca7f91000d02d45452bef89779e01e9895d72e4d08c919de02eba3906907070e504b1ae57848a544701b508c6caee7a04446aff35f734b32b8620f0ec79aef7f49998c8008a71c4c065b6e16eec64b0b59003c47d4f912fa2b1eaf1239e7b18ce77d397f8720933aa34764a45062f39b3dc556dd5d9aa4ecb9ace01d52f18b24dcae74b72f49d7d610be034c8fd167f8cf9927d2a2dc715485b8bc2533243b04acb62ca93ae4b4ec458d51b8dce464768021d171cf63056b4de748cbf59807e27972b8d4930c7eb5158e53a6ae6ce401ed66c8e01fa7484af4f186202d468f13b4ae022198c8dd6cf503e426a3093e1ab63c0bda6cbf232b4ccb25988df2be42e5684a493f9162067997bf5ca1deed98dea971f45cb64a307074ac3d1dd8b141cb0e77fffdab3673440bd2e275e9d7eb28f20175b6abf05b306507cabbaaece43cacc4a1669ccd73bfe1ee1b81cc74f73717afca852bf2ee726c766518ccd72fa8d75b50e22919e2967a92697f5f5e4b83cdda55da9c5ed9093b54d8159eae94b4ed63bf3b96493be2a551b223bbbf7360095c3d79c1865a328b00c79c4f5ab6f92d1fd4ae1fa0ca4f1c0f3dc5e31f0fcfa683b9acc07a8e8324cdb9c24dd2e178f5f0b35c3ddf0e5724b826754bd6b4e263006cfb34c9f4b3ee91abc74559cd203a471deda4cd661f20efc1afa3f126c214f3918d5e17e10165e57299065c396e5ac109c1ae599c66007e5c34979721abf2dd8ef80628ea5066737dd69b7fe354027dffa2388950b816b2375e4df253c8cd04be8c48d186a722db5dafbe5f7dabb069541a8504f48af77ba58a5176fc8a1128e42de0b15c7be9a9b2ea38d3f2d374975a627f718170f40866e6c5527037cc4e1cbed1d0ecc0a83b77b04d10446fc2f777bc0ded83f5601a4dc70456deafdd3a51a83a3143758a9e2ce617a702343c87b00cdf4d55753cc8a0c26bb9f305bea6b0d9a785dd20676598466e723d482f81b8fca7de22aa19291742861394236977acfe0659c1179e6fc38ad1ccd59fad8ecb4d6bee850ba6dbc563d427fb40852f10b632466fc5284003b19104ef30ed1601feb38a791efda03552e6907d50009ae787b6bd5560b56d6ab8fc50bcfa5ee627b74c7c60b3a0e25ee7c8c0a086148640fb4d07f115048771809994d679a66d978d2ef201276b72d0eef033cfd949f7270ce70477914e5885a12a4a492f5c7b991b015b99e4709b4488c60c5c6eb2201bb94e02a54446c28fe99cffeebdc9b3ba6603b9d12edaf57b99b4bf0fb7375ccdcc91ee9245a6f821b988cb42db30c4c3758078f2564d1d9898d48eda593c27f0f6b27455d7337711a6cbe2e94be354bcb1151323b51c072591fb82e9f88f75e0f661bc13207398c294cfa760c03c3ae489174c54be6be94aa1b9e29eaf92962cdd2de43d3c3928b850834e3582d3c10932061bd801a2e08044d8140367e95b911e2624980b70bcbc4db0643937a58da1861ba67349e22cf2522e634c0b3cbb32ce99895035aa353044ea588338f9e867562d879fef5166d246a468cea4d0bec216a75001de95a21a146056e334fbeda18440590badf3539038150f62b1d86bfc44a052ec8d9d4fe85f885b8fb0277363e26ac227c0282037417dfa7f13fa025e17f46f931d4f634c629a15ef266d67e09680adcf1aabef3248680489b984f3ac590537fcba3e87f82cfe21cf7787c94027c8ac5385e7aa7b6c007b50215764415f34cbf5e999c7eb391c4ecf073fc9c65df74bc7bf650ac9a332755f2c3c590f82bb7e2059649880c942f6a2642d70ffa22df9b31772be2fa1fe904376d7fbb7aab77c53f3ad50a7a855b38985c72a409705cef58f2a092403876a1609a449129b0736b5f5b85dd4398da7325413cc7ee6151a77330062b1f85fa18aef94168bb91b6ed2574c186d2a0048b11f81879fce31bee7e8797597b85107cbbeee85279ea90ac161d13f69edd3941d5d8ba70db3a3943e6fd91ecf08b11150a58d4c750ffd4be553d17cffdfcd4e17c70a53be6e2be1c5bc989a51825d49d27b6c138f21f4790b5fe84681de6442d3bdf883b5156a6b4a4728e5e5e2f6df367fa08eb0b072e2b80efe10084d2c94f812bc5d3b64374c5efba7e40d2fc6af29e997191df482c461f127e211f07c5ac46098990872678871af576abaecbf9be0ebc0b7c3caccb1c79303f59e8963107b938854e9616c50497f20d0f988a9e0761db4bf96f841759f610ba33e3ffd329a6e1545d8f9801774c021af2792f9bc9805d49c7b0cad4e5c99de5763741ffc81cfe368cfb7affb185605765a19d206484ba0b9a07916a9b9f4e8c16c5928f06261eb0e1a12a97a84f68bae57ba29afe576cea6c9cb5bee13ece64f24fcba81518cdb4641db639ef0d2b49430ec3e5d7e0784f2b609f420676ad42322f2a4dbfb1f86f728bdb6b074688374decf32bb785257ac224a76bcb59e6c6b3ac5fef7dd849c3e0f7e338756a21309b53f84d233679a273549007319fde47651aef3c33b22e5c7838b22164913bc8285edb07040a2bf9fbac0b5b47ebc6561d50d53bfd803fd0de7708fb0a230ad6523e82bdde180f025709cdee22c6f607f99d354bf1895da758ed1b04fa69c4c5ccfe14403fafb2ad26d4d469c401b9977986310e0eb04cbf38b1913f886664484f35920a9646a4f6bf8e9da2f68a79e66efe892f1fcb9e320bd446fe3ddb1594b8a2baa1f3fa4dfef94a30b23b94dee7a26c900f450bbb61acdec68f3d0de15b7133289e386182554bb4041b24e23f3427bdff1b8136e506f48f24f065bcb22d252c5121e4fdbe4efdb4b17d273bcfa8e5eaa475b908db80f09f6924287ed6d79033db3c4543ed3e0d3db41daa16d6bbd88929d3ae587278154b8e963dd9cf31a6cef7ea376c35f7c9b08c704b49d300ae24badb03565f5e0a82bd2c4c46608d6f77d490e3252dbdab96b0806323a29d7722e117fdfbb1ee3b68c655425b7fb965a89e3cd71863337e2e2235b691ea93583bc10f12cb4ae81790ea2835d0b419fa829f2b31abcab363cf6fe80744a3fb678db04f2b0a1b0cbaae1bafa740504e810ba0baebdbd932b976cda69a0011c41c58f09ede6b379451980b928e77d67debcf568a292c239e98d89db6a8aca9581db1e77c0f994b1bf28cc4852dbebcac729ff329cfa03ce0ce153cdc6414a06beeb3b19e619dc05347d6599fab52162744a728c6df56b46d1750608c16c784dcd1b551663317d438a226c43ad824a052179f70dd949308677e0379a5f6ea4316812fda32a52e0e7ae46bd2bc1258c8de7ca4b950b807c02e7bee03483929266522b19c154b4471c428a107f2b2aacaecd767804b7cd1d75b30f5e1fc19d31126f6e29b50dd1118385d2a8598c441248b0876606caaf37db5ec8a1f23de79a877ffd91ac537082dbdaee2eedc99ccf5af347a6d73ed0e49111fbedabbcbac8e3aadb34d4679cf3fd27fc1f1323bc9aa963c1c4cbcc21078fcdddacf9041e91a01fdaf91f4b2602074cf35bbca68ea085fa2fc121bf605b45c5f2d867ba51bea0451004315ee89be5208f6ec9c27719b0bb8325d3a3c384e44744af41049456edef4d984216a3a7bed0a2bee1f255e9dc3ac05440d6c4e1c16352dec321b6c76f433bf7aee8a59ff6786fa13d44e2ec43bbecab863e67dcadd2d26c693b6a48656d5c8188bf0f8b825f4cea8360fef48fdb7c41ef449ae6390ad6fa30193e69a109a3899383a0764a093f3833bb21780b093762e2bb4a8b0e0217abdf7855a34e27d0b1da1365b364f67607549537ff36cb3ef26ffd52dc47e89994d0706b8e3f885417c8d907b91a05e39ecec0d9c0e297018dfb36c86f8b554f96dfef21732bc6e93311ed6b45df1425c1caf5596ed08ac4e2f6ae8933ea2ba7c191016e63bcb479b4f8caf2f8081684af127cab5de890047f12ce7ef9703eb4b6726378c04122f998a0a33f407b3379fad7d6982853d979ad86bc50dee500eeba4850485f607e110f151b0aed7f4f4072af5d11453f5ce3efb986e70e025219c0bbff06865f93cc4c7bfeebd985a74b6ecba56cad3e0e873cab75e80a7ea55fc9e43cca63d1a4a0d81d320e5f55961b9054fc0f0ebbdeafd32ad4078dabf2887790922a9afebe5f02f93170741144b9b359a43566bad58a9ab253fc0b886c1baf7d0bf0f8c1f168a16076fb697a71963474943787f208eb173b1ce97234c6a77a69f65077776230e20a388ce0012112ee02f738bc6dca17f61fe1b31e482e38f0a687dfc9749ef9abbbfa2cfa5ce6ecbb387435948b9f9fab5fed544d592f45dba2ddb7d14bf55105161a3edb850239f3345270bbcfa16c42138b885b95c36869b65e90d5df537688263f9f9a27e12f84c13bc17864a7aa6f9bd000c6844cf88fc81db5b263171ead29a1a4f69030f3fc8625bbde561ae3fbc739ea892074bf541f508c618d2995f299fe1a70c0f18d50e36999200bace3ad604c0e34f9c588d7ee3d8fd3511f0cdcca325c39fa6436634384d1b4130966a0d51435db280d0f7c5fa77115115e67732b1ded881d5d557c2e10757b7acbc948d873ead0abdc3b75fdc27e97f140fc5c92326a1a981b2382840545cb1000919a6f958d3d392f98bbd815b1eeaac7d57208a16627464dafafe2a184ade7b9725e9e0433214f5b5b7ea476;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he47863d220b068c9eb5f55cf8cf103fbb705a7c6eb56614a0d3e4be659d46f7b11078bac0722a4a9e58b2f9811a5003297798cb60121b314312a52b71486686e81f6097a2e793f8bee444e3672ba9c69e22556026127ef2a5ad742e91e4b6a122520c704da23049f9ba7e36e06ba5a8445781c6b637fed1b25182a22c983f734dc20ed4738a3877e199d18c98b2acd000c245b5d1119ed2061745b84e0d5b329af8216d2e011e9c287b55980ea0aebe5a571f2b32974330926480fce80feeaf311de8ece947f8d9c4da929163610d7ee6df46baafd7729a7dd7da9f05251c5326fe7972dccd7a0c876d6b429449fb75985632e1ebc14ec75f052253c334f27e7b84d6f03e23851fde227751e4eadabf4dd81ae496dd467330a30a2a06a75ccd2ec1b0f2b97ec3dc8eade19c81df82ce8e06ec94262437ea85c1d947104519d497d29d69f77ca4755033648a68b0215c1788b16b0cb990fddfd42a4f29af0c43555817ef4e989e371829daef21aff432cfd0845e02d0c8fa95961414f931c48ac6cd43ca9143ea030214c5661dcbea17bbda04a026834e82bca1ffbc32f2abeb25468f47632d5633fe511b077a750a52764511a5b97cfa493bee5e245792fa64b6f8342f88f7ca20cae06d6d253d5ef0bf078694db60b003efd2f8fadf3ddac0fde09cd58427685bec46eb71f4a890b1e01ef2bff872d73f69ccf919da7d8c83de6a0a2759882cc8b55ce11cdacde5fef27ab03f3503a64e5259cd3b4332fd7a159f28235e1f877ae841887f2748733edc319340516b900a07c778e0ed916513f276bae78c835c33c86a24e6329372cbef2a61ac9fe1428e7e3632f9734e77f1de6a6b69fc5f8c4b43809f18c0a723d10d6b724112f92831bbca0206b786a4715acf38c58e5fea2674abee06938c1f1f0f34f8e2da9f46f9bc4cbba83356fbb06b31f55aa7d025f8a15db7b025e33c08c2ab7cde247acfd347a977ddd1dd273ce7965ca88275f84748e0959cfd985e396fdf01a24782fff9de9989015f2613b775a1461385a034e95d9acfd5c78dd72a7aaff55d4bb6c7c1d575e1fa5cc5e0345abb1facc1cb2056903c8a68759ce0beec7b92bc7936b6a0628cb5c85b7fab2753791b14f875233ce159eea32520c550ba67b466ea04442496f833659028ded3125319c3e05701f36b1d7800d10c143babd2787d0b26370d2fae879e3cc1c3f7ea68e5b1d07960003f8fc27d2e23448144f16b9010dc977e144693a9c0ac2a7595c6f087006aa7f88e82f24c65b33397d33dd1297b3408786206934d708050948c5829d7482734b2c7c1fc09e762df9db04caacf80259ddd3e965317535f851b56a6422cd292b658666db3d6d1f6680601ef68a7f9e9819b6d18eec68aaa96ca3f126d1d338e7ca2b0223930dc81370a34c1c690c2411ae14337de39e8d48544fa66008bc5f16d3a2b5d68383a22f64faf6fce3eeb5d86ed5a92de984457478ba280c7f83216488d65d943a5995bf4ae7ed7a0a813fde4d1804cb07a88090251e4ba4b68bb301cfd2c0ddf29f97cdef0eb94320ea433d3012d53a9583d1410964be9762533f151b3ef3590d01aacae586acc3f09e50f0aaea4db269cfeb5a3643b34b3787fe8a6fb00bbcfd1c6f0ea70660580676dcc37e89afeb6e37c946a4bb54629115f48ad3a149d56abdd368143b6c1be8f6a178de46a2f8753fb162943768f8dcdc7095c5845858dc7a1b3919a665301829dcf5a63a7850e8b98c1b3a1b2dd86b0902fd2a28e2d69fa06b55e59f10601fb1ea14069d25fa91f45dab354d00cfde5d6e1d51a809441c42dc10f51c9a275dfadb4cf03d8b723630cb65fd31feb832e28a180c290ab0e6029b5ad985ea913d026bcdee508f6c9a95b73e76fffe57db621aebe06e8e33282f37543e3bfe95507279cb8761e56f350df285a245ce3d59d5f6991e549289fcfcf22a39c8f5bd8ace02a2b8a3fd615e181d55c7a19d93087fc16f19ddddc048117f51199a4c33134785b170c93ac9eaed92aea122e04f04f790c9771730a9e42b6df42ffe4973f850fd20a8199db6443808e3a11909705e52ba2bd88a447ac4c69c0b68c4f0e972d7986ed1def6e92ad9b075d8e228e1d7af65b4bfa7683108d50a2556595c6f32be23a8b8b8c96a1523eb0afdbdc20e3ecf94bdd0995802e352f7c208d4ad50152183196a255f46a57a7f1e12c58a4073b6b07dcb247d51e21b15093751e1d90aa41897e6c1db6b7e29964964c9c865972ae7635c7c797e28251232d2da0ea271fe98937fec3925201a5bb7a7a35106e126086ec6f406cd0ecf2506b909b123c9ccf7ce4e3a9c39a401cdde75a6ea3e0b51db7db0adc6a63d621eb5665cc5988a78ec054180d5a799e6ede5d0c4b8c82204bd662b49d2b0f8327df1d309eecb53b823231be585da4bf46c4c5ccefd40dfcc56c4e804b688fe8f1e98c1e2cbd0b6419de6711d1141c9c2f4ba189fc294f198294a9919ba3ad81205469dee6fbeed318b96a4e9f036c00735de19b04583b40f1146bac01654981228927112e41522081b3f933c08b3de87a0de7262a1e117024351166ab73341f5482da0958f5e2fd558aa5f662b66b05da9123506b66758d93ebf3f039203f7bcb8ef2894b450a70ff65299c06ce5b5cfe5fd66156e8258da5ca6359a1b88c7b27bc3cc92b3e57b884a6e5abd66a1a112be0eea111479206bfdc873670274bc9db54d21fca301fad144343ec93834b23d7ff511880399135bebbabbb3c886a49e46df73bf273eaef0f4251823873e12df033b98248fb60cb65063cf03e72805d9b5978646f474d699edae45e2ea94d627419d5da45a8108228add497485c31a5813750ebf848e14d7eac4e78d619b7c945ff2222b3c3deec5c231f1303669129569cf07d8e8451ef8d5ed98f49873a7dbe3cc61010820d60e78ab2a4f1f74e3c8a5b2a9a0858e2086cd8c4f8c167663e0388190229bb0b4c6cbc9a0fa3a08252593206280fffcbbb10623f249126550ab20a0d89b93f70636dca36bdf5b293ef11a8be511d325c24bed38f25a1e8e44225b5301ca9e34656bb43dce6ac0886393a4784d073e43e2871d8c540c53f0ab0215f29c3f4e85c33496861d976a8ed533cce01065ea080c17be53f91efdf3a87777ddfbb3b05fac31f36ba1b87b9f9be81614fee755dcdf55241b87435acbe15bbea24244cfe114805c95accbcf2965246852f80cab75caf8411e1d8ebcf71f16ae27b05122642f1b33ae5aef9512f427c61bd1614f463549846082976269b96e31594a7e1b88f6122d4be8738228405bd82d512fb69f2a12d2beae62d947ff8a211a954f1a03e01b90568305dba729fb5bb9219ffbb3aad0b5e90f4637317225b9746182caaf53003ad289e044cf9b7b61f1f37ba998bea9f576aa76ea7746907f99e5967e37b96bcd6b056c4062ee5002b6a183bfd54a59d8188862b6c771aa4e81af84a862e59b36aa2719b00673399d87358a78d6de1b5138d007c607be192dc97b9b156ef9d03ec2aebe469d40a0dfa81ce4c2a4b72d5b66c9ebe1d605c962e8f641a0e9717f68ccd55ebcb1a1d155e5dd3f556068da6315a835a7aa2ac278ac9ac5f35a7f6bca2a966516931f2fd82ae58f1f2928aa5d881eede675449754ed676c257281e55839a3339fc2c7b4a44cf5c2752b540b13fb49799088516668050c7d4acf5c2f89b572648f5d99ce29a5391caa9a92798373f4f1d3e7583880643f6d53dc2ed68eb4d4a9c64be7e97c07f32ad8405dee00e980270fe110a28576e154be91dad68f0f5492f1118919d1accc2c937bf954c876152782f1115e4f4a7493a9ea69dc534670c42b64897054f0411b4f3f0285b8fe864bc396b9f91194cddcdd764a7b502555c7b34c266581bf1f7b088339b678aea8754a502f8987eec0637ffae86b483c38d205f67ed2811a80abdf19acf34ed2f59b69c607927eb98b5572e669bc203cb1c426f9226772ee3424d121add380389077941436bc28449a3f93dd1b83a818e48f2f8328d25c86a72b042157135c0776e30c9c9fd78ffd68760b6bf6c3220de13b43c5ad812da9dcef9463b14d2452ce50b8d13c8bc109d42fb2f4d4e5676b1168442720e1fcb717c0d8d6ee1be8c727f3d12c131ef1cc1b9fcce7efb00819e995b5aa09a8859ee61abf8d213c2b3d3c6681ba13220d8807c0af138f525c8583ad931b4e2dbf5589358c4afbdf8f0935130b8cf6250dd248414ef445ef5c83458438bd2c21834faff3008770ad28e9eb577205f2440d84ebe6387f9d2660905aefd51dd4665c93ba610a82b021e94e67f4c50c9514fa46ed4a0bc1a5c9247050926b3b8a7cb5699364067be574b00f4e091510bdbeafe21d27c506190df05a7b2fba570d6c451a9c52544848e6697cfd2784cec39aa5d42e67d5e596a3e818885faf733919e7cbbe8bb19ba67428a13aae1b3e82eb4d22ffb4a2cad482eadd97973d802014d5f92956f09e477ed5e0e0c00fff25ed589b733b481f9c6c0f3326d51d9633bfd8c90c9fc3866803092324e2ca2d533ffea1c1424af5789f89bba913e0849f0cba7ce76aa27f95bcb5f4566e011860f57ee92d186f0cd1e7249f404e08b17289203e18341d086896372fe8969a1411af650941edc4b5b69f7ee4fc5a8cc27fa5f5d2c4affaee88a1cfc39be8dab070d26d108f2888282fa765f896d48f4d2f621a3334dc139eae9bb6e4f40f765aea4fa1d216e46a9eafc4faa60378296463ed22c094a56899415f76c9a41da802305d8e4232ab818441bee16f14a6be7fd3abe56563a11e1b075f9bd2a1127808a06343b3c4eb5cdb0941d4182abf4d351d77017a8e5d822a9293f984c9e043217c263bfc080938a6f515296a63d683a8b974a7fc473ddf4ea786ccca1d518bcbf5404e45f7724dd7d632a809bec509c96f48583a132f8a51c75e3a5b18bf7ce510032ea05b3fc68f0cddca30617a65605bc92113888d547bcc31498b665505dda7c72409cd804ed0ecd4fd203de572ad5e889984a699aee440d1bdc595f2b97b969e1ba2d9eb4e1ff3b8a7f4932d9048936d15971905ea65fe343576f2d323ab7fc131677062bd6f85561bd1b4a37266ea878bdb0785e025fda343f9fdc0eacfe415f0e5a8571b6494ae2fbed717f47b260948c96c84950d25bcd6fc7e6eb58ab31d432458ca4398cf39e0d3f069c493470f6cb5515b74f6e759dd1cc2466c99f4379eff8ceba858fac82bfd33b613a6c85df0734db06e39b4166f9915523f064f0c251ca5cc7fc2554857cf2be2f7fa6c7b32e026d6976a22a79b30ba126883089e936ac027869557d5ad7faa35e211425b1a8bf2437b48c9a57875febac88a4ad2a2e38689557e1faafa01195a4299fb84ffeb1e3e27d0e1fe578116abef993c194ff55e45d6189eebb707c48c97e92e75cc57eff1b148d897099dd51770e0e5bec46a000c96fc9202114edf6eeaf5dafd59ccb700531522d7021d4d9d040c312d53fe1014b218283b644b4a4f5b1be3b233b500387d64efe08e4e576f0dc2f2522ec47cb0984f7ca193b56ae7fce8fe9989d12e6d3c38269ad9057fcb777fd6b9e98b740e83fbbf953a1301cd27dac229173835aa156e2094c0b5a343dcc2f9dfca54cfb5641f9f1ef499c4c246bf7a877f39f1e5cccdcd48528cfd3d2385aa9ca40715c56d68427d2536ada06a5310788673f4bfd7043c126962517ba5d9d41128a5a7a0fa55822d46b061219f1034c159ee298cefdf8b3ac4af9b5097a45dd0c40394fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5990e0949307e8bafd55b66a95b9d745f902043f7f4cb2d1198f9b5811de8dea2610ff90a93037e09fb83cef4a78cdb18c829da5db410e7eac8fceee61adc3fb2b74c4c41fa9cd20dd84cd8bdce7b5fac2350e91717b52d474e63decf310a27470f9f1cc0787ba60dab643aed15538525cd318a72415afb92ffdbeef32253901020d9ec7e589bdb7cd6c6405bfaa3f7b83d56fc58ff360cd54d5c7b5ecd6c139fa522b6df69cf1175bfe92475006c64d913944d3f5249229de4828a85473e1de1c41a06cdb657be2228818b703d824580f3b4256eb30fedb43cec0c957405e9ae0b90a3083e278c52b1dcee2e4ca8ff6e94ffc3fde674ddc9db1693b68b479172952b1d8e7f8f31e7a455e9d901cf98b024012897a26246b032f48a953364cf68e61b42528b519d51b75a502292e90e66d3c43a6e91bf564227cba742c1c2d8a28da63c6caa968edde0eb0d46bc281173db9957f60fd3f13167c259746102588531fd32059eaa4e653013d5b17f62117f9ec466413b0e309bb151f3c1777422d848b769bf8af574f586e464803e1b32bd317956abe3d52c3ac0a1d49e77a7ec909e9611d6665075584f0c0708a8c8be7ac5e71786121f6faaacd3534f06ad4682e70d3dd3d32ee239090df7c92061d7e71e2a2f36722336d81b7737295a01a7885fb39335cbe41cbc5de6e763b1d01359ecb4e27314b0ef63a2c7a38dfa3180873057833597eebbb1e5414ba3bb8d87c58a80013b3d6da66f5d6e7a1536f08a53064e8ca9cd2534d4459557e76d31370bdbf9aae9dd36e3ca3dd8b379590d22049857cd8bae93a6b8a390a7819aebfc639a1ae1a7f8a1f9ab34bc100a378b1eeb8ff0edf319cf0e02b95fb3745efa03145d0596ca5244b425afb27ef67b9b3226204696656dd6294ced9cc70ec2cc1121f396a82b109fb7a88e49feed6925a08b918039112bb16e97c58bf034deec6ceb1239527a89f8c7a90b92b8c37bb4282d463bee13ebd13e3b4c79cceffd7f7404da88ef2ff5f20ad5eeb97766189d10aa338ebeebcd01fa27572e4c0bd13278700bdbf22ba087d5b8ffc8210f27f5902e18d40deca95dece291b7452b5f3193c6a05dc587cc6ff6337987d45d532c703c2c74d117a270bc71fd492e2261786ad2bf827927f3d12c79066dacaa6f961c0b1e057f615b592041e3bdbd771a99bf647076b232372aadea643bcb582f65863f6ac48117e1bcab6312c5ba15176c046e5834b43fbce0f5e8915df90bd75acc2cf441714ba63f697a345d243cdb29f4832e8cabd1e714882309730235ba95d7053fec32132a50ad3b17fe2b4e7b8689bcb548b348fb2a7a5e85e6e49b4972369df4ea091567c09414c6d4cc69a88264e5d72a6316956d874359c9670da0a1a795c9b0d3fb1a3bef89343e565f3fc0c16bf7983a437f15cd64d8672122c1fcb229a059266d980a2222fab3380017d4b22ccf8af63523ad7667272adafa08e250d523932172cab4d141ce87a7f14b1ddae7272a29935006e2c6b3697df3f80d25fe92eb09513a06c6ddc207a20b7de767e1ef897b29ce958aea2bf5c048dec84ddfbe25866408ba2fea6e33efca0f4b3ba3ed4bcfbadcb762e4022bc60d90b5e6c03305b1771adfd095971cda7b342c8bb142259d1c4ea588e6f7d2a74a436634a89e6a2f8f569787a2c7d7bfaa0836f103e47855d7f43840e988ed216613dac7c7a6ff84c8fc6e3cfb6849c3c89cc6b27307fdecbda28f8cf91c62b89bdf25952282d7184050fcbaef88815908cf81426f72de5c61f26ce52ba7bd1f322ca7174ec44dc21233ab000b485abc89015317a509fa4e0e9b114d9c09e8a125eb2cc329fc855cdfa23d31981c6b9c8964170defc67eab899153cdbf40c0a40887cb861b0831d73992f67941c6158f21ff46642f7905aba43b19683b109be16431a62868dcbb7e6ccfabc97809d78b4110f60d3592918a6989ee835417d3e29e6185343eddb80865011a0ab5d1207a12636cd11086968c9db08d0b566f3a5e652abfb67f1ecb599e2771a18dea4bd6ebd69e924784c705660f2ffbb98b468546c0d0cbf365566a16f0fb0cb3c886e0988b7ae5644cb66bc9803caec449731df031f38e6ca78d876e48701d603a64e1825d69c12e36b59b8272ca5ec3050fa572f86c38503484359a83898741fee8eee3438a4e5f51aeb5712602f723c49eb02d22ff0fa0568f07164a3bd6fe2f19ce171e4fb3947474d50215e0b8faf8c3fd59205bb9ac3492f5f5a4866f9b6ea70043565d806d5230a947050aa7705ac9338a43ec5f1929a96fb2adec0e9a42d60400eef3d195c8399ffe90d8d288d9495c6ccfc3f2ac65990aef369a209b17b4a4c504394d120eaec458b45441697d1a6eb6366e40935ae4ae16baee6d47cfcac75ab41ba969484f6c244f618f020c72dce56ad7f8c12cab12f457fa6b6d1d4fbee016be0b94257b426566bc6951bbc963744a5eefc355cf5f6fe7b4eed2eb258824ce8a5d776f573326c9ed6f2b93227eb191c0d75ff846968222ac53607816f30b14629df73946032642a9c914a39219ead34627a0efdb83ea11e133bd7919fbec81a4373cf626882f99f652b67a747289b4b602437a6c0537bf43233003769c910e2c7fd602a86d33184e7677ed12971dd363e4c1cff3e8e75ac86f44e70a23ac442fa2149b69fdb2333afe8df2ad811c9b9eb84215ef712c4e6855884fc9205ac8be95fb7cfc86a87a04bc21694656c26b42c6cd7d3fc4d9128b33f7d6a6efee474c97507a0d71d8110e0514a66180514023863064f8a3bbd4fafd26c5a006c6446e4dad1ffb1a7fd731e2d60c634322ba4c57401091219eba0e21726f972e2d9b0c3d1c3c11155079085ad3f85b6e828393b209c99bb07607abfa7f7a268d354067bf514bdaffcd6ffbb8a5fd49b2835b556a8878820eb9abbf07a763d4cdbe215e55fc5188cd1c1252feae21aab3c9cae6b2d8766b3f560bbe2a06733f50836a4d214975b05c1dda335fd7ee2922a7abf86e18f315144c9750d4ba4f98aca36b64c5387d99dc0324ab74ada6c551dae5b6a2c43873c1dbdd205e88e209312b427e109f1d1e6163944db229c65e64216ec51193ac18cae8b72e7946e7a699aaa195dc3888d67ee34b0d6c74fedc02782247a7e6dc3876b2cba2f943b76919488b1ae51469569327be478cf0fc3e9146894c150ebd38f8425d7443a68f10a4bdf1e054e1e9fd94340bd6c0efdbc8ceb32558e2dab9147158adfae375701390435ee202cf6c6c8527cd81d1eadf435e41bc139a014e27163e185b35c079a521373fffa39050881e1e3617f70fb5c4e4ddf87f9afdc0bd32855855b3171cd7d5baf43cdf1cf5507f15d609b9f2c914dc4a5d668fcaad07fe3713073e2bddee7cc0d65b5578c5c9d340bbc494425a25bf4bebd0399b19cf94eda8e32accd5c5c502e02bb54d4a9c9ab7bc4f2d99179aee4dd6a8a87d05163c92757bef224a741ecd8f68b184248afa169f9b7c2e8914ac67454783cca825e58286a444b28225cc0dce6b5f32faf4540a262bc09e304c4ac4912de1408d6e0bc1e5d7107246a8debef2070c8e9678d00a9b228d81159c54dc92dde209114f08a760a27952d418bebacec6d7448e1cb8c77ccdbeb9d6218d35426572c6cd12c501526e49a9c828dc8aacf075e25bef6d9c8c82217f01ac5c2fc8e4fc38fee9a6acbfba9925293f561e44fc43cdb0b368125a79a158c42879119ea041eb53cf9253b2e727043cd975cc1456815793eefb2282ade746c3ee1c8642cf2f259ed1f9453d1a964bda96df28b32b72283496c41c8e815f675bbcc612bd0235419cf23145721de3a9d7bd994630865d4fc778532106a88637a6b2e18a101979d1d3d92bc9cd5afd7b8755553ff05b6ef98d4d261c79a69e392b8af12cd599bcd11a50680302b9e1bad8f0dc156ce75148eff62c74973c5e5a57517fc8e0cc24a7e2f1dad09b9e1598b93915be43d5a712466935fa9e0fda1009de6c9a996d309d62ef128bf2fefcb6b2ecd57b237152cfbdf0dcff88d9f4da7de51d6ced91729c704c2943b8811af644b8bcd4aba574da18ba616700d71b73e331851450fb70258896979c94e746582c79fbf20227ab81d91d927536b9379032ff77a9037adf15d76c9adf0f47553e4e145efc07be2882ad0a4444a6a7a64046bae8eb3508c6e32c5d7b2c9a4e0dd1407a51a505121a72f412978db77ae6472d6e33e8a19085ad45ecb6a36c1bf8175aa007b43d0700f7a901146d2f3159f0aa875cb3f410018d9603aa169a936b4d1528caf693ec42751874b0bd7b8ec7e01fbc72169571d509dba3ad0a588d8454646932c8c48a3a7a5856cc0714d1798558e98f2a8e542373c3b55c426b6c3c604a606ba70a16451220fa89087598c807da56249bcc2f4bae1ad480f289ce96cf3b5eaecdac1ddca8ad39e002139c8fc4de09689189ce31a6a192619b6b123b7470791c76a382666addd885682fdf53ed2e0c39d91ed58a5991cf1e66e91ef0e2a433ecee64eb9de9bdabcab083805abc68b92e4a1c951f73f4fbac09a9fabdbf08c437123581574c943b613c0a515428b714d50dbb1be14fdbe3fc6f77e5f799f58f17bed6ac6c95af9810ef025bd31171c06cd188c5c7dd628f2c3c95fd1e30a53043a94d703b0ca0f522804cbca55e19f56ad363cb1467e0dc1a53fa643c4e9893778c464ebe5b78ebba531a0f556b0f88b5f99ec10c682c40fdceefbb4410a8101d88029203b8a47afca019289379e53368b951dcfc2d4d7a4855f81036012530a7dbd5a62a434149ca983585422faf65eaf38840be5c8caa872a0e0436563ddd48c58c97b9d734d9fa773931e5629284ddb0a69cb068398c47acb7900e99bbd802f12a51cf0b4842993487c9b8e5eda971f00ff8a6f626c0456c054ecb6eafbb6da95f45edcede58ca78bd79a500bdf1cda922653bdea30823acb56d6d440a2f7400ee5e881e652fc36c5355c536ab26939fba8811bee3e328b07852b4189e19c444ff377b1afef3a730074083baf21e742c0644f334d5710ef87f9435f5dad116c5a7cb8bdb6ddde3a9b1b2eef2cc62bd6b727a80edc19e8f4937b8b455e6bbb1420db6c77008e184beed71e0422e6e3125921b40566b0bf4fe256590932b90cd14c81660ba8dfa1dfa4d07fd9d294910203cb02d65e01d5ee7d9683e9578e55e4877e05d91858e7f2520751659dcee51c07a819bf5e701d5cc9635c48ab1b614a5a697a3cbf6c7c5263aff0a542fa0219c071d66c30e1d91c268b43f770954c0a0988619edbb51f23be87f5c2ff2e96e1b50128b2ee5d35dccbcc0f460842e9caefb47134a31b5a11efd75f9d2cffc20bcbe8420e4d311bf445eec7dff4e8c18c5081580d6d6917d1ad0716a007d2b89a6d1f4b9a03bf596c3e81c70b4016be216fa3c83f216af5e570805a059d83339ce0b48e8571b114e563c18006c2d4ed0fdcbd7f8768fd3ef95cd0c3cb23f6057e86ed2ff548a2d8b0f30850d9c1b266753461c68ca56e461051bdfa33b70b6d330be59fa2ca8d546e1bf61430d9a8d8300569ca4cd27e1ac5d959fc96c3532e6e52f99f94d4bd23772df938274164fdfd1e7b8b835b495e2540adbd110ded78cefc3c644290a3f98031c93fd5afd4bc10391fa7fc924edc0e6181b4f82cb4c5f80b3b3ff175f8fb0900ac73d02b729dffb68c323bd8631e6563ae0d850345a9b99226b614d8c67058b2c05e726efd967ab3ed94b8d56ba809dce90366dc6a94af4f89eaed;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hed99e57f9eb98ef77e17ef86953d9f7f440ebe9da5bebbf734c594fb0c22a3c6632b4fa7c0b365ec98a6d4f1c247a3b178486690e793ca3ba5999472c837ca01440d9b63ff08234d29d22e92ec82df0e3756d93b47bae0fb2ca13a98fed4be9fbd0ed5f9222a0e7c3356b654ab08509f09a8b410fde90439ea43e1e2f2bc7d74c573ff5ea4d2a506f1e6c7a4f494cf5ed32e8cd1b4c0697fb29149fa9ecb101d25aea7c6eaf0fecab0705df0ef36df7950ee33e8dc9a30707459b41be311205d9ebbf3378cc2568e1ad07333531f31b1f023f9d812aa5a50360401e2e801c2c1e9d8bb0cd3739efd8ad0f16460ee918c5bd7aebe5ca0b743446c8e1f71d81227a5df249537604d5ff44922addb9080cb1ab709afbce54643e9060c5bba0f7dc0e9c6dfb752f4b5f363a00e46a4aa01c755f230be4607724c46fe1d3fc93cb57b99a18dd4ea143bcac7313c40dfb5e376bbe93dde1ec4ff46557071724e284e12c8cd65cbdd1f487cdc3ebeff6b88ba965bf7b0043f8beccde74cf97bdb93beba9bb536a1dea410074815d91d31aff9d65755e4bb7e4161f68e3c61d1403dab569d4d3f2b8e4c6a4a29fcc83e96e601d7d3df84663e533c3f4fd4a7904a8d84fc8be7433edb8c373a46cd9e314ba89c13020fdc75ff6253d5d2756ca2e2bf0b46124b82dcf55dc95584116a7bb7192a317ae5a6748e05bbf4911c9ee5e3de75be55761568a5b6346faf9247bf04efba3fe77dd0050a24b2a4020b4d79024825dc05823f765e5d24adcdeb4f59b63920890b9dfa4591c5a5b555810b7a19eb5c433e06c8ae08de7af61aae9f52ea4b168d3ac1056d62343a184f94d8aabce6642fcd651fdf369aca460b1cb28af7ad9487854a2c18929fc202243127a7608e0485d231f7fbf059d1e31dd3f20b59dcab9385227b36f451a5bf751c811dd0db9ff412d829ce3250d67e42acc859acb31452317e94a5af1680c90c6d67d6d8d5a78ab83185ef35f9739026795d49e73664f0111921d37ac48d26e3554751002de62a9e7bd8a84d2750708ec67924969b8b5334a04f075d34b341c320f8d1b7a71258799da2ab5197b8cc0f3b6220690a62edd03042c8c8d349feed2e2cf0d1b33f546fc89da8b7b96fa696c5de0debb18cadf24dbe3432b3d05078b9fe2e0adfa72e20d983088a457b5d11183ba980fe2ee959bb45d1719e36f44a2dc6f211f6c94957adcbe8b0aef534f9f8e60adaa799818b1fe5664064e55bbcd950a0d3ce8130bd74d369a74dcc366b1b383fd37fad275489ac6e70253d4962da117c500e186d2e329c4c2160a5e95c9b690fb6c77eed727712a825e8cbddadc43722efdd7db2305d085c9d2baffc8cab7c4c24e224ac8f5a868cb0e5766867f1fd4784fa53ef086b27482a7266e01b8af98c00d1f25e1c2735280b790779a4e87b86c7c8925d958096e99ce33fedc885ade4c30fa87b78a53064b9fe4f086908b77dbcdd68ac6357610dfaa80cb953dbab669136dc36160c7832f9de0fe19af865c3c52a14170c0dc4b32a5552126a2b604e2e6b3388bed521a0e49f1979de59cb4e6e68b4aaacfa897081441edb2f99760893bc6b3130b51b6db03590a9bdd52a93eaf039698d943ad31d377846634eedc1941d041f207b145f6abc443a1ecd3c9ba743519c53a4a1762b572b22d619df7bb0cbb4380a3c316ce89a4bbc36855167367b1aa807932b4326738b8d6434340b77f9d1623e7deb3376b553fbceac6e9cd1e4a23ac92f610240e7f0bf3a3b2e3649c1fbdfe885f32820b84cacdd2be4693a1b82585349562b7ab83b3ee3361401bf1705e4f61d7149cc71de733a6473702a970a1076aedee12609a858dd983d239bf13482da68689dea72a7b76ea4d652ff6a1d8bb98586eb676dda9dd1269a8f723df4c20fea6261dafd6b9ff996cfac659846440ed35a2d73af9068a29c12fea307d1567e9b63c8d0721fd68f0d30251400b10224a39fb38192683c293e4f09dbbe61873dc87114fe6cfcaba460cb21be91b1101ba0c1306f25e3b9176c743d12733b23f7947e8a6d5598abc4d30a907476a6ccab26982e3081df6d0e12eff6cd1e586b5bde04189d3a1183365d080ae1b2c3aa7889870fe033b76a73818f270d6f586cc383fab5076370538bab7049fad90c0ebb072c8fb3c1300daf8215946966cc3108d71936589ba973cbb7b91169fc496f2c3720fc13b4c1368183c478eb3a1b4a751c1a322c594c2af4484e8409df083babd2d4839f5b6a73a3b3292b496775f8da16f37092c485557d6ca45ad45dcef01e1af8c7743e003b47c8c52e665f3986266ddb32019df1d369955fc12add1991b06578c1394a8f865e4a911c7db91510176e810f7b8820257eeb0cb12d1f0a9b0d45a998d8a4ed77db3ecdb1ef50b6321b11fd2abcc081d6624727df9da4f2f63e1ebac548c23601fae731da9d993821aeed9ce3c3320ccb95e6349488a78a70b5ac6b3778ad01e16175f23dc96f06aa09cfddabc2ddf7d4e4481d3cade4e85de8944cf8b62cae83b9111af3907ff9c77f13da8ff703fec62ca7d7d688d17995c9e56e1099c01afc2948dd42c326d1583edeb2d9e8dc2b587b7d99753b52cef1794d2824c50994953bd7a1a0dd327609e0611cdcc648328fa0cb988495e2204d13b8f87f36dc96adde6d68efe17d1d9dcda48c4f19be3f77038adfb93820ac1bf77440ef8bc6dd0a97cc7a800355467681ca6cfe86ce087667e1185429ab538909245359d0f6be16dfd77fb630b2c8d4b276d7919d49bb67c4a721d3dd065d5ba78555ebf40fd331f0fa9c2bd624774ac1d93a1280698dc603144d872e1090d38d2138646a5dcb1f2d718e69aa742980439a1e0efe046deeea50fcef25297f61fddd454eaf8db8f3bd38b71f9cf958605a2e2f4e3ffae3d13db2c390d64145e91dd14c6d210f715e92da53ec092f5eefdd1db967d33c697ed822114740ceb39af237eddbc36822d38bd619d2b41c9d7e350547442d65a073820a742d4cdaf7b06db7e32971f32996507eeed0b003eef93e64bbe22f94f5814a0af6cb9d75027c96bfff79b8becb7c23e5477f4890b9e70a341607ac25c13d0ef6ed1a7b55dd641fecdd3f98eee7e7c10dae1e1fdf590bc68aba2e40b3522d47208f9047fba1c3a5e4dedf28dbb1f741e3c3490bdc9412376cb709d423ccfb225eacf7134ed21e058bfe36bdb8204ed9dbf9d7939211be8d0def9e02237cff81a7dc7856e8d2642c0649a7155b2584a1b6a72390fc72aac7591ffd87f97b450f62bdc43e84db3ea33d91a877ba45bbf31bac5ef378c8ea8f6153a93ffae76d7974d45b129a0ec39ea96ef7610d7891ee48c41c954149a85846b53910c58a14f1e95870d97b1e219999e3945c93e3f6e02d02f076c569e350ceea0b894335a56d48d8a6b9a9b85029b67408d64a7da0da207872f4574581adfbb5e5c5f56f678fbd0bb1264399d5cd4dfb9856cbb6392234e82431f1bb1ff34b11369b32e04e8719dda05b18f88546a0a08245401344b306d2a7c2d6e4c7b3407e60f7e0ae0e9d029a1cef5c82347defba0307329a329191c982372b50d6595e0aed88f588eb06f4467a8cab9c437c553dbf0ac8cc5db5915edc00b3f7526f9213f8f2492c19f82fe19038eecf1a62ac228468694656b9d77d258e04592bb63a9588ee939fea688edf0c731568237ea6c3c56fc8e7b5292cf4c3e853c497957f2ee3c95d365ff758f5bb18911a1aca4b029db412d771efd25e75ccc6bc2d457d729349677bccf02f42a2e6ac882ff467825c61e18958cbc32b2df3f6093d8ad56b5c7c8b7062661cdb4b96dd18ff3f9ef736f409f078d5b3fc4f1261e9251a324f25d2597f09fecf0a3504eea24e5a206d8539f4a6a8687d83116cd2bfa8c907ea8bbf7a69048953eb2863c5487aab4d260834f790c7f8031ec4b462b871088199e7c0cf3c90758418165cc4f971a035804a84b11f0ac7c8e9b99a9dcf69c3e9dd07ce90f1667f42c59079afb1c55ae42b4f7a0bf6669f4371ec228d9cfe38f79f109f81d59017dabd409f0fd98b5442a3d0cd89ef1e32c74c19482baabc0210314e970b624b24777325262a1f07df42c26c9456f1407e82be18246bec9a7d2d888889c46f37a8ea42081e4cfd9427fe8b7b4923158ddcff9acd08d8b60c1046ffb89bbd37974f16b0a5d8c7f3113f8177b90b81919984ec9819d75067cb3c46f8cd762302fd524e8f0c65ef0dd2b4cc8bfb6af0cc7918d20dcfa655ce5a1f0bfa3b4da773fed4b757ef0e7e29cd886213b2d1d592cf767253dab54458360583a7352587404efdeefbfe2bc7d1f7a3d9b5b9255d67be7b0ecf4664496224c447fee030862df2a55fc9f51857bb6465e63392564a378c4b14cd4809108fa0787cdf5b1cc2311df1ddc8418893f0882c3b146327deb7a3b7be595efa0525cf0d145ce25190a6664ffa564a1fdce60fbd138ffb25469fdefefe4eee21b6fc12fc526ee20ea75a6ae88162d06b1ca3502fd68551bdcd76153c8dfbda912889bd888a290f67010f32b83632f701687e072c85b880dba0a238bced289943d158f581d311dc52bfada72165c1a677c8a104420eb9f8141971c6e0a24fe1478184c3de187593ed26a090a3698ad76dcbd719a623f8c4caf7a19bda73af034c2de668db745fa1837319be251fa632aa59fbe587756cf5ccbfbf6d5faa921d715b099a8f69d257c224f77de822242178405ae772a33135acdc8698d58d21eeeed550ac78c8611fcf915059fa482f69bb2a8512f765b596938f9c1d36c1672c98aae9e307285298ef1213c9e393f418843b7f3ea00531ac421fef1842334b6011f8ebccce88691182abd3232635cb2c5c33f4037db33509c35c73a0bc5537517c38d742239f856799499b821e6d1e43369bff1458a3ea9ca32fd6a6cbe5ba88de1d25e3691d99ff150cff5ff8d67c9eb191ecb1ebda4bc5255406c7732a5d705736509192f1c4e0f56f00600afba69c3eff55ffd8733fa335846b2ba693f9278d8e2735fb095ee99fe2d575494e33d0d495cc42407db54b6c3aceac4f3dcafd9d8d4f6662e97fcce28b51904982c7ebe848c82612de067382de7e345919248de43173489baed1c2f7a7e205db26e253cd55751764685e866953f2bcb89c76fcc20cd0f3b335ecc63f043aab657415f0dbe95f0d6133146335632b418480fd388c0c2a847a279790c3e7857490598ea63711e278a41aca3d19ab223235258e2fcb40188487c43c4755b5fec4e71c68dfa4aed9586669aaf278f01816cb90cb28c52ea20857bc1ad5dcb9485c970698e33bcde687dc664fac7d6f6aab09d50979d54bd02d939060b21346aea8896df70a8652cb6a4fc3764f1df1b4e7b542748eb7baa8081fc0dbea3823bb6f4c73915d9a48b1cdd72256e05dde089cc7b96326063f3d23907a73649af5b26f68b25b391c83feb556adac85c783f4af8cf1c9a2ad208f3b7a94a4fc009c564fd1a769e2c4e1bb24cd976f1166e13c5183c9829b86350dfee4501eba313e7305971c119f292be681a2aeda3b81fde3144b00a3206bf5e1fa648ccc76d849916cf3410cfc8c0504be8ed9416f795c09f959f82a32768d9b90d9f96b0008332b13c6f30a475dd455987d23c4667ed32551d2dd46b029ce592c1d57911b04b5469dd723ecde4b8e3dd6b7d028aa5a27dfc75376b9a2f67b691254310323fbfdfe02af7d752c48cbb91681514b2add4ce8e60e015a44d59cb6996d6286e6932245cc6d89d9b71a1fb01f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6861014edfa4f888e8d1d4e35a0fb575b93f67ecc18f8c1efce7e01493dc27b4f8d384cf1b25e5dbd2467d2cd926abc761ffe588668654c65027cf1160a2817b79d8ea2d64de19dfd3bb7b26310cae2001fd15fb626fa001c6a052fe736d170b15ab280335cd36cc4fd0bb0ee325895d497ec25b31f3b240a5deb9ee1c6ee3edb632021c5fe6d6bb119b5305bd765a5abdb946bd547e6a0d80fb20c0d41f8e9df27a9c9493344b5575ef3ed8a8146ad011e53dcb555d8ac635fdd4bbdd8b9e28ae8342230904882955f7b9b6682edf4869d2df02bb985fafb1d938ab37c1a32f210c6959f0eeb858db62909ecad3c43c33687e6714865e0d0042c1ddf9f0be221a57120b7b737cf6b4f9b125ba2a5b5178fa8bb628395387582b4d135bdda05306665cd06201b37891406519935c10e46764cdd234bbe57715a05ffd01afdf06e1cd23d8c6edb1d49a1a1c686ced72b0ffd8460910a6e44d5b4277cec6007b1fc87c8043b428aec44cc61f96f713a5ccc8841797c0ebc3b9befa2e17753f2fed16e46fb4545837471611f381d807f1c78608d570f381304ce85b7ea4818d6324c416202de93e677649f2dc93db7508cd5c48287f8f85ec63505a83c919d3ef2fee64b7fbcba9a097b6ff2d23b7794f2e386e2693e4a6e382dab44a4f5ca5779524c1ad52b08c87a848f3f37c7fff69a90636b2ccc3dc89020697fc1aa12bd2785f91c28d08e9bfb2a703d841b2921a7a81ddad22ffc0b0daa7d5dccdf17e61cbc325875acd82bf7986bd90d881161dcc1f544c05dff0220066222cdbe5c7c6395d29e191508e91795361509d098ad1141941dc6d6bfb1e5a7c4a719ac56a6123ba0338e4f33b75b64bda5dc8a8f1d7f85ca771c6d179c3f57bc68a3216cb2196734fee48151788d1dcf3a3297375aa5ee867b04fb06f877c60fe6d9f438708e6d97a23a640f8179bca8912dcdb392e65125649fb66c98d19e7ebbcf74d48b4de6429e6db1e7399516fb83cf4e51980e10ee5c1d60b39bacefcb1202d82dc955fb9b34f570734c9bd7a6decbdfd5d750de32fad33794af2e8d595935d622f077426db8d6c42a2099efe94a940c46921be75bb2de3fcf0dbcf16903feed869527627449c55577d072ebdb9ce0946faa03b3da78a9ca093fbf1750bcfb9587c23716a72d37979d7b4995be63838d470157ebf812fc349c3bcf723fa31486e2b887abd003abe26d9f9bf2a565b035c00c12936787d9e9b83d86a97de93477e699259b730a51acb717dcbc665e3b707c62511ecd3b6fe83fa5b444005a59e2d507bd225383ac60fc95794b97f09b8f6b03d7a2641c026a89a132a5651340fbe0d9fc95e91b28e197edc03abaab1c84169ce9e82afbea316dadc9db052eeb8e0406d241cb60aae9f16331ebc22b274ac988935895e57b74445f363602ec91f8928cabb1fa428baa628a7ed80ec1c3d372205956df658a8f865bf0cd8bfc0c7e5b531c1a9931d59b760e60dda8c38e296a715d32806d57b9630f22b7ca370085c111593cc4a113f7ac51f3966bf464efa3860995ef8e7be69406cc869d2c396e8a493563ee70e23868dc528e77c9a30fa2cdf42141f54003b853fbfcb383827281fbdc4581b5728b94608b7dacc51faf1633e0c2e4ecb8c7dbb9ecece22aac1ae6cb02f942813b56adeca6b9bd0fc687726b072ce71f1b3627eeb634d8ff34057bde7ba97bde26d4ae54dd4b42db673c980b73e16c85da49d580e9ac6b4df71c0ab88787fa0bcf22f8264362622f05d2247f05bf0e2c45af80b3f22ef0aa31dcbd70b2bdf798e17574f745a805caa28c5606904bac5710ded6cbf5186148bcf0ddd6408c69ba7cbb047daa934cdea5b0597b7ab439e7e23bd5752de8558c67014824426a409d43430cd2efb9e5836ae482497dc6623b2125e4738315655df9340b6d70f3eb383adec0be8d259af0e09fc793dce1c5f41b5eb4f3a9e0c8f46270e495bcaf92b8d620bddfa2dbccf8fa868d5ca164d2c144d471abb73bdf64830f84b1d99f6aee24a7e9171865c8a1c28ed3a4d84c694791900a0b693d1db8d9c053d1203d16fb796d697fff3f9985c197430bf9479c4eca3299367b98836e350a0968b7a1b36139b0afefe633b6b1d7527204618f297270d95cebefaffac3ae74f898bf5f9fcebdb48ac4c1f8a92af8c0f6e99ef3bbe1bfdd99dd16b830dac3038fc2a49f7dfbb39afe0211839f00f7773352633d374694b234a8c5d7da6fd16dbfac9221918090e8a0e1b2fb0a50fa7531a88b0939134af6d8d66cb5ee028daf97db3ebd9a142331c2c7aaecbce24e1e310f8666c8ce26476fcf274bc4a1ee885e7c0e2fba2be80ea26e2557df0b78d03f31d509efe01e52e9e35b1c9342e5944195e52e57f4437750cbec02773bd857b6e688d9b3077c029219bac294925f10eb138bb5735b70515ad60045e4db4184b9b2e23a894adc29d3cd7ec23916e2308e85c7b0e2083657dbb3d7295b3d56d67af91f78a0098176ecd075fc8ed917b6e7b4ba482983f59b96d4b10bd585d99aa46c9e9c5ca0708b71f0444ad61c28871ac4b88bf9ef971709ce5c38531155700461fd5a42486c1ed04141b3e7d02773d64c3598a1e30208614fe2ea2f4ca8ea8f068f99b42bd7678620482737c586bbde3c9e0dd96a46a006304bb6ddb69f560a7f7244f728a063cb681a9ec798a2fa1c586a2fc69ea94401c6ccb16e370ae58ac18755965a686a9347a669df984e84522918b73f442f0daac3fc4ad1dcfa7a741f90cdb0ca470394f9666aee83fb6648d08991dfc75b0d047fe7f4bf7a9217ba6ec5534ad5a9457aa51bc6003d222b557fe6598870d90e891d7513682092c6fb3496b4bb8edf004214ad2fd930dc4ada7a296395e8ec8c936b669243856097a07e77d054a0d871b41e1646c4516f5c5f6f92f2ac94b3177f1a90886717fb0c7dbcc90e30a9d68259ad6222b8801ea8709dc58d8708010f66aaa983191156892e75cbe18123d345f927a6b17fe7170f21ec6a7760f809454fdb3c5ab9748a3104c4d1f71fd18939d7bdf2ae265edb7364da46463b0171fd0d6e1e58103a1538027cd3ee93bc80b95f3559d3647e53f3acc1c1bbcd1336323dc8801231beadbb7d1510dc7b97d8b22071e69b44dd4c5be26aa738ec7f33c2477323be9a4fa50b57a99cff3bdcbc17320ad0a9c93dd713fc11e87091714d3e35903278e855e6323666c9786c3288a684faa746d9ff572fed8f617d5267c601a20cdc55d2e1b1f815a8f45e553392f14b9521581cda83cd96da3b87a6c68b5831aab599badd31f80c3b1414dcde48a70cf0264407ac6aa2cbc0ba2d8aa5064585043515ecd2df34e940d9838f578c411e6f1112f380a9e0b6aa81c56c2fae0a0d9eed15c9221ac1d1d81d5d7e4a8b2870313f78042055182eb51f50ec74043e721701d7367275658bdbc5ec69a1d2c135b9b858aa8a5e707af23773157bb86a1c98c69371bdb6fa03e7b02c61dac4916a6251679adfa74a5cf878de86094cf27dfca2d66dcdce4d93ee5054a0c1f7a0593dc733ec5856be17be5851a1f90dce108e8a1edecb1c3b33c8eb5bb3454c5bb450f4a5477836dfd6b12773310b2969a0568472712835a2c8d59d1a6acb90b0f84e5fb63879d38feda38d0974b017f5cd169b66536584d9aeb45430296aa6876f6da414f55523508d804ace7b32fc26c1ca679e90d561c7d01452c19443d0f29e937ad07dd3141765c2e6427e0e92f506c9f00823d6d7663bfacb661b0b886203df0164124b50cd042cbb93f9493b4294a0e66b1db5727cab3002c144cb7b5d9cb845f886e087b37d35fd37010b55efe970914f69447749af5d6410928344e1d04010403683ee729c58ef64d9be60c0fa9608f0d6748fcad240f317e44f3fd64cc2c2b8922c2b9b9445ea6d742b57e702a2bf28c44f822616f6df4cde637cffbc2cd812bd0135f69b83516719755971731629b1625d827ff7b95055312e838a77f9fdd719c53e0ba934a1a774f211969fb61e21af05412bb591d15329db12074bd9e7cf5dc365e595fc0676465e8512af306b1d3b904e58ac06f38d652220587e02c7e2b9c8a2be392f63be51b44afde6b31d3261989eace6e244d8b9f941d176e9fe651e507bf4b0232ae4ef60373ddaf32818bcce20c1e3c11c8e2875ce6edfe3408558d5d4d5847e9f43cb81f6f8b620ad15fd223d151e43858743251b650b79cf4ab44b602417533da59f5e961f722bb2181bdf35a1a4781ac2502e357a16067fea4b21e913ba355dbb84ee54a4362d7c1efbab33b4bce3bcbe05cc66632df73bd4acef8ceaab441aa2a1b0e85996f8ef9d451d9d041cc8036bf7f9da9fb694af39e507238c5a15192df4842f383efba95ff8706f05ed271d69543895dc357d63b15683cd0defccd608b0191ccd6c7299054c011518e535f55893f338f2c08b582cf456adaf65f0209742d797e58332e6f96e863016c9caf5041d627a04a6f4ad9d56a5c4d44239655dc64cb87f4383aebf690123d684dbd374a5c3232ae1a4ece7bbcc008beeb75882482d84ea6fa7b64f91e69071c360c4aea11523300b57ef609220547d5537539a0675dd227f72b1b73eeb59bf74bf8732b66417df5022440a6b538c7537701f89f16d93fba25af1de1d6452a17acf93cb3f057c6bfdeb34d1d00289972f7d67c642cc89c1814bbd26ef1d464d284eae4a1ec1e2e48cc8f675577c02dc5be8b3997fc2a420f7ce3aad462364b12687e6ffbc70d1bed1e842333bc99e4fbd243a8e22d40425659cb4d5cfcdecdc3c44eb070060dcb8f4f2336d1bdc746e0634b1207523f9b0fdd489e11374722fafbe440ee4124543358a3a5e03e65fd6e79bf4043910a03cfcd8883d57b71be040f03303c98bbef02a90735bbd0521b10fa28b0eafac22e5d24c8b939900aa185024735acd7dfde8ceac39981a61b354cfcd825a7b2ec1d3d187e1cdb092ad57eab8b072a3bac3f90d1d83a15def6fcb7018302e16d8b84f69361cdf61f64f9f4a4033b9bf1042c7ee31fa57c33a61bf3098ce0e75626bb70b81840e5e3a09352990154b0063f5338d7178917bb2d087ed3431cab0d6f7b251b682cd0a37bfaaf3d623f16472713ae621c11f3d84eec3d4bac77b9bac9892c87735af05893f7331bb6ce4527328ed4a934439f9457c6003bce3da639d271b6dcfe8636eb73dc0ef32ec512187fe7226e47d9ae0247213651731fc2f14294c389ae8d224dba31649f6f4bc85500a38837f3d3469ed69cfe0c9abc14678afff5857c304697c9ff908e9609bb1703703c321e128da27860c15100bb00028c0a59965aca307d9ffb25e1e043d210beac85eccc03783c155906a544815701397a5d021753c5acb7dad44fd9eec8576a98514bacd3bfc3960fa63499c3df101d1b938f9f96724a63928f393f14999266085f4ce4af43578515fba246e4223834c80d31d246a329b0c12fd996f0dbc2c438cc70859db3968cfd269fe9c2c7ade128846e0d484e8ba8691b43421a6137ba7b94bf2e8b925773ea0dce0e5355901e400f42f0eb53184da832374e7daa7299e4950ab48eb1cc766b40b3db4dcb88032e0d6bbef5563d9a1ff51c9d6f757f11c49533f32b479f69c87557fadd3396dc4a925b9c346024dc2b6b5aac18c02a186eba758dbd9fe1f849ff91f25d41424f2ceb1ce531dbf3969c20af8ea54aad8b062da4b2b98196fd491705edc6e5b13db1182b96f083129f15fcbcd26d302800ba37026f0b69550758935b9e53;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha71ee0f1bf192d1b7093a4b2bb18477b0b22acaceeb31cbe957c4eec1657ff8384d53ee839f9ccfa9ebc82da3bc4faed5fe6e81af568c18bc478789264513fdb5c84467861866ed9c702f205b9a47f1527fecc940573b0c8098b393780f9a3320a8a913d34b76ab55d32975bea43df605f191c5380499305bc027eca3037085643c28cee3c8f9f97bb9b239e7428ecf2118e150af455fc8fff23edb1ed4ae9cd9043da8089272fd90cf133483748e99f15d0df69e57441cb60b647b9f8ffd8da7ffd623dd805395caf1b0866e2e874267c23e967c4def04b05baa260dda54fe2e7fd8c19d2af6a62923d001d3175240e8a36fb805ff6596891d27154a2649af457561bf26cf3c5bc026e019e63d9aa25c30066b9172d83934c9a542ae1e2aa9093efc39060aa7c9ec3fda8c26f39bf78bf340d1eed42e5f60481747fb7b95cf92d76778f08cc26141e85499b2602dadffe1937caaf62ee52f08b3eb969a35ec41c31bdf604b418f081442f92153628dc4c3225d70ccf6b20df3b84899e55913e6c14038a5509cc6f3c0f333af0a69927c28cfefec106ff672b52b04bffdb37fdbf8233cb542dfb7b4e6792e6ecf6cecd29b26a254ba5ea3ab786ac1a8b44e55657a7411f0dd2bbc87b74168de54e54bd75b0c73c8c3ba42b30baee2249479d0a01a4c74afefac4e41d349ce8f8b4c0a1af9629ecfc14bfc1a47d4960de4de8edc6790b47f7fe83a4d5dbb555dbfd6d50b6d3c7b9eb7eca3d70336a3398bd3df62f18193d6aa4c07e69a2e2efd59fa10afa6d70557aaf2c523e7c3acf7fa2192c8c6a42e5abadd235f4248f0be144c3ec21de0399b8f629010039ddc65cccf877eaa57fa5203900c99d4202d2d49c75f7aa17c55c19a18f0831c790e534c0d622d7e0f017bbd458b12884d4c0c60a7097cc81237207be054431d48de45402fc7b0d49a24f4be7a18db38db96ecbaf2d4a98950cf1ae9c5b605b64beda4657878300f51c4fed76f72d962942482cd160883c6c12410b6e045c55c301bd50789cccebad2b4869479d144c5f57469d752dea53be98983ddb866b7153e4f5b3b797a439d358ddd8384169961cbbf2d7a7107d35f777e0df33f7f2df145ed957b1be61740f62b0bd83bac9d183bdd9a664d4a7a179ae8e08d1ed02def72e542b4656101d64508e833ba53c1047503da20efd5ac4812aade2f341ed92224516333b01e0d600cc675bcde46d0e40c14f0b0d8b0fe5aa5da27f11bbba44e2e2b01e68184e6b8ee5b4cef17831e8c0f29adbab607e27aef40cd0bf77b0d6b71fb0a2daeda40f49b4b38cbcb4deee71e2c97d300b8dd9abc046c90cae73611d26ae09f8375db1a36823cd1ac50164c6485aba0e517922097a7b3b9fc61943ffd1eeaf0dec9fffb5d1a2ecf13bbc1b2235dd5f5b894c8542ece3a0381e97d525250855426254aba868599a27cd987ec58e4a7e42f6aa7e009b392e0c54ad8b0475787817d508644fa821b95e8d263e4aec61e364c279a461ade53bbac3b0b899cdcf0a44cfda0b7da258934730fe6262dfae19915aa801c9d2ceafb1664ad06f04045ee3e3a74da11ba83548b86bcd218f4e2e9894380f3b9aee945df95bca59d806700210d48fd56e9e264603a8949bfa44ad43b2cee2823bc2306e31deacabfddad79534c89320c1c3ecfcc836f1e2c308664db279b6309584718d0a8afbef0f4b7bb33e3bdb45d4c5d970c5463e2cddbe07b3c74ce3b30e365b72978cf5e85f6717465deabac0f6eb03a883babbc351f8e172a7bcec84c70b8473bb9ef2d30604b33ab93f6fd86a2d96bd4ef32445488dfee1fc19a0b512d5767c0cb8f5400f54fa6ac7066ade509a2834ae5552954da444ab02817a84508fea74dafff7b4f14e0e3166969cee150b2edeb5c074d322198619d47ea24a84f08fa480e20a8e058e021d59523e363c4d375e28cd24592d43a9e75e20d47c27c4b481bbfb63ec202fc15574aa1870283be416a02f9f62ce557cbb6f597e07df687104fd45c8d695a4db4cf126bcb75a1ffb19f595255508150409c44a0380233ada3227a8e420f41ad1207c74707a3cc235d2cea45ab7745e600a96e6f029dfcb7fa1be45192f295804fe9a518f539635ab875805ff7907f93fae7b731707334262f5fa9ea298d5546cc1931eb878406e30114f344c6f8f681d1c1f476888701770d98d238a15def41e1e30a8a22bf3db42f917b7418539000abe83084fbf3bc9d2553333814f932ed90713514a113f2c8be05259096703e5a8a1d34d354682d1b6c19553bb22a41a9dbc4369ab3a2cd1e15fa202197790e44ab4e86df0d9487c556d908ddf735a8264a38f8134b1a5943556b21803730b091294c5e381a60f9424344a62cc4f5c5f880fd564d25fb89e69131e3f1ef2c7fe7ec7277c304d7bef80318a07a4f5635bb65c11992e8746ad8faa25c09fceddb9460f9da1cb776f96e1dcfbfdf737bb6b7eb0a8fec501938150528c7bfb2617f2977466b760d93f61b432c2e4f2d6a43b7f506e5a7f0540998ff43afa3ee1d20c341966f39087ce740c364165139ba63b832f18f36f18c000d718690719c5365dc62c79f624d3ebbffa5cbc17223a50591ababf24b7b654b95745e3827f083a95c8ce1ddf59fad26a897b2e1855ef91857cf56d6e5c22b9df18873f1780be059a7a17d33dec496d129bc84cd1143fbb1e90aba75099abebd446fcedeb770590422b08476e8f525717de8b7bc8f087d50ec1acd69a6523b6c888754f58c84780c1d6baee7c9765b697ea75b57afd83b6dc901a0fc80b62b187a5dbcc7927ecb67a1d45e93ed4f0a5b68c687e8cd40dfd08628d16d2adfe1f1323ea9884260bbe8f08501b1d1c7931b57b6915fc62a726a05b4d64867df4d2902188361ee32899c5613d65e599739f67548229c8f87abf6e35480aac18a87fb639cf78a2c9476d91e933e4e646945b91496926dcb730b02bd7ccf635e8f29c085973e92cc21a6562d31a106a955b62a37ec69f0d28c59c55fa2278631772fafe1c127f5fdf18a6dc420c6a33cd9f06e20fcf46130c70e8714050643735ec7448c1eea365707ae679530e4f281c2804d2ee283339465cc9502c23f89fb61a5365a5e6e32506618c6385a1004c6951a095ebc0a9b939b3a8a122cf17b5c6dd6a379e122c2b3458d3f17ffa451359b361c07b2117b794bb7ad303059b5044ef9c63967fba9177ad1b40f1e926f51556d145791138f9dd1234226f9dc7757f7f75b2afe6e31c26bcf2ff856e282a985144dfbb2c601d740b26e854ddba2d217e08233bed2dd7367f00409ece73fae0223a1f1f9a9dfe4028b098af70e9f8781d20ef4b393ed67601d222088669fe7491bb6b35d7da9e65dd160608e88f7a43a06739f0613c926c202fded4be33481dd2feb7dd3673f4342f1ffd8478c04a63278c585beac436d444e952189e85217fab07c362b14454fcf2c858e4de8f302490a6a9ee0d8fff0a061dba961f1982ab088fdeb989405d89e37ba6a96db79e8315e4b190e55b2bbc0e08c2d4d291d8b2c09c458410f893bd59c9c3527179b7928ce572f9d08dfe38c48949ce7d661f57e9fecea7d87ef2fc5a70df684507c5ca2d981a1b53c8b12d2bc2905383c09decf1bc18fcf37a04ec4bc22046d1e9ad8355df02a988aeec4879c8fd8352c8f60604215b74b5339bcd46db836964d0117221de003f6cf9f6300ae2124473c55552585d473b61875abe9b46ec43ed4b8810a69ce0720aaf447e51d3cf8a893d9c81830142636cb42cb1c83cd44951395b2b0dd0012ec5b62ff7f8c7f867670e2af944763abac5d24d8526c2c1bbb6021dbd56aa15711854e9d17c91cac246a1304abf8cc135174964a7a31b64e3144da440b549e998249f89dff53fa83499909d4e4f652636de872f4438523e6f67e049739a7e8d0802ac3ab64c660d86b946b5be78e4fad2909abcbf094b86cde9359ecb326e3621e5fcad1e504482acdb1bcbbd8045c2648951b45007a05a50ac441fd3878c8eff1cb7d79a4ea9505dc818b417959d66c0c31b878d601da437e591246dc98dd81a2b2524b6206a0ecf281d48be2bae1d9f0a594c6775d2dabb46b150f73d277329da51cdc976937a8f37997822f29de8e488cebb0d415885a65361880edd9399840facb578c5eb25408b16a97118771e8a78dd20f343604d42b90cdbdd1a86d6d16054253c5eb83535907209612f268df7d07dcc34a813cc38ca31efcfd47c912d0c6a0d922de6f73af1cede6e87c0012a6d18c2c5eb7e5bec42c46588e55923ea83ca67b3a06516903bb8f9689dfcffc3ce3ee0267b1162152b40fdce71fdb103636f14809d23fa18b6c43ed0b70897ddb222a613ad492df991aeded618090e724cd1435d6f4f9e280ab6ec4ad7cc9553e90b333c3d03de2e63db46762cd469d119383c0bbc7bb5ca61e6f03361492ca9b4dc4e87e6d8dee377a03bb7442a66ba6fa1cdd15ed6fc4f30cc4431673e9472ac6cfc4f2b969e375f54787870697dbfe253a9a52ee2057f3bd665a653d3b7092187f9c0d4e76286c11476cc743d913910ed5922f4aeeebc34c0b1189307fc6df51fb6bff5d6c568f23df1686231ad73bcdfc8738c51539efbc64af95e1539acb81261348ff2ae96dad1cbd5da43cf42a186df1c5b31a67435b23063d36601989b3932c8bb743809f0a785a855a2679371a990f8ac63d5d07e5533bb026a721ae6e748dd798d6792f23bb5e056b9159bf5ac0149f472f92605021e1b1bd20b956498544853f6554bcefaa4f836c62fa0589c816a6e589b416ea3778493c817fcc1691ae8b289c22b148fee4443e2f7197d83e691f5cd42cac36c6e7511b70da9ff018afd570c2f5028e0447862a9be20a21bf3ea14af9ef0f697e8803526cd6903498f548bb97120515f687bd350e79621c6f791c10d758cfd94be05223715c8577bbe543de3804c2df526d01aba30fa4994b0f0adce937183f362c2717bc0598e9b1ade1c9d3d0e6d55c9ae6f9377094acafb88e2dc8184e6afcd97e33b687b92f128aa2e051fe2df2ef52afb22f420a2fefaa618209ad451c50fd6a00cbd884ce043fa35c9ba9a3e4c1d1096f212dcf579fc163a3632caea76c2e03559ddacfb6ae68b5841f2e7d77ae5ea195e0362fa3638de9b8fe8479c805ebde31dd9c629d0c8abcb9dba41212519aa7de16497f223035fb591e43a31500385b47ac4a53d744e295330215d004123aa5a4bda9b588a45085b000cca8263c2a781c417cc51260ada3d05cd7427335e2b2c557218349bdd42acf03033d2f6f5e638ac7e0ef2997269e657d45b8c72837cbd2d3474e34775eb686e977a1404c960a807a23996c54720a0036797e519f831a54bc973a7c079e107300c8bcaa8a20d7196985f1591ddc9985f8f6633f225ce05fbb62e25563ec30286d9de9f48d3fa97d210ed21a80e5eddb05875a7e7e4d56fdd4ffa8cd3733db73981b24b7981c6cb7adee2b569cf538e232f3dad7055c1d8c5262f679eee97fcab447a02b266a03ef16d451842ae56cec87506bbdbca1b67d451c4343c2feadf4891329f355b87d1d57fdcfa9c390ebef5801a8d70370a2cd234441e00a58e3f31a5fed180a5e9fc8d157834583f1395e314c1a9d5660629b4453e030fafb5788b031239f8a1fa65026f7d3918a0846503d04a1cd9f96b5f56f670c4f534c10eed19abfba09af5aad8db044b7b9a04b722166e1d85ae3aa4b8907df5a853f580170056131dc34bc34754e468295669652de818c754b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc87fbe05d1163e734f57ed7c82b00af0a561c4b3d47646e3e91b5b0e8498e568e4ed871b6550f5821183c43bfb6b194bb6219f9c4621299ba81a8ff868f5538b2f88f53fee40722cf2fc58569ae4ee72965fe69babd362553f5d1554e65dab19390a9ab29856936ee3c1d40407f5d5d64ee9b896c8639dff4e793e7ff95cbd2eb6fe1ad66fee5d5201537860661b1df6480f175712a43f4416a688f92a13c069178389e16ffa2ba514250ec7ac039ce46b010c0a7e9ea7ee6035e726f76f2222475a632590a3e87efe5354278ca4e32039912401c5c0d2e02ed395db5931147f32924bcffa81117bcc20d56b5deb1edd97a47db3cec97ad8019fe8dcb6ba8a633d67cf178e168d2ffe7a2ada792390bf2e853f6e289b67a694e6d0a9c0c32938dd940ee365095ec827ae2b8872dc796faab2fabd086b20ece053145973a70b1b38bf1e8e0c09daab4dff6cbec3d567f39b015b0e12b178a58624eb3dafd069a241d17170a4c3d967ae91e27a12a8123f50e917e2ad0ae3180af856cd7ebce22cd009834dd7a85cf77b93dcd81c02ba2d5e889cc55942ae2f1290d09d32783606c703a4edae2b520301e2bc9aa4b21b71cdb41b68c78da6f4fa8cc6949d891eb62c9dd7f0d66daf9c103184960bdf63409e823de1d294e5fcb37bab4c1dbea2c674cdf16a81ccc36f6611a1bff3a4221b445439a37806025883aceec065d5c845f5395323df226fffd6ec77941c0e3d7ea12a6b136fc229ad7eba1985d958ba74dfebf3612f4ee60a7b185c9d4b005ededac9c23433194d20fe5202537ac78b911a499d566228b3641de230f7f7ddc32dfe9f627e93c2b3518cb7ed7995764a10134d61c6d7de25ae9191c84d5a48e0d20a5aa6ee7527970854e6be38a80096c28e843cebe03ed6a61e1329e86cbaaa6cc8469a3e47f42943c6df0c1c9eca91d7942a94d0ab6740d0bc470ce5440dffc983166f3460af16102a0094a85fb53cbfd43cbed3cb1ca9101e8f0c1cd8ba9e7b78e290372ae2348408244f132e6c855808bb10b661ec504db5fbefb31fda18ca07b29146c31913671dc9daa0d848d45b7436321b02277410be48006df658c8d3dd066b33fec508f60134606905fe18b20cc96c562e3b180bec49cacfca70610b2979a12ed6ca1ed5490a2e04b2648da6f4cbcf6c543620983282df878775a6da6228e3db1de155ba4386032a688643493baf615e11fe2e2f69da80774f0d5d60b39ac646de66bc87ea237a965c07d361c1b140409c20a3aa7870d3dc04046bc1eae5791f4e63cdae7f62f6cd3b333e6bea148e0ba2868cbfda83e0505c5841c63ebed0692a29434761fda35f9d62ff25fe6386fa89962db831c25b86bc88bfdaa888ca3144354b9b7712abfbb9e3fdfc9213305d68271f15aeb847d101c8c62ce8d778198b406d98f0a3eadcd76b5b5be6d62c85595dd684a672a418ff98e340c7e556d4f450be2c30a903eb13ea5f43fe283dc43e2a82976544d8a62be72e9a879ed62e7e32b43f1004e02c793d45804f6578eef877b64940612feeb27a1c0ebf021975b52fd9218a8f14d51d552aecc0a00b6176bb0ee60a5a250798fef1efc62d0425ddd80508018f2138332b7b6bb87d344e5a3ac4584a295829166c2dfc90b7946eebd6b84c683db16130f81f6074ff2fddb1c15a498968f27a9939acba3f451111786a725431bfcfa4c9371cfb49cafeddba61f3ee6cdf388c85e78524925b1b375a3fef50c1470c5524c998136ab2516814ede63d2598a9c74afbf76c73d6ba46df389834541017c4c9943317da00788f16ce810b9157508e1e22767c3d4f83bbed56b1c58427720ad98c11eae710c8def944c4149e02af42eec2596d99dbe4bdddc4324d7b5c0485ccf02488f714662be1658f4e5ba2f011ab3591022f96abb4649f70ea9d53d824795ec08e670ecc198486d2dd32297b8bf0e2635b2592ea5ed2272301e761ad7fa8da7832eb5dc8451c22d4ad76be695e1ed901767ed361c8fa860963379a99ee864fc94a86244bc0a3b366c55a4ecbf638404583e66f578308f5485138ed71f64c2739675a37b0ce2a8450c748f75ee17385a091110f3b70c88f0c21af605cc98c460d72158671bfa370d6b5fda9adf1f10e58a1abf39d317b64544e37f4297c853f565802a6b252ae57fb1955bb7a31b35ef5fe953d0bc1f9579ee0fa6becdbd21b6c7c664d034d1afe746242927362ea81ca15ca444404788fa3bb8a610d6d2fb3719ad8044e6b32b4318a847d66f24ac119e2b9cdf6d9ea3783e84c0d6a473674d277a9e26e32f191378ce9e617106fc7a7339e10a0fc0f98b26d0c59a358888526f2a34372ddeca1cfa437e7a0e300c74e47e16d643797cd0e71afd7adebefa9bb0c70cf560224ac19d8fb48b92b78a478d709c82eef54935855df47dc0af1fda6d74f344a3b8a5d7266e435d80b2dbd37c9542728b95450d9856be465ade3f4522292e95c9686f12714ce46286e5dd73ea3879775c29dd391c7b229d7bee8afe1d65f2c8a3827c3bdabc4e3f0cc455a696e724a496e540c06ee005e26128e46010ca6c81d430d7614f4b00112284b3fc8ff9db95e2ed0a115db85c619df7dc06f4823b0e1170a2addaa6a34cf450988c1a943d76552e0a1d85c77b4899167c3117bc4398dc63d1558110c6bb20aa49021b6cc28f577e36cb5cbe2ca4834d3eb73e55756debffef811265d7a291b20f3e693152fc3a147eaf6868bfe8e595f6a8fa717552f8dab76a968115a6caf5d61d10f3a45efc61699380c53944182aa1f995b923f89eb67260fccce3ecfb93193d4159781ebce8a6905989bf5bebdba8d0e66af1a3daa39ecfc97af7ad0d9b59f67de724114ccc623115d7329c8c8c33b1032a8ae2726282194d6adce880eb692846235c5412d36d2d6d5780dbd1734c7d492af657fa82b2899eacb3b5d4bda177639ffc575e23801d7d021b07ebba2be427df56704b5cdc52166f1bd44d52d78d474d8bdab7c094ea04742fad1cc77a00a2d28297fde731efee927179129b700a8c996c611006d264d4ddd8c6ed7dee18901c769f7ced47f8c58c125514555a796b8d53e1c209a65aabdf81a60447d88603726b4b9847b39f31803951df81b1bf897fcdd4122fb70dcb364f448795ad27958e1b0b6449bf348a7f03a3e1d2fbc1fd199e88ecef6010c3b537abfbca0701bf74032cad0544d20cc614e60029a5cf688dc8d542b2d6305e9666a06c50627789ac6bb526d792383e72910e7193e7698f130381c13cc2bea01cb33af7e49f0c9d37e308011af2dd5b245bfbad1d635a9da49c645ca40b9b85fbd55c6c6b17565edb3cf92d8ddfc71640304c4b3e1aba338e54aa18e367749afa47e23dba17ffd58a9895606ec508ef92099a70b0488d95652352c29dbffb42b2ee512aea4d6b0883091129f3a278f7539606c7da173b6d0b9ac54e161b7292f4688e309893824d2335254fab332115b134ebe300867457f027ca1d0d1a91aa22dcbc9847acd0986921144360dc6594f99296959aa5abb9cd691cbc59b9a9d594c688c66985b0777231b1d74b0a0ce17afe92319992a1b193245fff282abd76da13a54cec8e44ff220d813fa9378a3a1212f66b089c3e8f2657fba3d9b3e0270803fac6c2a7d66513102527c10c89859c1850d4d139da63c6d6e5e670dc88884b6c449ca9b33bad39136e7c47f7be1c60ba4240a0442d5ca620d2bd695338fc59cf02b8959fb243bb5df30533324d620ef92d5764c4b6b0b591ea929617e0da12bf2c1e2a9752e094156e580867147affced28448fd0f4cd34ba860e75e0c7a446479b47e3e0419d0bc8c718513925f57803d46acbf4160b92415af564a68472554da50e334c161320da5c65377638b504845313b15e72750b29bd9cedd3152696ecfc79b579393bad96d3f1f7a76ba06471c6bb55edcb35c47c173fe57c033ae4fffbbe027ef2f5b43a8a8c2e3c7ea08a16f600dacce7ff61fe3ee5e1b0d9893dc4da0df5a4855753993abc4066fcd0fd13a57cfef49068a691f40e0d148a41588b5c92968d93d5d83b8c65646143d29a21d0d4e7c4e9bf9ad3366dd5c01188e93c67e880105c765ad322b16394d2cbd662ee07327c427cee4cb8f33061d1caf3284802ad8f9e40c7d417d808ef03149c283a168ba133d8624571057367fd1600730dcd967179e84f09529de17c372a68fcbc07a8890e558aead7bec616801887944874fbcba53a0b588540c87cb0c5bf3ae137251cbd544b9cb2cf14a7f4bf7bee7f7562a86d2813c342f32fafcb9651df434375622b1afef9d175adffa62e309a24cd175b99ad73c76cca81463a4bb312174115cc588649804c0c0a72dbe6033e4af1e44449ff15d8b9cc3b91f9986fe9ff78caa21c65336cc7afc2dece2c6afba4059a842af522852bef6cf63c9cc7b717f8835b90fde0e57f6b9e04cbec0bd0e9a1bf2f25069f1e86ff3d7e3894734725afc54b3a4f8aa21f0aded7fa2ab29dad4b7142f4de04891d4ab81f9132541845b689ece030b172aa31b72c522f447bfc4ae7d33fc1dcf3e3a06e43dc0fb131202961e7c98b34d856efc7095a6d1f2f297e6265d94aca6412739e75b5f565b0245b16fc4f84a395c31af0c28e1f45691d322273e23ad88e5092a73a9b041b133e5c4783c943051cf5658cffaa426fc9411270e5794867b2a827b245c2ee8dc100d67640d79ff13e8393f438f449e4a5cc958f812f35da2439672c74e079675802eb6b31c2e430fb2bf7e38272797fcc845aa496298cef3ca0e1a2213d538420f9820be87b8c5752e0499e0162f8b9195bca0e2c64764e75f321c7f35cfa90f1e152c7d79409bba63f96da7d9d8c66783375d2cd8b73221be56152569a03d2dbde2c79eb57cb2dd4fe5bdaa11fff81307564bbdcdde027df6e3554073c5ebc7d9a2e3159d6a2bf7b051b2b3cf10465d51bee36f5e1025a2ca3f985bb6f0c540b96110a2bac2a45dc40a49c0c2c7937f748ef0dbc714e82e4b22db6f46f14433191d792615e207e8c418cdece9871e7586c37ca78758072518973ca50f3fd32c8ee803c0a536310aea1340c8d109692a250469fe957883703487a93a66a61135bb2e03d2a776f33ade29f43e96ef068640833012d74e485b596798be5c37d3051e9f2266759cbd0c8323096b37ca2497cb068c409ec2c25325b188d65a3aa0de558be09d0f8d144eb7becaa1e322c4bbbd564db333354899f603ecb5a791ae090597ae4716a468500d1c4521ee1412597306d955a92df9e76d861277ea6071c2e7ed4e060020cf69c04fa928a333e130cbebe55e23756aaa04115092ceb27a9f1a4821473db6681786c2ce42e76336312fd6d3edcdaa0a23770acee58c74d88773f3c40e5e9775ab910079c112584e04230df750452e1e1dc24b0e3a6b7ffe552318f40c38dc534abfa08b144f11c72aeba295a205c83ebf08886c0b4734d874c99ab9440dbd074d23ea2bac83423f57d9a6cc8db605892691b6b1d51a6213cc74b54c6064a344a34faa152ce31d04c627657b8bebb8184a8800e0a7d9b25a71b6dc6e6bbbd6c07832a6e3450ac39b1888b492fcce0d150c32bc538b996e1dec3ea594c369476c75ed79ace9a2d4df5a175756127eb9ce7e49ef11932edd2a095c15d359942950205e3ca725fafece45f42e1ad1c80a9a9321fd2ba900b9e209edda2128f25948cf5c90b5c951a08ef47666220bb68cc6a172fa1a09bdb297576ba5a8832414ce637a95819f4a6eb9727cd10cc7ae24c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4fc8b03b6aa8bd8fd3ee05c88e18d4ee8eb8788df66b7b80912beec66d3c71ad02ea9de66fb8d9842e1a839131e1ce0507b950d294bfe508de349c68fd188b398848515b84b964e7b9f7b440fa55ee4afbd0bc9139ce98ac2bef0bd52c8ac5457a8f5a015a1cf96709b9226b18b3d37c8ff01e902c0bd32b4d30f6ca6c8baac2f7ca7418738131addb4b907b1a7d84900108b4877ae0d78ac8682a8991d4b75de9f7a7835a2bdf5a6580d35c77d39cf97dca89e1057efac781dcec31286d8c4af4525376b49d946e0f8014374c6ddc46192050dc59137f56e7c887a4d0035018ee078825aebb2fb1119abfa9828895bb32b7eb1de40b6cd9ca72e047f46041c23437ec051ae89b98a8a8ff51fadefe6bf2b8c654ebbfc0b05ecdf9e56830683d7efa6fbe9ea476d5c141f4bc2aaa6b4cbea7a6e18068354e4b9481d920e9806d92db3829d118689c7b74aa84783ac846a009500c45bec4f71f77dce71c5345f33fd9429bc4d64ba1e7eaadd453838ae228248c5de508de4a9d9c4b0bb5edfb2daf91a4a59c2a28629893e2a258b4e543f81fb6453de897e6676a36faa8ef9060e071e866cc7f30a112801985d63701bea0514315be03c14477aa759d24b10a2ed3969b1077ed5aac6911b6cc1094e713db6411a38a2bdcea446d1b720fee46e0154ad09b8136eb92d85379e13a196c104fe38d60e5f8ee94498cc787e8a0e115b3a3fb166cd34bdd8433de5279372926ec8a2e01ac8dce87fc4e0a91624520b7a16bf27fd9a835f0ddc08205444f35c3133e286a372168143f264e9a89b974d111c56c2be5a2c10cf8dd74707217e096515ec096f5bb22d24f68216aaf6201a9028fc043549e335d3435b64985eae4a142414f028a8cd394231107e76d759a1f9e482cacd07d1ded675a00efea83a66e43fc3adb8cadb6b63476d60ce19ba2e9358db3c5b8dde39a205898dfa0298ce919e0364da9ce56cc95fbd38082b67d388d1b1ab4ab9811df1fa8c82fb55acf3d0d8a522ac051d2005dae64eb9cf7ebf4e2094e15658b33fec275ffbbca05fbd6102d5480216a2bc199ce7c74758b15dbdcba022bdd9d95ebc1a1510da8fcd1f1ed08a07bb241a10a024a7a2696427179d406a16c6b889f90f9a30d6c521b58c6decf66a9b4256af195368a0694984d1d8b6c9b18b008f8629d4b043c0c42a2724b56a3cf2d9690b5ce3616f5ccbe1907068d4cee016247c2a61b4620529cf2c09f39fa6c5e4b2318c4fa48f617835391f625ef3e9f88e38c6669768bb8658750bbd2b3f61d43359c27ef78248b1e2bafdd6b1e23a1369ed71192d49b2b5d2143afab0956eac8bfc480abc21e8272279b444bf1c9b041196393bba4570bdd35a46d461d0505149752453d10ef0239b01e5dc3269a4643f1fc7e5b3fc442deb3b1f2f42d3c9b492a5dd96514b4e32f24d90a252ddd2ed865535a62ce706945b899be1586bad71b6d4b62fc2f88a55566827b8df72267e0c64d264e701696befcbbe98900daaf9ac8706d4677475bb129bc29a8484db6f5860e6e318eb2077b29e24d13fdbe403a2ab9982e3dcb9ac2d021877e909b112612430ba10304016ab209577d19a58ee28a937653690b42954f2bea2ac4989bea588198ab3b39fd70dd62a5382ed7e5ab3d5e7c224a1989b9946a0f8ffd4404d840dfe38b12ec8f1cb7f015ae8e9c9efb2b42688b53b852d9b1f55defe6a39dbdb9f039e146b837fc0b04d73a7cd29bd6e21ec043e857082d3bd0895858b8106b920d2053dbb2dc74077922e6409536b9ca3c561e2571f8e68ddc129fdca3d1ccaaeeaafc31d5b1ee4c6e3fc2802ef02cc8fe0ce20cd4432577121346fa5dde943fa53cf0606e6a1131b1878b2c1de95802d737928c456dd3f26ee21319d2597f7a883a51c9039eb1956745d8caf5f05651911370bde41de976c7eab2437f0885cc8a1eabcd6424850f14a5ec2cd5eb4912c7f46688e3c233a635bcbb1596e479caec9fcf7d12fbe1974ab3daa21a33506a3a10ea4d51cbe29f5987e8ac76a03af01e20e71c173c149076a237e5a23108bb2e883e0246db08ef6c21aa793ded65da187d2fb49ae93cdd196100f698199af159430e230b64926a4ec2a55dd8ea427b9e697f922b7b2b915db19f77e4f480ddef920cc3d999fc58a8a7ec2ae86e1a98c7cc32ce340c0e3a6e9f6e333468c6ca7918a163a2d76b712dd81bf8b0b4843c21d1163afd860c2be1d054bd976ad2cb0f637eb942312323e3d966d0788038d8cea07538f552bd2a6ae8e4e8c99470bddedf181f68b1ebd469de6b4fa899698ead96ad6b9aaaec0d2faf8208e067185acd95c59823cf4c25ac5972e7d6b6d4df10432a609b7535a56c6004433bba2d51cccb8512858d7e763931cbcea94e1aa108422510d35f8f0a6922bafcbb093bd302287a76dcaae8d6f6872a266bafdc3fc39160503e5936591badd2c23d7a4c4202a285e2dba5e869dbab2074c6e0e98e67de3efe6db1efeb5c58661b249ee4341280e584564efe8c5c6bf599a06e25fff11226a34e0f1c9ae8f25e957cac5f363867fb9cfb22aa5dee830b8057db467176ffb89776c4c05265e5d5265ee811a10fd901a67a72e799d51a8e4752389b16dd2d717d7b560246c7ded83f2dee945b2abee77093a6cefbba9b615d4531ca50dadceae6ccbff1cbcf5acfdf98d5d23368e28726cdc797a3a112ee3f7630f6370d6e44a6c03e4701f32102b70bf71dad7e45a3799ad0d9c69eecc9c6f073bef3c038359b04b09e32f456eb808afb2f48167d3b125007fdcdbd5f3e082c9f25561d09af4b9289c60ed587f4b216d8e2c7827ef649263b0a3f5c133ce2de8e0f5d7e995334a6d8c41135f08ef29b9339c7f8fecc05fdeee37c408ca6513ca4b7da490e83bd166939384be53e38454d9065eb114fd8a792e1da6313ee98b4d81f20feff84985f830b90747a8a7342b69c287c616b6cb326261f8e838762d085e855e05e7ae0eefb5ebe1010d5fb50edb22edbe78a6d634da0c2f3816e3f64b82c941d09c798b778e6fed5a3bdb66e828b2e97947a7b45e5cfabb8234db3927c5ab68e60fb3dac4d3eb9bb13ab69d86881b659139d6c80818afecbf52539d39b8840a658b1fddd1162f6076bea91a3111a6cd20a9705d6306dbe68ba1193eb81e21b890415d609f4d1e6f34d59f7a41ad822bfdb671ca1fe17572040e5b10960cf8c8faa49e775c6d348b04de7eb0e7522de255b06279ef8da999b43ff2f1f1f559ac070ec5f0f3765a04cf64ea3dc1169bcb3e4a0a8505875f8321879c57007b7553107d57b690938bc9370b9c8f9386a2a4dfb3b035e77fb1c553ce677e36ebffc5260cd2ee59a8ce1df9f29ef0a1931e1329ae22d05280bdc4baefd7286d8e400c7277f156c75c48556751e3d1a2c78d3afd0424622943ed63c877b714483bb6d3f76f9ca6db14782fe72800c5513108207d097c0ddb2de73158c98240c19a25b13c20b010d2fb96ab546e108b30da6ba29c2ffdc9ba60abc825da1a3359384581fff7901b0de353b0893b619aa7a4cf4bf8b56ac7d0c47a681405503b94720ea0a029fea265bab628fe7848098845aeda80f97cbfba987dbc756628b23dd3b6688a7b81303c2c547c905489d2b54ccf6a4c0e03ec091702886a535348fc22d808c15b2b084d7276ea73a427af82a53ff52c2498910b73dd90abe2f55ee86d5fdfdca8c03c0d22eb33da6781bf9f4579159617e87169ec844667529931b534aed86d73617e8ea552a92604350ef6db6a506d326f91746efa414ccdaaf50b9001480190fb6f86f35dac7846ea0a4cf06586a57202e205048647d335cfd9cc4e0f4f0a9b52b61fd6b752631bf12fd65e2832b722a96181e9c33cb68d877d2e28951bd937146c712ef04542acf98501c360060614f703e2e7b70f0a9db9460b925ae69232e2033bb16fdd35c80352b80d41873199394cbd35e609efd12d64992367768be28b894fec8ed18b0bb00c2dca0047220c1eb331c151785b44cf0e27bea0103e00f95eb9b607c3bde16419da2e6dfc9939ce50db59ba34f0634d1f20fdc9011d97c2ec9508dd2117b68c27b75c87332fd007f41698844ef772cc0c83f738787bddab5c070cb8304ffd051423249c6c1b5e2d6c02204087c1f3feee61d74ee569671f812939cca6941f52c9a58975da1011f4e6c94241963a72144aba6a765fba3408d1bff308e0f9616ce325f7b2ae10393dbdda65bfe9ceb60644039978d05c879ad0db114bc52ffe6c72871cf5557018b33e0941f9e39d45cfa6eb94cb361b12a3cf9cf875276bf8c0df50412303352f0e7f2d6bb2337d10ca13b59e71489ec5e9c334e2377ded290983e19cd381ccb9bf76dba392073fd5dde371b43d954ab8b0d7278ca9db8e2169fdebea636ff78e49c4cd1c9e046cb8ed158fd5e3fa672d2cd2f8388ae4452f209ea65927fd49fddbc9994378c85138827bc14f1964aa0433bffa58c8cde3e4fa02e2d2b4e25a2e92853f07de2e304b2f82c44663c965af2a1a43c3d86388380553ef3ea1a07d6b9c85e6faf597ff1e9d4510903b31a4d747ad67f210133aa067cb09117d7809a895c6150ec4de105114028665e0752305a725103d024d861904767b5ff870bb4efd4cf31c17cbee9715800c90dbed38617a192428e7b1c83251ae92a9ce4cb7d78fee4bc41d33a6d1cc894fef4bbc2def2f98ce2d3e04342c0229e283f8dc4ee9855a0699b64b21b2dd317a2a13a20a759c654cef9152f568b290ca44cc160df9e05191f7e08ef51ffad66a942f4ad3f541f4d9f44964e640de4b1cacd45d1a5daf9853cfdd0f58637436e164662793570b313dc0acbb14ffcfae26538c4424536d38cfd48a37922edf8f95e3de5e38e3f696ee77e2b7674914cb1fab68cbd9dd48738f6edcf09d04dc60f5fcf727c5cc907e661f03d64279f4670ec1d322fd875b79b69a66a844c5c79d9996e67785ac3b845e60a9d2d9cf8c5321cd9af06659f76db0ef69c8acd21c4d0bfda69c761b6d9eba1c33f051bad0f0110379e1bb294e87661dda5e37f3e37fe8cc26ab9e9ece4357990a3bf7dfc67a1e7ba4a154f8538a62f8604723e130c61700f0336bfd1a64f303e190b37d7818920437c679ce6be5a58565ea92fbb679e675a56ee8a4495055bc1a6f53c15c4f307910d2732d3f65259dc1bd4b8ab9caaa93d47773891159839b2a69f1ad7b13cc5e24b78e1234cbc9d6b3d77f3ae051fdc307e631515b8232a105b996b617df115c973426b79c565d83f008a8eaea0067ac0d585731118a9ba769b4038a9c71ee52002066ebdc441ccd5454732c6a37df2faa20ac04331668752703a5a1a7ecaea4f22d0b4947c62859e6bc10c21dc3bb282e1adc83a28039502b14b666e9bd5d8c112116afa7413b335c86e689dab6da1ca16dc983f2469cbad76a78c730a74865afa1fd27b16abda5064bb5aeca303d38004a6ed6c3f8fdf2893df4da84d80f03f65c25027b692e982dea88f31a2a5b9c681f3c2ac8b3fd9ecb4fdb777e65cb6db464aef104f2c6550ae778d90796bce11c965225a4dc2e36a4240fadb13da0e473c78d6e393c901a7c73f4438430ce9a688b6cc578142af0128f16ee945b696d21dd88cd5c694f4b585007b4a0f7417cee5f8e177e296a633c8ecb6579c3f29d15462f53b6f46428890c9cb82c61a21aa841d9450cc2d971b194fd50c9a9497514625385ffff4414a451a2c54908269598da609818c6d9d4dff440680286cb633744a2ec30a29e1202e13;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1fda6718782f66ff17e2ad270d8b415938ce833c87d07605bcd200a955fa6dafcde6d7e7d167145e5f92308f822362eeb5fddce0556eaae2fee415a0c994b85ebdcd268ebfda45e15b2ac173ffedd912d9a5aeede3bdabcc4b51e553e7b6d2cbb75fe1200240b596490d74457873272586ee5c4a11a3f26ff39bd4e0705f1923e817701c469a572bfad989da5bf6fa5bb38ced5dbd2cc7367fbd5eeb1f9c6b823120c687b8fb3d5efabab0bad846b13d8ebb027e732358d4ec4d8814426490e32a673f8f022376618276d6efeea856d23236ce663cfd326e9fbb0d29f4533a8f21115f3e779efef24dab794cbdd24122e32cf3eac5df1d3a55b6f6f2e1e6cf011791124d09197ce231dba534262ddf8e6c4b6b1c5e1a7167ac0f22691a286a6d3f713f9b37012863896251222cbd604dffd141f69a522e31b8291ba74f55aa19329bfdbcee4c1476f47d8c883e0863977307db6d72130d9184fb9a95bf83942290f8159328d7937b63b28e93e227e4e56718837fe05afd85d304714620585c7e9d096dcc60d63c6b5f77bc5b9c76cfc290171947758bd9766d5291a31c0fc5688084a48f19adcf90fd4a760b727f0e5e8efbea20721c1fab4c1055a62b6fdb3548e21f5e191c71463ef95c0b69403f10b5104f30e6e0788746b1326bb3566150cfda3a1d7152d7bfd19c2800fcff28fd92d95d285f50dd9f692c1e622b2036960ff1732de93a54d6e9df19ec9ecaa9ccc42673cb946af44ccd3e6b58c902de2967cfcfedfccff9802b859eee3ee7272dd8d18c6886e4bfe6f721650c24489e29abc80196ee0d9790506353c7f852b99a23555c760efaec5e41d4e7c98ddd45a9c83c4269add85cc9a8a71ebe81275ac8c1b216e93cf6c40a1c65d7d7e039dad359ad5a680fef2d98ae113812c909bd85953b84be7539ac5c52c27dc4d99a8b032088aca0fb6ca4e29de7654afdfbb097bb215a152151d9956f8126554a1916eb6de7f669d8285d75ce2af1434fa21463b633c370b56c11f1da2ef36f21fe9fef3d1f81eed8c5b12a0f9b2697f5b62aee392668ab0f0a849af40f1a01a6de2de7dac3c33e8e30849c7d02b766b683eacd32669c0feaab47864cfda36acfed1bf4b0c6b52a85991a503148cfd9fdc3b81092558c2e6440c3755f45ee0664b1d417f65bfecc7305696f8b6353cf2c442b137dc22bc6e3cf8104d282b61c91c9feae7cdb6be89e8047e2f7a4d1f8f1abf97053f57790e507d36f7fcafee70e6372a5ea74b27bbb507f74a9d4fcb7dbafa2d3777beaab6ebddd52e55909ce358fbeb6805ecfa6fecf19b7c39984ea67260539d88033ddb85a91015b5e9733cda04f76069e3dbb2c50027f408c71cb0935a1a872484e54d520095baa29e395a1ed13ccf895e2b5e4e159be64ced7b5a54c91864f8e2f0d68282f663c9ea4eaf0b5d56b89420629988fce135d519371f8f0913b684518aab982d061606e49eeb124476aa637936a3954fd4871eefe1324dd28e8964865399600abf13c45c9522f4a80ce7b6205a69a832266ccd6388f45e40df309739526d21341ec01635f4d1fe233151d281a2c4a82cf913023053ef0ebc9a9c221c03da298a8a77e6a555dd182149e01a9ce57f9d89fc38a58ee5cf98f06719f5d4679c48c4b1276f3b8d1ea07b7339f8e28cae8684778422f43be6351e94c765175152152b556027befcf7d7ee7e420a1b6c1e2e99c0f5c54bd99dd1ae3d76c8fb51d6a900873a27801d232fa143e044ffad2421fc1ac7542fc1fb817b44f798c0f3ea4af1593dc4131878c32169002204024a835368f49e1f0a41e5e2a2d88c503ea2471ea9b4fff8349093b00535c0c2607c8092102cf49c4a05e1daaf6914df97d8e143d63cf43ff892bbbbdd0731ef66342e0e733f859a4181f8163a6a54968008310773c973ce5c59a1005433f87804bb720276e841a501fda2e3b17aeb8d8bb47237da22c05baf10bf040e5ab039cb2f6ce83e2148b02cd55b31ac4d6b63ec02ff40a48317150edff3e9464a7ef6428d26dc200f4f0982e2890873b4989d1d8e85b9b98fa1cd0fbb7eb7591dacf5839b2d6c0524f273419d44041e88ef391a21f9868bd6fb70d5089490fc79db7cb12d73275a17b0d4d94b07bdbf491df559d16af0e8f105243f9b8b71efdd92e4e14ed8a9cd28e367404a9a7811b945fd6b3d7ed58741ae6bc054e1e0cd1372e69e77b2d5704f2a68d85e451a1b22bfea9b24cb74c09d29c494032bc452fe40fb2262f4c06dbfd3a820322bd278ef28cd2266f67ea8a4b347cf652cf63f2b1de91a13d7247753b98212d9fc8b973732731321ebe9860031dfb9faf28f9af9c02680f7aa800fb287e8f6b87b8388bc793ceb74661c2ae5f6ac0ee94d9182b256f6cf98c33a3829b024b34fd99a335b348fbf6c3aa573d5cc12bdd40971ec47bbb94de9e3a6d82cdff47f08b41333f5e86bccf36586255a17982b6f4967c63696aecd98ec92babda9a7e9379593a2dce0245ef9be4348b0663876ca18c693c48fde88306b56639e359699893e3dfd476bc6f56470fb23728b7a6e1aa0c57e10287a526b7e74c06e570910106a6d5587fa8c1e1a16df7cad49a49420671716174cbf6ae93c5e0445d1547d1be91e702068f79bb84b3af15c16b95579ad4362f059ed73fdaebb1a1e8b7edd52ca27b0582aed8d8ae9d8cb91e2223777261a65b9754b713914d05598e32fd82c4bc97d858e34c1baf37b05d34ae107831df1985580b2bc76ddfa4e00a6558be641409ef51597ce0cd462312efb37cc431b545a9c4b06eede5c08ba1463085912a8b10ff1b245b6fdf2f6f56df54a2c2aeead11fb6744cdf5567726ca89ec00064b682336f52ed555ceba81f5fefd6e8edee1e9ed537ef428d5b6efc63ae17486e032c5228ac07001b95b18393b3d7828c4c0c1dafa45448329a688a0803e11d7d7dbcda73e2e1b07642e6f8d3370787661de4ed8962bca3f817654379bbebd2ed6c37d0cd477b352877dca119e5b8f1432f3b0180582db8463957a41a77bf52c9b1ebadbf7a4c0fbc005f61d1352f1efb9cde35d9c277bd6742c0e35a22eb948e5292ee952de378d46f32780e5ee0195fa8e76d8e06eb7325829813c5b4a8a82b075c46e6b03c37c3ae489385d15ac77bc04f14b4187e8947d7a7736abc4bd50c908c95c5ddbf381c699906aa34fca2901d2607a4d8568c66c236a53ee3a1909452d8433139d752741f26428419e96860b32bc0684dd696525ad0add9ade79b94469ce98e1dabae86a0dd9de7308e9531d0cc9222a48dbc9085f2b8fa2a42b4d973a4db3dab70bc5816977a49c05cd52f6711bd7791f7eab495a87f26719d20890cf7badb070bf970d06c2d59f0448a35b767e14a5da223ca68a4ccae93d23e1d05da911cfd4b566c0305687c16cb68fe9cca4729f536792e14fd315cf32f57271737a6f0c0c296197d3def2858bf06aecb7f07a1a87320d34b2cb86936c1a9e034afb5dffec4b95b3b7554a906747cf43a65b1167d1b1cf0c8c276c8b197f8645fdd31157d35df87414870014fc0e9e2afa2775f53c533fb2a15a056b9102bfbc847620f864639004a34773564ea6de5dd75478f63606971dc02b14a09dc7d3b849815bbc682160d52cfc46ed4f0743640c7d4d981cdb07cb3b06afc6c89e07ec6664d039dde9ad93a0422b49dbe84871292ebf34fe5aceb3a41958030eab98bfd6ec5e47806ab746fe0a8129af2af003ca53c6d1f9443b1f4cdb7289863790e38fd840c94dfe1fb2910c979c2aae3926aefa215b4b6d984d53d01a62aa45046689c858fbfb313daa24857ac9f7cef89190e94b689c9f19a95516a87c479d3e604d6ad847af6edd575f89baeb98dd9fd313829358239749eda11431f808930f6b17ed4c3042bd0bfb6cffdc08ffe941128bf662551d2037c79fbee38ecd64eaa871e524e68549025cd33c21de502eafd0f1c46a5be124b924c4181f2cf0c9390b3b274a6d92c1ec5b864ef225eb48d716d2814ce92d310066e7406cf13fdb3304690c98798f38b0315505da047f5f88bdadc9ed9f23cf7b48c3c21f809444261f2bdc24edc8a847cc23ccdf283ac00293b41620304786bd326a036889664873c4331c26c79408f6d4dd080647c6e5e8301b19306bbdd1b985ae78cf364df5e7d25ccbdbb4ba2798475f14dbcb0ce95c43eca60eaaab1d770d2752ea074356a2e171c1995a9070b81a92c9ae8a67ccae27c3f6dd9bc8c858ecf2efcefa9d5f5383a564e7e684402f1388ac4bc2a46fcc53e064d8ea3c328b3ef256bc2ff55ee9787520e2b50d96df7fe952b6a867364a3af6cc09b93f0ed7a96cfadf9becc1a470ad12f22e37714119e59d657af14ea9d97a0fc358ad0c8c1f67c9a91c23629258ef4c9d93a5b0c77e48905438c49d9a016747502109b982b006f73f974afabc6ca8d6cb292df4a57d70c90bc479d903c7134c637f36c07d7c1ffcde046b59fe0d29b0ff85b08cd3e765766f9276c88d68263d1b043dde416f4f889e9ab3a19f37536a7892958b26ed62a3c6d94d341d0455fd319e5b3b95865d9e4615af9f31b4c0f4fc3641064455bd3e3b7010f09beeafe7f477301c841a6f64928a9900ac52202cce661e1971e223dbf8744d127b7410c536b72b3eb4f4a60f8f45e209f2c487eb5e66648b2b6b6720802adc3424aa58642240374018f32cee5f235c3d8469c0ac63e1ee1eebd071b0ba52b65193133ef94532bf2028f805fb4049e6c7a66370c7b8201f0b7d57b395c9361f42da51004515d83eb40c5d0e91812e7e6c37a3d99a1db1a8ab3f0fe7d70f2e28329b1d01a7550d60c38ef44f56aabbf185504c6ebb029b8a8f9700524314910c1500c923343834c3135039b8ec5d443b352d5838acb40346c884767eec2d5f845f3a197489e7fe83c03796d36f9cf20420e34b0cb651924800e77754b5360c15db3d6e3ba25fd2bc86cd4583b7c0cdd379fe34bbcd2a2f40c269db2fa3a4da271606b5ca45f40d50ce220ef476d119dd91ba534d012dd2124a94ddb0bc08ed7ff25e3009986b85efcd75530108393fd2ec5e9c8ba4d76941f709828764ab55439535fc200130790e6058ad0be810a7ceb9f422c8938f5f7e0f38f4da71aac57cfbc400ceb4f4334b0e2da410a5a7e25f1f0e9c164a21cf3ff8e4bf432edc515a489a88fdb7bb6ec647d233781f6a5781d6895536582708c22d18b6fd9746b4c83dd0ff9053a5da99f49d762fd3942525da63515f62c8958e5256eb4a76137b584731d9c43e62eb594d803cb082f18c99d811fcfefed8b894a1ba3433719ea8648b2e3706ae246b1954f36a7fd560e55affd9997dc5c17e9c103db6a74d14a13fd34e4e0f53e6db82dd9392279ce503838181551d64194c056e22021c5a52d9ce4fc915f1cef755a2e5fe3c141c7be87a2f26ffacfdb4045618620a02e84c56d4104eaa1c5415c6d0eeeeb06f679fa29476e1d3c9cae798457ac4a44b286139029a41437f38b68696df9da291b3e70507fe5c553adc37852d447694245133e4ad2ab6f3df5679f01fc5a17c3c7390bff3f0a94834c9c799409659987b1bfaeb3e1025175913a438a8b4f4876f48f980a609fa78b0ac63151d80b6531731b1498452b126d2fd6147d7e85e5217b2596286105de2a568d46673c4b8096f8844be15b1cf72a89b28521e2f6412e71391b0f3b143b6ab2eb7189537a5fdee34825e0510f54a20113764b6101078e759c3c3599ba6c5c7de01c16a7ca4b8c55b6dd98dcddc5662cde;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h912ba5d70927c95f4b8a28d905e0b660a17ba2fec58d1eb80d854246bf83c97fab5694b37750486fbc4e0fed53bed5a279baff0f2bfba83dd277ff9feeae691d487d2627d109694a25cd7ea8630bbb2d33904aeb7ea00f25d4f762eef2723ec8416bc8e2e7d97d12be9784c8cce99f53b11ed8613eeeff22e24155671ae72ba4ea6850fd0e440c1e50126f3dbcc7a56ad82db32f2a265d47867ef13c0417066b5ceccf32cd8d672f033f285afe3e642f2650b97069c26cc748717993fbefce2f9bf8e04132921e8b5a1c793cd37094d931d3bc0155bf8f7a5d87f1061270ed72920ff2c09e6d4aa3eb445bd6cc11b63781efbc2a41652bf0d84bc7541d1b386532e338c4047cfe82ca139f782d38927b3188a90734a1637cd7a226f9fc308b8950b810d4a144f0536b3b0d2aa5c8ee4150af42122b8ae721c0474381a6fde34c9a5491bc095122956c4e6fbe598e600fd5d14f69cd39e6dbab1776191a18c498b45ca052a716c446f2c699233c558343f3041bb88431b0564f2cc61e036da8967946c2fe42e40f4d781d4d4bb07edfce6fda0938cc808946be4e10fd7aa73249c9861d2e090e8dbebf4be7ea535013ec5101ede155503806869c9c96e7d0175925505890504e8f3f399f89b9037d88ff4cc863d36a7b090068cb45d55b1b8e2e54c670fe3780a59fcdf8ac092741c57e716cab7b53e4cb98da137ee08c5e78a5bb0cf88c39fd16c6ea2f147b9983cb08396673267c84ee3e0d32ce27b3a21a078449c4d1e225a4eab0e6265d5c1bed0e878355582fbdea59513e6defd26a92b356fe46a994488216c3dd8783c0b0265102daac3f5779bc5ea65ae34203ba8b2e6537eab06c35d41f8c56cf00034448301724c6694203493e371e1837f94f4581eb832319c4b6607856ac1c3c493cf80203e1d09824561fde0baa01ca9d6f20fe7cfb759c04f758541818b22fe6b267994980d5297ff340219c37da87b5424fff755d5ee7d9d8d5d78b4c98c47be8a701fa78534d9fbe56bb5363c4536aa2528c95d4f784583294299a220b71f919a331f00d5abe8e6707910cf637ffa50f33f706873793785f578b075ad465d354813569f9e8513370000c4cd7ff2c1c814dd637e832d9dffa662ec220e3bd9aaa5a8443f3703e30471908319f67cec9fe124e3aa2b2f5da11b2c4fa4d0dcd28c5ac5c138cf8e320fd940a52087eb68bd516f773e387c9dadf6b3a8b2828468796a3b61b5cf72fa7f5dc8783ef636d8e6c385affd41263bca8079ca2e0a35ea05d8352088f18b9ce5d9dd729707d5f307f3a74082369f97f85fb218f281dbfb8929305cfdbdaff2b460326ca6c9abaa0d57a4e1f13aa928f262c2b6a57908cfe12e639f0a0d6c93e0a3b0767e42426a513cd9d24f7e091275afb8279926296a33ab445b3fda3c134979509999d404a7b0b72f4e942c7f9852d77bd5b3048304c029b5ba4067c9c5d58a0e1c53a37d768f87561769707c8ef39fcaac74e4ad4bebfdcaff74b3ba2422298f23bbdd99107545d918128b61cdd3569f81e4e5a3e5f44b3c7565c25727a37a1c0837ccc0e060f969dd885c0e0f311f1ecdbab91deef35e7668d12474f118a82e21ec9f168d5ff241542d11f792fad5cbab474e867b4d4f814273e345bded807d742990baebce7a4aa6901d967b32cf65bfbdbb7f3bb3fbfb31f94fa728e091e5dcffe4fac05425a4b1c3c1f1aa10b7c6b48a5e992ba8d16fc74d93ab0d08550c2cf8a68cf1d0b65699d025aa409016350c23cef0b00734e2418404aa59d702c3bb3d5d59ae39ea9db3ac047c57837d13c6a7db89fc0f49cd3b2ca4b5f896f55e97c46c113d7b83db2e75c5aa867569259897b9e0d7f1225d9402158525f5c76b7e3c742276119b4e97d843f006d99eee5f09b33d35def2d743cac0f7d750c8ab60dbeb87503d749ed5cf966f8eddb5e16246b133ff994fe94a5994ef3002ebbf48d2ac4a0bc4c12788f202aecaba87a32aa87144124a233af5a01ab1367c746846add9558c8c44169b15712b8b6c8ad9027bc87c3ee70f486caf7daf86f107564e14a2e0a6d0ad863713fa24a5fbd40329f62f494f2e39f28ad883bdde2975c03aed66b5e230da1b4cea8914e2690bfbf99d098c4fe69376863ce2d246e49ffc6b17876e02b277f452783d366625d57408a60e6648bca5bfc77e262e04866a39787b0c140aa89f421369379041444d3e136b1884d6f04eee0f771e87304f2dc5eaf84d14227b0c99d881a840b72dc92bebf146d6e07b1db42efdbdc458240d07377e734e5d0db2c1f1290490dfe1719872381366eacb06323fbfd5a482384d512631bcf2fb34d503c51210473eaab0035543484bde853a0da886d3e60f6d92d6c1a314ccd2a67c91ae855757f3cebcc003b50026df598756f1b3648b75501f563aef93909f702e94ff713516a0276c19a4f2a9d9a7d194f817390940946c064418f26b2930443e840681de15704b8ae9efdfecee51026c01167b9627e0eaf53e01f9c06382aaf879f4d0d0e5771d99c2aeeebac66fbf2b96f2ecf2701155e78d7a3b89d550bf3b38fef0acbdf525e0e1b6308534313798bfc241a7b6653c858d97b0c523a9724ea1d52ae8fc9d0d00cb51bca34f6fdfa31be82e96e842be44f59a8a9a91301e03d09468e209bae548bd027c9d663a3d3bbe7b8e89130aeb2bd497122c9d48c91d6a72d2cb9a2d9f9ef33185a6a11b8b8a2bb40d0449f159466431e1c74f244ab7adb7b99456a69c9cf5e241b3b83fd8b1ccc43c8f154a0c7637cf2c31b19054799a4a1ca8f462861a5c583e82ff96202d800a37e52e3c19a9e1551ea6630db34c01b26fb928b1006a1db743be3e77e020bd6d9834cc1c49b31bbead5e5e57c4868625dc2a088a44e24d4a62000b57983bf60ae516a3b34e98c1459a698d1a16c101e220174a7a8ba43b4fd65ea95a148eed0fd477aa0d3a3cc4f2a0b879dfcec1a0be67c1a5e9c5ef78792986dc7cbe41333df023b361d5897a5c6fcfc9f076f020a9e5c3b7d78f9dc2cf363a26513883579dd9a09f76578292b8b3ffc564bf7e164b35f40c83d1d3dc11e369a33f1c8d45be8b707c79d08d29cb704e809116942cf9fd8757019c6be6f4fe44617a194bcfdebc61715f8eec36919be9e4cfdcb96a281d2e4461035cf74170df8a254f0481fc88b37260b439a36d61b36b2250c2df4fa6102c01b32610c57b75663ae8bdfbfdf47f1273037891c2e52a241fe5d73a3950c32e57076725970fb29b71a770937efb5e6a7f57f42ec155a46aede09dba38dc38b6f5cbe809276e0c2de5131a5882c1f91cf1e36e7d0ad2396228946eb3e80385b442e28f59fddd132e74c4443073267401766edc3d12e7171e958e093474dbf3c8c1d87c41392e72660f8018690d2d1e05e6e4465321be478bb32fc506b85c09169b9128bd32584011e6c630eb77dd1b67ea1765bbc6bc0db2489692c7918858e2f3efbb8c40414a06d3920cc414bf6f6acc0fb9e3bb74f087ba237c6aff95d154fd565e62e90ef3f8c33f33e6a96b1e4eb651052183f09541662edbea7add6830262ecc3a91798bf3ea65636b247541fffdbb75fac9ddadebacd7be9d5f84c5b533927b1e6b07c436c4fd2e7cacf1f6085e1fd7071c0e66f7504643afe63a0364fe4f09e3f025eb70c8d3b036e0f5c29b73e28f888b44eab5064e9e5c36931dffa5d3867419badfdeeabb266883743d604ecaf343759ed64ba034adfc0cb67cdb20e324ac0cdfa935020da12e4db75961f97a2759c0c4cc3f2a5d4c5a62eb2843892e214c640ab3a10825285c37610142c3c8292be7f5b3b71169f9be5ee8bf9d7f07bf0101d0c8991cdab929db10c248b88dc9e8b2b844440e18323da8efe4d3fbeb86e879ccf9ac852a8bbc77c00d574612ae9daf255a40729eec06457444f7a2dcae485ee5d2dd603dc38b398ac7c946e206dfac63b788ce512363a3221a21541987a7b461be9170e1162fb67d7b8173ee3dfb26bb5d8ca2f341724d39f448bff89130867a84a98d326fa5001da783b39d1b82e960b9b0b837362cc32f0658eabde990bbf21447d2d31cf7b0dc24bd04b0799057a3b0ce8da892d949c7ee8c3c1b4594f31441d8d599dd5e9387ea7799cbf6758a71d50e5f137c3494e9b5f52e3f8b3a8254f36b5073568ad4f388f7e3d92796a769a322f7b8f6e9f4ade0470d733974ef35149ce7538a14ac5aa3f72b66aa4636733e27bdfd245f6c02433cfa397a9fce1b99df2ac65f7c5f71633b3bbcb1ef2b3df1e71f99e32d548d2d878d3983d6edd30dcffee0c2ea20ad28ed278eebb40c0a43b62b4be2d304a2b46fc33701a6b2b6d56e487e4d0849e45324a3ed9deba8eb0394cc5e42ff500f0d7a50d49b14219019a6cc13f74174b4d2c22fca34b7574922aea6270aaf38c50b60fe1ceb2523dc87bb055a108bde134171ae99941c6794a39c91569395cae1bf00ad48d4fa675fca5c1769f4845904464236734fdcbb89c6e2f54705e3366400335f2ff3a442e7a2a43a77c38aa22f408c66cb69c2cc02c77de83308ca2234e34654ec49a37f15a33eb33c26a546bdda2828772e4e7cf27254037d1ac8d5305bf9d08cf61e1236fd618d1f79c365a542be18b79bc0a25784ec0bd9aeb32f892abf1b6973a1bedb99cceb8fcecb69fbd841381eddfa6ed1d868543ba3048d49a057cdf80913f3760d0379a3d3fbd7b243103cdc25b6b071f127694a551681483b3099bdcd0f85849990a1ece36aa528faefea99404e2a230ca246a0aac9b89da2a7ef8bcd37175d0da882e15355739d108dd5511a649de7345da1d139de2c86bbf5a2019d528dba66ecb9446312a4ba6455169299b0a38275665afb1fec07692469d8cbf855dd0360184387252aefd376e24462bb0be993f7b4d35e6c386126ec427e1a37fc7e3a239c646d3be5c1c617000ba1a53552722b82b116fbdb1ee818588c47290a837f4b2b2fa622ac12b8e0a86ca90c7ddc7dc50c20fda33701333e8dad73c1fda0421815a7c7a408668ea0e27b4bd9cfbd45d330b9da53bd6df3e77dd6887271ca3e2bf53f9f0620935e03d88c3dd4af26d7dd8a24b1aa77a679d7ff5be9949758a0e5e75b12af1bc00bc1a5e86442d391f4ca4fc724d080974e2cac40489ba99cc689da92e3051af7d13a6db8e3454287ede780999f16fa469b4a63d819261a153aecfac5b84e7bce8177fab0000799594ba7b5bb2a96786e28cd21d2021f50a8a5933e9282df237e2f9223e38dee4db0bf769d17a791e7316f2bbbe6c8ad6d3021900c4b4a018e259d1c397911dda953e5694101e9a7e8c10afba9dba4738bfc892c268e42a03faaaed33c0438fa749eb595020be37a34311492082a6aa2aa8ca774ce13a5c24903a2b16aff64b75cc19910c6ac139eb58d387d66e8cc0fd056e46d26619034d919fc03ab9d44356a4e782becce77f69e8a20bfd2fb2fd2256afbcd9269738538cee5ad9371b40dc9f79db8ea1c6b4b630eacad085f4d50f01940e2cfd5ba5649e61639c0d72d47e90ff235d3500b2d46de7a0e63c371743b535d69914875c49832f5aca027239051423f13719345142320ed1858079bb4d31af429a881a85eda098d0713f677f076c8c5cbdd9f0f51b47c3d5e785aabb3988be6e727a658648e624ca68a8c63d665c8bb0aa8bf3190b159356d3fd8a95d51e373ba67a855f1bb3d6b6c6ad02907d89e767ce9d049f45f4a7330e1c08e4b57081eceb7a92605a0367d2ec1332f28f149eed523745be40cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h71b5297639eac042e7d53d3adb31d2b08cc3ad71c2a1c104e10a7ca94cebf54a550f5bbb7be31f45b0b398a33fedcb1b6850e54e177c53c78c8c57ef40a47c0c06110e23c1da9c92bcc0e577139fe5255484fae500e099b1d7c27237a930b44562442b2b2af426aaa874de8287218e09661b566b4b9f40a62b4c63f5f11f3c26f5430069ca6c13171185de1c410228aea764aeb7cc643a6f60246bc7b798fbeebe44a94f130bd49bd98478b79a924b04594ca1edb7ca77295592b48a4b8cfa28d30fa6d9f8804c4629a888776b7d658a356797240fdaea93ffa5f52a3f125eb716b813bf5808771759a9b23316f3ff2047b04dedb43362464a5fb677f3ae789049ab751d2cc2ce7f207afbc7b458c3fbcdcab3378fa864a7eef4d3db078bcaf2bf13b038bf0ff49f8df91e7590bbbea99d6afee72790dbbb247d523d600e77cf245a6fba0dc564cbf2ae9a418ade60cf6cbfc22fcad9f013d669fa0f2c7afd05e9aec70af247df8228cadf605e26c6854619425ff754943a48171e0c2bc9bd65d0d161d52daca8c59f0b1fe15eb1d4de34db1ce422c14e80669d3bd47b2b8a24d910d3943bd9f9b9335e59f7e728ae1dfb23843d75038863c7ef2258375e383e631aa69e97f301f76b322885e89e44f3ee267f2c8f8cbb9c4cce2dcb22d0bae18d6523cd620c793859b972e5ff6807cb4d6271b4c07b8e1e767e10c83c4e4ef2af8dabaaf74a344641da409ee4c7b1a3f39a669c76e24aa3426ef09a2c49ef9949cfe6db750d6b511a7e0ab36466f8a0bae7584176160391a71785ba82aad6fe3d7ba31c5d0534dbef557a57758e0cb7a8659763e14ed02198e31bda3ebc2656ef620bbbd4dcac06e8acf8f7e60adbb744e6bf5d2baf5772943e357757f0e242bae409f59b67e22bde45aa71fb377d472e27269103048ba3d5bbad8ec8abe67297c142093b6408265505f755202c95423523ac31ea915ccee8d7eb833ba0f3b277afd1f84bb69977743d720b4af788135b8d39c3cfeaf1ba3e8d853c88640d5a80b209c864c9bcec53c9925cf96c6032dbfa4cdc91d61c03c1a6b3f9c817525583a63d13369c478dda6134ffcd0035713d0b1bc617f2b656afb089163af26461d57e31b9cc2f5aa1efbbd7f9ad097db676226e522eacd72b010dfb2aa4618e2565f9ad59bd4ea13ccd0f7cba9a20cc0d652a37239c98cceeb23d9fd43b2207a65b6243908aa4a960038cbca4ea73ea1123d0507eb21aa6c184821ca671435d725ae01467d8048e2c3e5f9132257fec48184bb66216e5b3c8f7e60b1904f006214f35cb5a354c43f0612e13b3ff158ecc20d4d4643b67f6208e59d8eb782bd95e6f4340d8743183800435e63529dd27ad8740b8816320281d3720ef0c43376cbdadaa013ef902bd54348c50f2a62567b2944ef1e49433dca30d6c9487a1cbff75679b7cb40cf5320fe693d8f45d826c7e010862c02f893af12f0d24d285d32730dbe78f663ba034c09c41b3847ddf70421beba3c5336f8566b036b53d02c5d793b49cc6d99654b50cd55c492c522cdb9418c6eb7c5b0f9b096964206dd5cf9beb4b1721446ea03666fed00910a8c2a4c6e0231974227eb7f183aa9fd74c339a9957e20c2f7f14e0ae4b567ca2ad660d049cd288f0a77d31dc23b186d92af5a1cca538083d1e8ad74b64bb5936db851592552a81f0a258dfceb07b6074ba0152d0c90f68b32a4b1ce76786267de2edaa735b66f963bc56ee01d35ec04100b3614c05e3d59f92d510d252fb8ccb96394d356d9ebb744a93657e9ca381bb6b3d77b20c9840c70435d3a4a6a9eba28d4e5cc0fc3cc1d4492c40bfcb915a326ed2598389048c303ea214b73981364c38afa11323d0640fbcaf535c5942fa02b5c20a64b3a08138ec5a150ec8e1749dae4891cff5746899c9f1617102df734798229cd077ec8dddd4d529a0b33fca07a034105b62869c7cc5a026b727cb1fe86cd1f3f7bd5cca50d2f4f2c61c288f8653df5179353919cd27dc7bd0b99b86d9b3174697e6934862bedbb07eb049b8998876b72046fc4bc98487191d9f54980e9b7a37caf6a52d77130da0373329a193564d6673ad1061d560e297ed3f77a6e37d27fe19fcff80068f92fb42dc6545d05cd5cffba2dc0885b83ee5a8d31b599e2ba6790a9567253258f1c38eb3f4f359b3270733fd8c313afdbef35d7047abe8aa77c93f9f16efc64ff0b8b593a2202c29c464f271f41e5a33b62f8feede758076e05437eba41ad058ce5bef2e0fde27c131c93a422dfb7d0d080028b360d5c4082593d0ca63f332b08a05eff74ac109e457784a675c89236255b838a7a1d0e71c1ac61265147ac93b7623943d3f9a6247dad3c651555fb83d39e08a028640d69e71725f431885ba36c99c6bf615c47a410c5d912711b6c486db272ee3303ad847dc86e9cb3019e1db43719fe372ec869d08f3893b664cd905b0cb560d350b79a4236017d4bfd6db89e108b70e026de6cc1c185fe504c37da82e588ed3c03e48cff6c9f65ee3152bf74224ef3d2bd4ae22df0be6b7f9d8c1fa5cdd31a79ceb307a48bf75103b80288c19710be1cd86185ac84f6acf2817fe4a2d9337c47379452ffe8e1c25386a66ecb7552f5fd03b3f34ca18f2cbce205e7841ddb22424da0086055cf86e3e7e20804d2aa857310d28b4e090774a3efcbb63262657912affcbe4d91325e41e7c22a893f37bf8b0d9c526219e0290664a9352e96406ad768831f28f452ac676907a2652575971fd696d25cbdbafc04ba39cc4385edc0f1aefed167a63dea929219c056e57b68a59a09cbecd7de8333f03ee6c73051e5d7fe697af7ead2583e67bb2082aeeb9555e2a4ad37954ac40116e696e3be5f278184911cecd92531e4912b604d650a5d8809653e004959eb7c74bb03303b36a95ada6362ffa88f0a54a4778c63bbd43e60a7ff456961eab7f7239480083be97064436aea920563d841d2dcef8ba80184aa8cb4c7580c58b2fae684ea1520c5879052627f8ec22fb2fd2e1c7fa831c2d3285ded9789fb044f343e606a51f8d9056e5359e98e79b6f079d67d9dafd6ec64e90f254a6dfe30cbd54e2568a5035e28c1bd8f771997badf5645aa735737104912dfd29e51ba7577fbad0e9d38403e5913fb213657c166b4af0c2d0200b9e473e2be69c11c1134a5880144a369831cabd0073e9894ee227f88fd34082165aab06c745939a8c3313a97215fce57de805a9f585242806f4b4e3db83e1d1c9dd80dedf505028c755fb6cc99b6635695a597921abeffc883c80000030d1b94b87ad5b89c29caa6b7649d729505cd46bb978525aebe24723fdb412ff2d0cded4d5abe727a82a437c6970842d67de1c1adc1c73b4cf10970d6337db0791fee0d8513d6507b67c217f33f65a9e1c750f3d5c503e105a79668e2fc9b5a7be08aecbcb8d1e347a1e6148ecd7fe8b03d2caf06fcb2166f9b7b583ad35567a97ccc86e663ca4aa84fd4e6b57233d193678e5f26fc4e9334a4791d98c6e5ccdc0b0994ff9ae0ce33e819d2b6df2dac6dfc788271d0b3aa35db86026f5f8ef77688416098c7d799078dfbe7f3690d36a3efa72fceb2c6c58f73f3b93d00d3dc0559b60141cb36d3c1fc27480e95b489e4f0fd407efa7fd8203c33d76f5de8b5533947bca3413c5d1bb5d5aafcd7f0f499de75a95d59e410e00321b44291e99d6aae8df278b1560d44ccb63713088361c66c7d45a44da14ee1882a18990b48811c95a974d4084016d797bd6c90f1858bab6f6fa6eaff44f52e9a7f5756544b9b0d8a8659855c8e7013190fba43623787c28c4c70415c82095f798e3c009ac312d068a8d8bc59e89c1eb21c6430a39f68dea0b5458a9007d6b205165d4b121eddee561c6865f87c4194ba5cf1e552e560ae37ff3e525f4ea7d248f78976c3b9e0c5a4f19762269d349f089ef6f1980d5f10fa3d5aa7cc41df7944f180b8e4b0a0712007eda2acb42ccf4fdc87922de05326fc8f2fc5ac959dfc339a3d2bad21eb2812d85dfec6713a0f0572acbb46874f7c321ee4126d02b8d99ceb95c08b357133dbc2e5bee2bcc31c444ad658e011cdc75a68ba55b224094e83302851e6245a4f593d950b7fac824c40302b0397d31436d24c79071136212b69dfa60b7927b07d54cecf6b93451714d863ef10a469eab8d8a532dda0234b1de052ed0b8b1a83382c00b52b4fddfbce0f90d4edf9f802b76966d49a50a80115bde7b84b57cd0609db743157dc9fc44d64bbec10472835a34edea75ef1c2a9789372082da0ac2316b57a4c651114932cc098c5204cce76cee4f6ffa016936da322dafdc55a088d47ba2d7a97a44433ae8889f29d60c695f1c53af20c2d27205f9734c6488d1b1a3ddefec1db1e2adfbdc25e147805f8a2108fe75623fdfe3c1115677c0b69cc1feedbb975337e2e717222345bb361ad85332c5877a6f0d67f84354d4145d70d578e46fe7d2aa0ba4abf5574bf53111c41b0db3dc6965ce6b30b1b1932fcc12b20a845af2f7ed7217ab139d93e92089c1bbbea91a7d123b02e65c9a63d39110bb106e90a6dee6b1311a431890a360c5942d0b6df15938e49a4e56fb59e3636deff71860c357c89318adabb40f6642d66215e4bb4a00d7c6af8d2f262e03cafba1372f987fd8a27acf9119370d2e69d05581d3bb0f4c3a0d5c6371c598296cc14bcb61ad951e0ed2ab8bde01a293f75b33e547920da9a0c34238d69e14c8e9934df0819690037b84041067fcdc0a1092bc448daa4d9f000667d3ee7836d7e73bd7fcbd5af4472785ceb2bcad5e3344b1f2e9e886fa569e4ff8493e7f4f92b9e8559db05af9f009e7ecfd999f69061ba485c824c33047ddef61feb7d3d8ed00b8bc6b96d99582f6540db2ce5807b3e13d0d66d32c8c3508f3cc786ab7cba8e44e4e5ce95646aa1c341aa2f44eb81b334f1a9696a243cfed676a8891ff7bae4048662e1efb9a1e8ecd5a4cb7649777fbd82c58b9edcf8208d9fd7e8bf37d7a8bda9102b61fac76fc82617267f2f9ad4314f9a4b2ace479ff252797e8272b13588e1f28e3a91f05592088a76f154082f44eaaf0e52cf74b93dc1014451c8df9948b4da0972eec3c11ac3f65dd9a19c19fc9d0b649aa2c01ff5ae544889ddb5275d6854e5a956f37e177dae37c39ab6ab94ed931108c8918dfb651494d5c2d07c5293bfe7897ff9be9b880ca40aadf1cce4a5d2bf1e92818d5ad01d29a8a1fc198c6feae040b7da8b8cbd0efcbe67c3b83faecaacee58d867744fa5140a4223f1e154b7e9dae96fefe7a4bf41b441d26fc42c4eb916057c70225ea3449057436362b2e989ef2ebe9ea0626bd63eaa8ac6b99cb0d31c42e39cb810e7fe435474e1113b88efd8157b540ae47e7602202a68cb6a4b289880430662293d5ba709a1adac06e9231c1eba9e5eae61267fe20d6f0c7dbc720ac4d3bb9e1c74655b71360fe669419b17f77f2e0d86119bdd9ab9bd5250bdf936738ca7af16c5925dfbe8b13b992b003736c09af9d09e62838c2e6bf7aa24d3c6c21e04af861154c1df5f395c4c68b9f9fdc2f0ccad4b428bfb5854b75177e2dc11d84fdeb5e796570acf56bcc6c161dd5a48006a6a2f89216bfbed6253d03d706d83864f676d868ed53458df1b459f97f2b3161f2affae18bb05b3bb5efc72b6ebc37d6c34f871c939c75244023c719f457db435093838049190712595d2b8899122d1937f489335a6016d86295e691847ebcc35752b6a1bd22f5e74247a4fab9bf3dc65beec782cee4098e92;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h108ea73955b81cca2ac23ece252a2402f31f32b6289261fa4a532c02d8bc2c1854d2e27be7a8926ab891c42ac2d4f1f003e4b6041270f1d0f7f16cfd55f85ccb8ce2967da699c1b6062da227a8e7f468fd95e55cff66b2605a563fe10369f7aaecf35424fb882eda80b2d94ec8bc5c920f30a73175e1d4f56cc22e6099b0f0814095fd7ceaf0fea00be3f8db2170631cd5c1096d2ac47db298b8c8a4ad1cae0b175e954d4d192eb9c6a74c2394a1952384a9532558bb54febe57ed8569bc20135936e3b2b92b97e805019db19102f0669da5b6a2a5b1ae0b37440407f51cbbbc4a11df5c1118f83f4ef383d93a8e64c02bd955c0ab2b85763ca53dd14e96e8dbeb9af6f5fdb74c9c980cacf9bae9cf7813e55b5666e06d5b2cef244d3100a3a79b2572c711c6c64485c396dde32f427daf76f9fbaee2048d35662609fc5f2da36aec22d11b3bd0c8c402373988840b1e1b2d26ae83705960c67c860d82f94cf71602e44c8ff9d42a33a6c9d2c1a98a3fffce66b443ffbfff7dc0458e2eafdd599bed35cdb34f206e8017e9d00f0e93e09aeb5ac95da8c19debdcc883c537dd74bb1e6ef4ef55a254de5befc3b258db6f553415cf48e789461fc2d8b36fa52d1ad097a8a6d2820ce0744604e034a3271a37ed0e1269a5a9c9c6238afe7cd25a88296549f866e49db76015d686b08dd02dd3ccaba4a1ffb343cc4653707ff6970fc3d4b20ab57e114718c4657ad23b7f768daff32d5ca9175045627a8608001e5f41f5bb2c8f34526fa7e47d66cb36e67f9d67463b255efc876f2e3ffc2fb5afb53542b2b7a5b8e8fcecd93e378d00d33089b4ef84f18ed482edc234c3fecc11f2e1cd13f8ad0bdb2b1e989e774413142df5bb284eeb9cfcecd0b3cb6d139f28afc4660d1eb28015b6c406a84753175bf0ef8088efb69efbaed5f18dd38c823a81aca4485ab601edae620c8fd1f8e195ec17b037c47747a132b0a19c61664fd50197ffc55da0340202b8248d43cf9e9f30d5480fd82963cfc590e84ef776e0ca466eea55f62813c7e2f44df8d47d304c586cce7c64bffb98074752df37d6945fbffa3f51e8b724ed67b6e364f37c54682a67ebcadf23f68104e8903c7ad20fd6da4ca7501f7a328d5e00029776cc1045b274f8c1467eaf28a7a7c976ddbd77df82914619978f95e50f22c3d0dfb738e34acd99131fee6e683d64cfcc70d508ce4aa07a3bfe2050734fb46584afb5706107ddf31d07421e8ba8a33b3042ba6b4869ea8d67f35380b120ad7ac6c2456d265d4eabd824975454e61eb0e62edf21dbfa7a52faf99413653e2f098a736bbcbb7a0ac280dcb6d2be256cac8a5dfee868e67493710eba115f4a27c6c1eaebb25b1f9be612f902c31975d9ec2404762c7e6c1d11c462f1da3faa916a01a9cfabef7a44233f1d588f9f89a0a48a5b82c19cf00f1ff6ffc78170d2896a34f8f21664be32f11063e1c027a70355e6a2ff46dac51e812f1385212588a66646fa0c30cb457357f66284b634a6cfb0f6c913659536a21b687c888bdad25ae916921726f743fa9640eec29c5451d5b3f993ad786cded5740bf36d9bace6709de7d90f115e6bf05612ff2ab12c31046834fa34aabb35990702ab81047928c96ab28bf363fae53629859af4b3c4cd0b5fd7c042a45460fd49b62d2b7fa9ca6685586517454dd9c57749ac2237a08a7b04e8c255305cfaa1b9ed257fbf18efeb64baf4750d003efe8dd7f80316614ddeba3bd9ee77c89a32867bba552c80575e5091aa8ae0ed283c654fa184cdff5ac74570f777f33a7d5d80f491980b57d11ef7e3a72d91cf0a0ca5a7d642d7efa228147ea1272c4ef0a2ef65fd15104297a3057ade2a3095011a7574c4c251a8b24d07232352079b449cc15762b29d6b879f5c6cbf7c31e8cffee41e025b8d439ecd3cee9bd17ed01f2988c2caf6da3a2e74e7f7cf41fc6f219cac7ef3e9f105b2f3c7fe774f7fe34e1cb28e2bb00abda0dc92ed92eccfcf5f8c354ad72ce2c6cb061a71c898a96ac1c46739fbd61043d1f42a47b86478327b68dcc7192428322e455ad04aaded046d0a74fa0088abb8c330fd86ab5139b106299effcbf81abe14071a8ad1c74443d44c6a332cdbef88e912b2217e7c1e9cf00c13109a972946fd0f990cdb2911ee320fba00f8a50c6a16e64f29a681fcc771d928218a1058069e1cfffbc1968451aa99fafc51cb61fcb24b05cf245a7d67ea665865b22c6d0bf092153f067f0aa347502e94acb0281c2d96b9caabcf0bf28bcf17528b6cadf47dff1e5ee9533d723ba69c92decf48b8b40e1cfee57e53835d6e11c578ec674087936b9a1804fc36eba9b063f137e1cbe6765660ad9d22181501906c8d63e2fd18c7bb0db74fb34d1c72f1e7514e1f4067cf8f5093c8ae31a5112aec761aedbe5f02ac072c3d145e095d9a707f43a8c8f14b96cc228a56a0a2bb67d758329316f5024b9749ab6f8474b8af580a67346e3f1a668ddc294d6624dd262f2efaaaf61499ad559677e1b8215da688a577f517ba060aff1ec410ac71e2d2ae88ce21b0244904792ce0a6726b8c056ec7e2c893bb758242fa63c6f43e1794a1b62ca294ff3b399c4e41e4fce1ee6e941e80914ac69516276de38b72deab73d990f203b10abe64a902d6fd5f33abeb1c458353d17af4bd97fecc15cec4f09f15453ab4e8a60fb54b20aeda8ab5bc7682200d65d0432335e52f4b76a2574590a35ce7498cabfcbe7f70c32026891908298f51025cd0cb21c8d1d8b549d1c9ab99090bca2a6b8cb75f59cdd86037b7c80ec914716be1212ddebc0049ff09e43a9b6df5d2f933459c2ae11a25a30dccb998dcf3488ed54bd0a439ee0e74eceed4db14baeb5c7eddedb53aad0bacc024a847c3b22245002df1b001912b838abd2922220fbc3e5023cfd8aa725d496f3d9db720cf5c95e6f240c4317935401bf5f91ad3f84801c64a843d2193ff5d5cac344b5dc30713ce14d8da66fda3b0ebd19f03b05d7a64e3ac00ada0ee1793dbd099a7e1b265b93fb8f8b94154c20f48eb25710104ae2729acef96b7bfed4a9e65a0fe3cc43071833b26e457638bddf2c8701d9b1c82200b52f92ad89c76b5b9246353b34ae9c586262a2aedba4b120089f01db019827624a6289096a5e2e80aa263770e0d75bf46bb15fa8edc23aa5c303acb97fbb33b6ffc14686b9c28ca21ea581c6dab8ab3a01caf3cb59c0e1adef9ebb2e087bd752c875fe333e6828f3661f19abafd0292e0b82264cf83361d1cf915a8da965c7e7ecb6dcce6e5089485af45d1c6bc557b6c9324659ff2246c2a2d8107a0ba65ade40e51f5ffa0c523ac5c50da0496474557b0364f85b52a0e298de2ec7f062dabc2f300bfe1b3d49d8e2ae1fee1ffb3a9bf5093f45038e148db7fb81c376729d8a5887429d171ccac40525fd1b4821bc5bf2b2b1a7ef9cdb961f2ece594d9769cb2c42a1509b1ee3460ea75d991b40ec139eba307eb1ee4bf437cc7935b8cd4a79457259fd29a8f161a9c69894e97f46667186f558f3fdf08f0aaf06548c80f0448bf9ef9f8ab713efa96b89ef782dfab9aaf855b157ea9fd6953722782b03e2691a973838195e73e94634cd361db31ab9f4e1da15ac11d997a4693f48995c3bb339e85812696cdcaa302aed5f14d163ad5d55c845ba46e2161e5487138ecb0b1e8482b5915fd9654332cc1f9373d3334a406cda85c06d33a2739de01969dbadae9534b6b8c855ec3f162d5fea46b3528dcaebf8861e15e7c84545e3b439f7fd18d7dda3bdedea4c843a044add07d896c6c16190e27956142cef29065a42d89254f7cf664b6d1c3e71ffd0f89e4b2edb9ca6e5aa711fbfc26beef5b7ffbdeb2f18e3c56d3ca1d5b5a19a5ddbf3485673f7c57882d489cd073f8682b79b3400088d54d5a0f822fd631f97e53aa1c9415d34295d30d1e0c3ac7bc302ec1e492214fba15eb394857c3af4c1173c2f5886bbf6b80e3413af1e7f83c48cd4f6e65ced66f57e1329795ec2142f9413888f2633bae76dc7bc3ea1c050b172aeda9067afec4123bea4d58f1e08c5240658674b6b2a9c56498446a154787efb85e9fca7f7a5053f429a2d9b05082048a6d81d97126a9da82c104e806841de0e14762806df35cdd08d77459cbe3e149b539889a9e37bfa719248bce9fd574b976d0ccb7d9be2ab04138054fd81108839749c86792516d5a1b80045fa7697606549ee34d6bb35d70d8f8be44c0ef160a37089b8a25c7f95620d0e4b0325f4553c09dc01b89556670fcb8e54ebc40d42b1eb8cc8495a6c1cb92b3b867b79616306bbc93bfc6ebdfd24fc299746803440781300ecb51abf249c607bfcbc9a52ad2ec9506730c3d13f98959d63c2c4461e9c38e1f6ff66fa31b1402eda2c0fb0fae325b24724b74ba17efe793df4e6b531a91ea9af1b3c1f0ae2f071ddefadaa57dde253b8f948f6f80bc8bb4f7b01be01c997532250b1fb180ecf086ff1a680ef311675f2b1d609aec0e6fac94160dd319c651728cadc0816dd9f9053447acfeee9a266e14488ed693c4e9483814c91c175a39636eedbe0998812f0dc111f15119b39aa4e60d326a50657bcf7a6484edae8fb0ac8c1e324257cce13ffc92161c35899ad89904373d597ade1fc95e0ba603b97ea05d5fb9e1c33f003f31dd261fb30d7e7b63d7269d620d3f21aa8524c2b65eb84183ef9e87b49f278aae1c87b9077449528c0757e2ea20131222c8e41d547788f79af2ecac097bbc01b1d4f222bc0126d51ca50a2d84ba99629aab07e0982fdae041d2fc144eff23fb99b08ee72ba16190756e83cc266bc64bd09de4f148e733eb91b719b2fc1dabbffe381266a1fb23458b1b456fe91f833d8d467dfc6320fcdf0cf9fa0f8f72e69ecd896569fdcd78153068f9ab2996c99bb1ae3224c0e4df45b1b1531dde42a5b8fbf532d141f329416809f3c136aa0c6f626342ef1eea88bd740e62a601e733230f4beffdc25929302c09354db916995f5955105936f3717b9cf5315b54b7c4d6057d80321a7fb86ddaafb91b462fe429d0a6497945b0b74a945a255a296990c37f0e80cf9de8dae0b0794a7cbfad0471e4449b935bed7a2b3ff327887c44295f3b8734b03342acb97adccee61e171cd3b7e062bf0f6949cb1670765335bb22b5d0f1676dff1e1e0a9293837a5b566597fc3138dfdb0587302e5984a5d80d1200845271b070c55f9fc11f92de7230b0d25628489befe209d790aa30190b200fe0e1b4396773a133f7e26f5a398a7692ec0d3e3a0803076de8b1d1540c5162e860874f507ab166e7a22b66208bd32135f6f515721515b2e945e93b0dad42fdec2edb5c81e029a69a02a8d7f584a4d3da1ec5cf6149e67e52a19ba0b95e30d450962b66a49ca26117f864ca9bd305dd5ff92cf3d3b1a874717ce1f3adb98d40281985cd28d29f2f21d4a87a3132e75e3f78bfb9348530967bb3b8f68044799abc01ffc0c87fa69e38a41d5b98097e7e5a20c298e819f511e9ac5003cdbe2b73ac6d37047f69522a9bc33868f574963564e41b5677576a359d352e86d02c4209a09e2242f5e5cad5ee5cc0a2ca8ff7bc3ed385140f2bfa7f1c506dbb60468f7de51eb7a5945455eb557e6cb102b77ad8a8c640b28c8650e247bdea9fca5ca74b822554f418f50c7e3c249d8290fafdb477fa41fb1876328f425720aac40c47711e4772565823319c2cfd2845888a7be5e77b207bff26e90cbe4310e2f6312728f605502694b2c104352c7e4e36a18dd80f471440c9c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha48c8e795f228cd9b9d28f943189f55af20f1af25cdec5a178ca37a5e39c573d075b17cae10b6e03197394ee7e5b529416e7631e265cf05aa767490db813a269175f9934e0dee2c89824fae54ae3c6e1e62e47ac03d6f7eef041eb9c01e13430882d087411b23db7419d05b9576c8bd0f3d8cf9c60d65e5e3bacc657af6599a384218112edeafac4989a9050e9b8833f0f318f1f00c8f13ccef32163debd93e09f2960399328fff19b82a5c1204903cf7cc92c9da2e7a96860bb20c70fa8f132acef866256bb8ae4e343302aca3effe7bc74cb0fdd06eb7f0befa81c6325ed70fe6f4cffbade79b604952875acffe9792f6c394443759618b4cadc1d6079857480bda15cc1b9fbf02805c9e67f2c3981afa4db0d4b32b09e7e44f5479e91f88645ee89f38bc08125bc9f167ddcd83a8b8b6ce0d2e943a1419171ff7610a535096a1c041c2f5ceadbb65cc2380c640787f7e9f04b76eebd3f5554f37eabc27547c33a393b4934bd10829a4284b0201bb6b3f5d19857402d02aa5fdb2fd733bfccc3287c25d8850425d35c06f4e0a7c5ff0d6fc4b384c8bc26f6db105cf70bd9254a0e32e669295e83e91d92669909fb98c5a50ae2bc3dab9a9dc073dca94e377bd927d75ed37a88a2fc9ea04ded96ca4fe8ce21a7d8e9620dc0716f52068ef268574822a1cc429eb4d31575d225d08e7f9f34b5f04f90e475f7957f33c3bb06c4e608be4b3022c2805e86106d1270375fc47b1f1adda3667ac3a890650de918ef53fb27eacfad134774020981b55693ff6b5e5579fd96bffc9c53f12583719c912a110b65ac031faee2e1f0cdc68663671e6cade8a59f96888b7a443b1febcddd8442403e505833d0f40b7eb6137c2b774c7354e5a788cea8a3cca6d6f97146be1cfaf2398d9eeceb50fda60c41f86496a40b06fc6f7f0f80ad50dee8da34a59086af3cb6728783efd003dda9d38cbfde8140fe77ef33a6617a3ee8a4dd34be22145dc046351c6faf72c04b071debea8fdacf22a3aeac1ba24200df05c99419d1ad403b9ced8bf0b5a26118f9a1b76507fa6a6b43a07b473dfa5ed3db8f4eabedb2790f872ac04461a88f93682c55a7416baeab2ee83864c3d1d7cdd92f61f6d16224f32a4083fd3f47f2d60e70bcdfb50297689efeeb4aa447c0cc3b49d95766305e6437eb068a5d24d0a9295ac6425bf2eae212ae85ab540e313733d42e05f4b64e2f8096f0a78a3987aa2829d2c36b8d0faae63674f8a49d6eee6f1747703fdc1dce21e40533b773274d56b28c4930c5d8eaf06a840acf7ca5b9ec53867cee846425cf48cd2b14bfd9787e160f5f055ee0f29356f3d055858034dba4e1627affcda8ed221dd3c097c51bf2c76d7676ecf0fb39e0ba706bdea88737e10e1c56f19128c9daa98bf41706e17a97d5470e027543559742e19c453f8b4fc44b82ecd31003c942e863e28ad45aa44ce6b6e7aff9250aeb8b2087f123468746b1df149256db1234374a3815a50d664a175b777e4ee95418218af07874cd02b2792428d4306f6fef2e33239d74a301720e3330829f46553519efd2d56a50f868f6eed406b2db7296f4c456ba0d8d04bc11e3daf301aa80db5edafc0c9720529ef01530c35fb2857ad18e3f4ad286538abd70dda452cf2ef668df56d42837444fd76cc3b69ed84cbc01d863833499f59351bf4bd9334319b3d97c6f4373abf34074f0b98ba2ac796aa0bf0853ed743b4588ad97d241664c0aa71f98b7acf8b15b3581dfbc9019fa1e6f86ac20bf69b55835cd0cbeeac47a98a3c4229829f471abc86ee8e9d36899b826211d38474b1977eb957b931a302bd2d3e312efcdb692ecd63d830e64b1d67ef18324e4cfc52b7b47863545c355901ffb161468b1bfff7629f3068f6a11573b97ff575f0c67a4f25ab124f5b4ec63fa859dc5397efe1aebf73c4e32b8854e63bdd9e42dc5694196de2f5660b2cdedc490af96e9533cfd2c904518282cbc83cc7f24ea34e229132d670993c59de91f2fd8b5cfd007e69469cd9b664853e65dd3d6d040b2274307365d5880b36f020274cc4fc959a5326893760f591b2a91a988f88927ea8900eda7c17ebe7537b21f23bbcfbb93679d73075e4a95cbe37754b39674e06dfb316d7cd83d54b8701193f552f0911e143415e929d9a2db5852bd1bb9a8b911176b2b9dc51d46e3b51cae1e27c69e524cc3523684dc07533cd10e677d93ee6ec209776b24efa9141df4e18caf27aa3a0cdb4d97723dd28574e3c6c915761f1c3f9536ab7fb584d9b511ead9c5c8d7ef91b1e433326e8b38a7ead78dfd7e37663aa8f84d8c7ece29650313cf4ba9300f00cef3fb0cda299ee021afc519ecccdae0c1760f65065ae82e2cf333ad11c6db40ef68178645bff4d39ec27ff183f4eea77c8d0e766a13c12ecb6b0a62e0eb9915bbb7a6d2fc01e61367245537ac0de82546e3dca4f0f0d892110493da46395d8c54b50d2607bc253efeba8a5a37ac241b647a13136ab1ff4004cd0365a60ec07962867a83b28d97113200d235047fdc6c698d3f59cd4dfad1ef42bc0e756c4b3e81e54f501623eb1c2e3975f67d90fb4aa4cf901b81314b698af5e6f8584888abdab9f93ee699954db4acf4887210905dfb88e23909e470be163f44175db57419a7bfc128da522aae6c045dc28d9ff288ece74af399514d106b3baf8f565a91d09128356e5f617a757c96ce6a50dd4ef8502acee1d6b9b73838b5feed4d78a7834dd84afafddad6f8e5cbda980fb7056fdc4b123b73b47fe5bd905836d97f3c97f939bbcc5635e6f7a18a0c935007f330a753563d10695aee7c32cf9e8e4aaf9616422fc6670c04b88e36bd84de8b547734f81437f3e518c5d2f24e50de0b206b1882e2d4ccbc40f7b01b82617758551252898472b9fabc1d6480446fa37c9532b50b957741e90283cd1f3b4370836eff2112982cb01b9c08b9ef8d91e6e97e6cc0bd7c04071faaa5d4cb8c6ca14f73355d78ea1919d0160ae442a0386ee0b74836d432ebb897fad3b8bbba1cc44644a801bc406e6a930112ce03e82b35269e8aca74bd6ed40d4bf4f70f4bdb610b0bc3d1f6800b9e52daf67e6e734ba31a66413aebd1bac7fbbeeadbc88e5a0b356297b1827662843d8974447adc374bc803ac39c0b526c3c8317c89b90420d178e7750c172298b9a2b037fbab2a7f4d32e7202ccf2933abfbaf17947bd6c5dbcfaf649502dc2dc29a324870a8bab75dd699a21b2c236425761f0d3d5d97d6983a98bb155a5eda482662107f73242c42cf822f8d2e853ecb810679b87624160823b355cbdc2f13c5094956f902eb3c3a29fada1b4d3d556290460854eb15d0c3b4609f000cd0c938d589962c7c29b5e2f4185508b70f17c5a81dee427a1e838b80567f000267d796c1a14ac66871523dfb6aaf4f403bbb937155f524701313a78a4c9eb8e2dc01980b95c1a8855101d819c2610966dd3d1d0d736fd111dd828249eeeda9c112ab168567b9f2707f01a12591c94a7ea63a860fbe91de9973d3f5e82277ad74cfefb6958996ad771f0e9622a25f692069057a664f1e7c00e6da4c00487a9a6ce61f60df9794ab43950741e6ca833cfd9d2bdb576312d7b1ed02580169b21365130282a4820a36fd324568a71b5dd43151a005e1dd3c5069791a4c71462c921ca62638a152ee94f68a5ed6cd8d1a3f83d48afeaa00cab734aac5e197f16921e7729e73f0a5135e458265025e1a051e8060e885b912f4a7450a6927ba6ade0aa169ccf5c0b50a4b35402d929b597b18c4d72ab98cfad216d7898b9cbe5d20efcf128a5ed5d98bb830176a9bc2210a9e3ef787f8957ec83f23d54d44a58a86325106aa920da36551e4f5165e0d727d6596c636759caee2d0715864ffce72cb37282ea1c68de537cc2c95f94c8695879046e31bcefb54545b06bd6ebf5cc7c6ad47b4cc41e81e61cf0a039877f2fc671fca52a059e68f5b94f7a36e34f48f762346602a8ecd015015723db9ba4567b5afa4c34f653b433480769fd86cb5f3b7b667ea95b3da937f2833713c2a855c06e20261cdfa2e10c620e306fbcbb42591b819e93de2725cf2928a236718bc14164f7adf3347ce99efecbbde330f1abfdc56e5ba78640259976255e085681da3d95a7b77e98622ec1df0f0b2bb3da1421ef9d8d253ce48c082bb9d1d1dfacd66ae22cf52ed9e8c2750189f94dfbb7df9b2fcba1fcd3ef1294372718c422a561732a04fd849bf95169dbbd578fa7fc708cd929fb9d9e1d5624b89242d01da270a9112810e4d2f86bfa7a11066566e636f69058cd38db5a4b072f9e8962ef7db72f712b9a82aacd54825dd708cf01dfd24afb77270856fc2afec7fef2b0bf49064a68ad37928d0d22e3b918ec590bf95243f6aed02f6ba8c9b96e2355cd825538c84843903dccd05d0a9a8358f33861643d5ff269e6783a82a6e503527a2fff206a3d89d140c4f6ba31c5d971131f61c4c21befd4ebd367c6cc8975eb740db213e446b3de14a86c7996f2417151ca5f76c00a56ba7bb75533491d7ca0a800d29245ffe931b8b7eb28d41bfeb57002054b0049621fd2fee2d72a19d520afca1b2d39f581435b5b9cbff40268217332f0039420d88c9ffcac8ef2d7a3c9adf2eecd9d6883c32cec2fa5727e1a4b96307c8665acd461006968fd6ded84a8304e2d71a968fd07dfa5a1e1b86f20b055756f11e8c11db05056c7aaef5a62f893660c6f8ec86bce09c82eb2c78b1da367df131e7850d6e2320cb59c780ee88c2d501393b8d43007c6451e2a74ebcc17342fb30c19de41561855502636481f9b9af8abaccabc58f8f4f019089d20b7788683467591ea07edf44352b927a9e33d6cc89a17d560c7d1f2a5831ff722de0b416fbe2566a9c2097fb8bd77d42a805a1f60e181129bceae09146a4c450794565012944307ae343b6d39fc29e89a8ad4c49229c0dbeea29a8ff86a680e12cec8470e6b898c9477f21275b69fdb7bb4d1d9f39c8f357d096a1f06315bd6ade7078480afb9a6bb3c76dc186724ad1133946744af6f9e8d23bb7ce93f921c74ea099d3470421203c603edbf3bbae9d1b2dcd72305ec20b921b076c6b368d0a6193e3359f6f8714b8dbe4a15728d09a25bd2afdb343e7977174d51ab02ebd62f253f85ef396f0286a732445868ca72084af099900cec93dc16a569aa9d1a67c7002a6eee150d505e62020d41922935302a3649090d2af23f86b6f81036e59a79d3bcb2737866427256ec116ef35d1505b3b069a6511d06fbb13da0d9fbd9509a83078f912c0bb3f7372700aafaf6b518eb64e97d2a9dba863c1d519d5bd4e36df034e79261e6e8cd5c58fdef61411f5f0c6a7aec37cb3c001401332b9187742b0bdf99a05cfd39e5f6aaaccfc62cab071a74373bb89b1ebd8777969104815745975b0cc89a79c8244d8ac559074747efe2a8b0bc6a7961b3dd78c9e2a44525fdf74578d9fe702eb2de3bc34d6c21003645865de6ea875d9ccf54d76baffe01bb9118ad1f5f8317bb9017924c92558212bb9da16c1713dbfb8c51207921bf806c3c59d5e91064c221a511c6899a3f2e9630e9d4ba3d0f7db12bb4a87a5a90ce9493a517b6373879319ae3959043bd95c01ece6a2d8bc14c8e38c30650129fa13e97b74e9d1d011a18169ae101cb738c05c324611ea38a855705c8944b7037592f820c728a736339442779b73d8cd7c485fa851b0393df38e635bf5c21bbf8cc1a87d875638036e874579be3f135230055ff8e33ff078f8ad26649ca2d9c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he3c18f3dbf41bab1c747d29a95fa6d76ad1d3ed80658f81616cc428d41947a26ee2022fbcac95a9004f850bf3a39456abbcc0b4a60edeb5abaeb6c253af88ce7c8b9e8700427ccb0903324b93a337d65a7891a87d06a851b96e9c201fc5ee08eb31efebc759fc71e1bcdae4aabc1c450f358cf19588f9970d5d9c5aa5163f9f1d4d401a967fcdb3f1bfec88cfb63b1f8aa0a259d09cbd951befbfc9e7abebd052bc423d12edb57114077722bdd4da734fc01a37731de174275705fe29c614e2d70f22f120cac7f98c76b15b7b4be0a86a65d6582ad6d7814ed4470d109b17f1783ea5421c776fd26efbc15501c48d5531ea699ef0cb297f2f2287f428072dea0fd6890086b1c935b870ef08788b429f586d86945e106702caef9e226012bf75f886fded7d9d1461e4165a47b77cf42950755ab7bdf97ebf30060154873d41a7f178a5009766fb0e1620a380dc3cbf7345a6441a285f508c1384c586f4795db2324e8abba039df63f607301a388c968f36e3fa61f669fa47e4acd413804e376941ca6b036911cde3f26dbb5990ace8c14a662903764726572801c1e11da007055524c272ff81f69f110fe1282c986a54eab99efc320131c9b1312020293e90bfbd739d258b7151ee73042b415e210824361e252176d03e593c8d579719771978fe7d76340cf355edf7306e70e6119cb825bc16a607bfc53fc4d5f374690a16d70d3df92b2c873b96e30a427a97f1df4b4950ae7afb04a5cd5a2252645887a302df4372b470fc5f2c9d8b1cab16854a71a5119f62a6056b994928e14e78984a9962a8cff1b2c7e6ca5d1f86c8b25b5ca9bcc11cf630aeacbcced493312c9b1001eaacac5b52cdc8a35f46a7908ad10498df4a0c4fad508462f3e29866df54c762f8be90218464dd8f59d41d41ddc112c9f98d092eae36161ebed5903d3ad777c702ca81c076d99fc7e25c9e3eb360b5f899eb138c3b57efdee460e576be3f79565d559b021e69496ac35a9f2f1066ab1179e28604622db71424e906097b4535378c014e5f58180476b663cc1c55c64023a6cbfdc651461bbef38380da41bcf47710af0d65a01620981e218ddb9f7f40b5a17fd8854e93cc7be805496bcfca7fb8619a1a5ad889d77b63fd2a44d2bdd669449ce168972a68a0de40b33787da0801549669edae3a841fb901d25135afd117b9c78c5fdb3c5198a77e8169f369e0572cec3ff18b9802f770047130699a540c3aea83d6517147b22788496a4b8944844f729e0efb86600bb147f24ccf45f48618c84a403fa09d7091dcca1618821a1f57068aea6c73748d5bbb7c1b117fb4c8b45b5544a53a8b05c8c5259307a317b4789464aa9c6b8fb436d6bd6f97d85d348726d59ed8537524d29d7eff404abf29a31cefdb09647220ba54aae16c89feba2278c678772aaae120c2cdaeb1da8c1edfed67dc43e71349e18cc458434bc607e7a67898e5b757e612f925cf1534a1bdfa6c40581037e8f5e92b94492dcb9fc31fa0c5697bbd61df5c291c4cc5d565426f39b57ca784916cf2747dd66820856af720f07180427eefb284a5e64e926d2dfc70c5cf475da2c23eb2e849ac479d7eaa5e5c937d10178a3ef4ebcef58d951714719dea0c00fc6a6ea0a38d09db672d62cfe15d8ed685c007393fab4aee266b8aa571b27571ef15d53e0bbeff454b69f6590d0459ea0c06e798f094e1f8f258a3c3193b7e76c0c63999a66f6dbfb9d898867ae14c7d6ffd0058cbf9ad8eff9db237c1f13a2155088fb09ad048dccbf227c7eaea0ca39422565e93881bdc55b8d841bb6a55805d3658e88c565b875a74c32dc189920cf2da0c7e15ecaea22244c5a68a36effb9f195fb8d7d3c76e554e1db79319957a044c322a3d08ce26a54de495179fe8d5c63ff6b5352b41cc92ed8d5d031b82d4cc7105359f9f9a81bd56b9024c80fe2987e328dc1b3ba48ac8a7bfab485cedc493fbf36e96b7c08cdca8ade6df69e0891824a13b29915a7a37ce763a90aa82898439205b32b83741a752055421a2ea5d6b7d62b8e32acaf5b95ad7ebfd24319d39281207ce8ca1ba652b195f862a02d4810ac833fae9cb82bda79f097c7cd83c36fb5c5b04512241a2e9d44abb20bf765fd9bdac3d8e0bdc8f590812d876dab1ccbca63e838548f6d48b636e8c276ff4a101428b863c73a5a425b0d827fa63af77944293e26b3fd1433f3942955e290e96a40e4de2cf55eb3984dafaf0395f09bf99b82525ff74fedfa28458b57491d1b4b7ac1f2691dfaba8658ff7ad6b06496c4681143278e0cf38f647ccddfcfbecc21ff384a37b1dbf61d2057c32f4615e4b967d00aee2059e47f8eaad37f7490f8984d8c7ff77e850cb946b80d948913ed483f60dabbe75fb12621a45ee2d3c58ad64bd346d192932a9c005e38c7b32beb48d865f6eb9fe23f41826943412a15170b0581150f99978a5e82a2527242020d119f0b41955c4788beb22be0fd16eece74ae79aff5063e269442179cf078ec8a6ecfcaddbbd72cc995ff0e867bc95fbd8bbbd882e5aeda41d0a8769e9c5e4847f2149f687b30913fc163320bf3b27bcca71f5d69c2685d932ceaadc2a2439de1b477a444f57967034d3a24990384e0ed65a3245d3823931f160d975b31e8f5eb8749ee318b6cd2632a268b95e5c9c375ea5ef7d62d28ec531f5148956af8d3b1ce1de7a26ceb4be8278419fcaa4ef7cb82100f4613e444972478067e7039f9f0176e92f92f9cc537cfe9eb739b50e23874e0b2fee6922b0b826882ee4ca5bd4502eb3b9cb437215144cdda6f6403657063b35d789769e453a102863b66058890392db1ddaa2e43cb0eefb7f0c611dd249311efdf21912a8bf457895d3aff538d68c0eeaafa799cc1a7ea52b31ced0ceb318532d8e4074e616f87584d30a5960b2be7ce056954d049b8de326d507c66ea2a123f30b8d9ced6516cdb78e9dae88a781461205d37d28d101383001c66be0219f5f72de530391f65fbfdfb1aa0a9e07c2af3b171acd747b8edbede22582d9bb7c01d1de3f01fa5a32c859e00e2cc63fb20c706562dbfd3ef7aef21d0fab9db70e4da3b7c3a4084ec7a3acf6bd8405cd2e6ba672004035e57f54ed6f23127e44821bca30da6f3450a190304099ed45737dbee73a8801a0ca8e96648d9cbf2d4062908e1ec9690c8ccab82864ff3d2efca82ec85cc844cb89e11b5346feb40b63d8d15ba2b891b6bbed476d16d78f8fb792e53a773cce5f3fd16fb68dc7dcd1f17b254408206f2d924941abfe026ac6c025a0de0c091153f9453b33cd86dec6a262fd4e02aec9f220a6cf31666f23f54f21cb1a4cc69fc636dec9b847819be38bbfa7d8cc9af504fef711aca74da60a91b4b4224b28f2bdcbe89e6fbf14eb86347bbcefde9937e35cc0177028efec8c3e63b6a5ec9c853a5352c2fdc9d3541ecb7908e4e8c60ca6986fe7efe44245335043bae17ad7f8584e94e34ec8821444412b01d555a3ef44da41fcc37888858c24780715f76b28244fdf4b1ffa86bb26b9a8839a0ab4f5f3f590b627cb66637d053b8b49dbc194103d1defefb872655474cbe3551cdc72d4f9aa4ee6c76bad6f55759496c77af9daef804c91b68593e1fba7f3bd14aa56ec5cb1b064a42974d1a1196a8b4c297b91cc3bbff38ad66090eb741f2be122fef7f7adde8e5827d100f49bf918201cefe1cc59cabb0d24201fd06e1dc9455dd73920ec02a5e1423c869c94b96ba53912af216d115ef3c8fed00ab2c5002571e7beba0f2f97647ee5c47034587dcbb618672289a54899061a547a56faca1f40416e62cac61fa1c0f01dca45ce361948cf55ed11a6a751165f0b1c30692d4774ff73f0e4c604a17623b50ee1da17c5811731180167ef8a95b4300056e35275ed851150fb02abbc103f1e8647e1384b6646800b60d8c3d9a99427d3444f11e67501c67559743d0b82faa2483597121e9ee4f8b765b9ff2969320341c4a746054e7313e056bd2915bd6d3b1fa1dc39fe175e00b77b3bdb721b0da13973e75d992900bb9f8b7c4261f7c965b63486caeb16fdf7b625160b796817cd2f75f3518bc7ff3ccfab7b1dc46d10a006849471011d034c57b6b580c8661cbea2f5736801837d6f0e56da6706677b1d6ca2891276898b1e9c882b147ca1f0d8dcafc93da63260972094b6fce6fd89f398f7d377b32fff777d9171830387c624affc4bc70240b7806bcc145750bd064c0c95cbdf3a73e7f20d0ce4b1273b79618d1ee99513d6c4d386e4a541fb0e7ff29f49565843599549e9756bc27e5330e0fd8c14d4a7267804b7c7a8c40573c34f2e048ded5ff6fa93701c8258563c57dd5e38717948167a7ac0581d0c7508c351b9f4231e396bdbc07465952611bc3d9b084415cc5136de14526ae53654c9b6bc49421bd187beda53b39824a4cbac00b69bb333eb882e159026d0261997342ea7dcf72318ce23cb38cb668253bf5030c771ec765da2ba6dc91625cb706f9e6757ad877f354cfb54ad50ba4f60a524cecfbcf815c7681a8e2005cbb0cf61abfb3422d2e12e8c0a56b3d4f14110e86b84d948bcd70ee602acdb83407309769ca4d7935ec3ea7476f363ef7c8aecafd07c9b279893b0b562e811859186a70c777ddac146b1e19cfcceb7fe4d260a4d862867a8a3aa964754849049a2e7f663df7ef2209bce49b79e5a83fa6482a460e9e36db4634bd9224e73266a47e3f8b9bc81ef3945fdde82b19b7ab033fa2b62aaebf773b3acbcb27e7a89138a13abe08b157a66d4b55c715af2edb871ed05bb1a0f9c40c4fb752e66d99ff8bf18929572f134ac1afb94ac84dff127c3203e228bd9dad6f5f3800de29d1a04ed2e14774793c16f87d09e5b39480a0a6cd1d11e96349746dfcb7d09d6638b7122f053d419648c50d2603a04c21ed6d12d66002250f5ae5bf4196cadd2ccb61fd7e4e8344a1db5f9b41dadb29d26fbadd37310e390b6898ee6c029b5cd2f312dc23420db262e49af4514f6db91a5da5c4dc08cfde0db4ee3437d0a49c369112645e8a5e79a763f265e12eeaae2136ffd1cb51a2d84517b52091527ce7e58cdeaa3b0193f0c8dff3fd217cc30a518ffaa5e878a23453db55c0319d40ca1e3c285ea36ec553e6594a1d47b082e2df420d8ff06b1729e396d48edb29cb1d3ca7f1a62b07412c38f3fb6f8f55a21351b98c633469e2f7c5b2c634e0003dec646d68b26b0f41d51008817b020c90079257fb78f083cb012d13a2ebed3bc4120dfc27ef789b0f6bd61ca0d896c4e1d785284fe5011aed5e39b39a611a03cead9ad81d06f7d6ed1b08c47b455ef7736adec2021ff18c6be804bace545e4edab7bccb58bcce96f53e12a2d7fcf3b3cf7d7477f04097767fb3561534166f296dfe52e947c18a78742d6b67c364801709ea16dba1830ffa79f8f8ad66fdf891e430f437536db3bc9230fda351a24b81ea6a7da9968af4bb5d7974bbd838d0e914563d4526665b68caa7b4183e31e80127f785a01c5adb230dc59fa3329a2e8e368f52c2840f8f2ed80089abc89fc7383570fa55be8a5a656263e2e0e331b5e5d31d1095b1035ccfd44d7d2acba1e30ea2f593f8b09c478891001b46cc5a458b3d1cb77ad01319624245e94e6e71216579d1b1e1d0f02e3735b0a7d309f8672fe021038c974d62b0cdeb3f0a9dcd2d6a0d093e06d93d74ff776df58f43297c62093fec06e5016ba462cc4c165c822dd1a9adc3205e584d8457b16aff99a611f1edf6f28b9a30428ce3eaf8275409a5878e488ab41134c9;
        #1
        $finish();
    end
endmodule
