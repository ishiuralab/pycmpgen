module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [26:0] src28;
    reg [25:0] src29;
    reg [24:0] src30;
    reg [23:0] src31;
    reg [22:0] src32;
    reg [21:0] src33;
    reg [20:0] src34;
    reg [19:0] src35;
    reg [18:0] src36;
    reg [17:0] src37;
    reg [16:0] src38;
    reg [15:0] src39;
    reg [14:0] src40;
    reg [13:0] src41;
    reg [12:0] src42;
    reg [11:0] src43;
    reg [10:0] src44;
    reg [9:0] src45;
    reg [8:0] src46;
    reg [7:0] src47;
    reg [6:0] src48;
    reg [5:0] src49;
    reg [4:0] src50;
    reg [3:0] src51;
    reg [2:0] src52;
    reg [1:0] src53;
    reg [0:0] src54;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [55:0] srcsum;
    wire [55:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3])<<51) + ((src52[0] + src52[1] + src52[2])<<52) + ((src53[0] + src53[1])<<53) + ((src54[0])<<54);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a2a9a8d91530c08514360ed93f23453c140826c17bcc1f8f9535978253b542888c8c005eecb0a0844828b972dd5f47b97a0888a2dbb8d0d88e07e16a3d0fb3d4c5226ca9118decc09c80cf74f8993602459e6d412394ffe041d7407de5b5ac2caa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57ae6b25f1fe56761e82c73eb2ea010b794910281d3ebe0e67f73e75f2103efe4d0d2ad65e03b48dd72e63be8e9187d2d55bfcf07a6eda39400c639de958f11aae26308184fa789fe6b032acf994e0179c8d46e58ca29cb79743f20c3e255964c9ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23b11052a110dbcc2a32f4b5c07f6a41e4fe964478315ee07e4d0c50aa921e013c6e099a249dc1884d6ba618c14579b7e7bd58d90fedce8d534ccf83f7be99655b448cff6a63954de20683042fcd0db23df0ce7f711976e2b3d797ddd62931c01782;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7b1eccff2cd59ffa4a74352fd752527313ce9416691874ced546218647873dc4c329ef52f06bb43e24d2433153e651568578fefa3dcd9ba314e1d4f011cd022f0b8812e307a7abe92ede3b0f54ce2de6509e4a081730f80e3120914e8cd3263ff56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a2931a9541213ed8fcef63b3be80cb572dc4d8118713a49777e722d99eb98f062da0430f02a9073a87c2e4a61604d9a749ebdcf98f25ef07f614ff92b03892e9ee601a6a7ff50954785ec1f6a965132c3431caa4fa7254842d6629aa1209d4a817e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cfaf73bf11fe24f9052141b9f08ff46c74eaff8f8413c439d77670c274aca6c61cc0e107f0fc14af49f791268540240836393e6834148961620c0c2fcdb4975216aa6a8b069d1f3d73ee48ae821bc52fbc4bd896e6af6dcf93c6c0756111ef67000;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdd8e66914f0ed31f29832149bcfe0cf0123213bf420989dc27aea79ec8106e27a2209fa4ddce6eac9e661ace8f514cec70b1105c0039c479d368c71a7e80aa866682134a8655b9fb8209dd29db676759ba22775094c8765a387f4c73d6f308fb952;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1839e1445785c1d4ca6c2a27aa203a47276c5d1c6a9e0338021aedeb53765b2fc2543460042c784619f70c82c4dd5779ea09681bb90a828afdb4a3820cf6aee07ec933b7c70f403e84344535742864f4810be925fe6f3aa23b79647fc2a86429c441;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35ec718d2203fc06f8a0e9cd08fbe96b9c049248733053a936eda9948ba61db903586b74e2d9e1dae3b32875beb0955711eb8e1eac5a99e740dbc8f78cbfda3f7a559049b78ac38829d87fea5762a413489b56e7bd23905d21fe1e5cd372a65f1b2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3fb57717b5da45991999058217d855809ee1f3f75cb56994cfe9fbbddd1186dab6f38075f23a5178d1f276f9b312eaa04d4b34c8c16a8224d4d7c5caa53295f66a7c364fa173dadb0aceb88581c69a8923c8cc7b25ae89c1ec05ece18f497daf89f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1585c0abe364b0804a2df5f1797c5860c8e8881ae1ffee38c9d5b5d132fa6ffc344bb71c414a92cfe8b8adf53b54b49658a6238b13bd25b2f1e8c96ab32f3eb9ffccf0a30d570ce645ec66cffc8a5ac7ba63b37a758718a9d7652c3e85df198e1a6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b46fdf1ba31795a903dc4bf38ec5caa51e86e6d634df0a1c859e792c68472a48422644452a7f065ea81d9797989649a5d72c43a3b73f99935f1e47fd1382696e12792f25b3460a395d5ab1a459eb3d870b2389adab16ef9a6ce85a7f04f135929fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd65a312b11363899bf45d4ff33ff4de8ac24d9aaae3fcc590cf3fd9c3938e067a038dce6de8a63b0607451c32fb543fd96e2d8b6b420524fda040bf5207ee86beb7648c294f52b31b122e24a07f03e9606c707104e17dca32e437cd5bd33db347b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb381bd3844f3c7d5655e7d5c54e0fbdb7e4ffd1c2b2e253fce7e769a96fe52eee8e0c3045cbb9f5443bdd7e81b2380d27d15a57a9e8e8c0129434d432f5125f4e0f6039aba4b16d650252aeb72f29563d005ef35e8e4ce5b5bd2400aabe1cb7dea9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h763387a38b669a23e5e221ecdb468510521eda35c2d2e03d91fc98b30b6e3dc65063b8ffee74ac1af4cf83317ecde332d06e58a5adb644384fb359666590738f9a83c49cde7e4e4883014fd156abc90dae32ad261a6973324a5a20d8a847918eb940;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0769ec47bf117627ec444845224f1769dbd9a8969b45793ad4643c08c323130a8a538666c391b2b94565917923e460015165ac3d49c7009abee14069517a90d9da3b6caebab16184a9ec8fcd167773c801f6933ecde40aaf3b864f42c3162792497;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb851dd72e58c0a03e66141c08221b88a1af33f6f9bbfa8f79d1801a4b0126d9ea2000d1af76f08363dc896f64bc576c6b156f9729fc1e4632b5895a3eb4a3c62bf959898d9608582ff73ab6fd5d2dacbfa6e4cfbb2ebaf8575c48db4ef11ebb4d28e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72dc38dcc360a90b1ebebd4b34b9c609ae37c795324220a9d9c82e7ef7e92b461af6ba1fed3d7d305c282dacea2615ca348f9b867d4b54f609839c114ddef177be6cdab7ee8b1d39c95556f698115b582a4fa97591a3b882ce1e90c1f20407b6b9d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8a97a0e902e18adcf640fc7dd5c19890447a6c9a8035e49787dcfdefaf8ea96fb4c1e96b6255eef0b3079c7e42aab1b5be608a96da69b99e2a1960794d9dacf1c1c09de51290e8d8b5406538ab2c1357b41c098ec34ed5c4ef33c89026b56fccc5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27db18a21d3ff54a3fa52ba396347b11e09ab25d3299899225d4a0aee898040abe6325a33350a963966d7a9a99bacac32cd3bbf555e25a51548369788cc312042bf024dec927fded11d0337c24c41295db6ba88f96af9deb350acaa8e9cd51b5a214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11863701ecc6c9aefb88c113152d4b76b6bc3daeb03e15d2040d4510ec3690cb0132878220b35a0ed9cf3e86f3c8e5d5feb1f2db3a8f93e67d0cd7d49690cd6cf4153d1aaebbc5e3fb94164804f77a02b56cc6d8fe2bd59dba400cd2685fe32d3900;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5938d85c454822c6abd977cf29271e811de7b797f87897f5af32be2fc0b602466e6bd3614b04e9b1ae9584dd3e4b3644773293ccce60da212569c714265cdfb32ee9167721e8519eda66b251cb688aded7b7f58e8ccb47d361b9382e9a38919497f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf07ef3021fa6d9ad789717628c9a8235910f408d9a29d938a1edc86195bf04fb099ad63a0f2e373c83b62df8bf56281e85e3aadfdbcc7ffc0e4a4c8c06961cef7bcc397efb3a37134df574336f7be877a40833b1d840ca2a2a297a3243cc25f9118;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcda35d10ab97a10805c67dc079a2e5f7950c19a260ad0a20f617fbc11c82aca078f37d92649943db3af865e773c00765c3572645bffb4e810b24134f923c607ef72a312d00d93ed3b172ecec63c74f77e77a41722ae062597fa6344b1e74a5e64fca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ecacf40e4ebaf75af7d9dfa43ef0b25a5beb39609af1f900382a476dd779bf1ce11dc82a47198a5d71707bfa697da49f1421b877b42fda0158bdfbea392c482127ec011860c5cfbaba75bec05f85e0017b0d078ac670f2232849805006a9af130a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h521f8ca437d9e8bf9c003b223de894e47605573c5a787beb73f382725830d381582539c7cba7fff5dbcc52b5af0600d42da97edd7c910da5b526157094fcd20a63b3bf1b03312c5456a810605ececf68bd8a424608d7f0eda20d96f93eca6990f49f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h967e46bee4353bd2711666b677dd702987242152ab6d3c7610caebca52261c6fa0f5a197a432b302521e466c94ff76bd0b175e7bf19e36e97a286987e26eb4eb86649beebcc797c989ace4e75a2d16ff7d4c10db02270af561a194526212e8aad6ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d60be1f300f9843f229edac67ec224d62e698f97f0dfdee35c002f2b6aafd9c5724a4d3817845d74e18148f147bb3edce6ce22a7185147590d378853918be2b6ecb094b1c8f73aba9ba662814f66bfb58174a688d92977db3f03461c098b4aab76a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18274a66ebdd53d04f293033a29fc710b4b7de94543d0a6b6d391a20311be5453f32a37fddc00391eb90b72782f6ebdadab5ab6960dd521b6262c3835ec6597b6ac0112a65977187e7529e67adf26f0dbd17c52da442011fcb5e59b4b873477db727;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99165a16cadc6114ade4d2bcd11969c505167086816c94b4a3cfca4f4c027dd079c2a05862b99b9e96a30440f35200d7ae166fcc02f65a48eb212d16e17b1ab47974fddb96654171677f27c52d727b77f0be4698754e0548efd29bb442d39ef2c2cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9173260c6d840c50d3ffdaa4b06ded5605d8b0b056a37579ebc5f3e284992c04057b0607992a23dbfeff4570e9e4a82c839b3d08c61e0fb99d7e70189b7bdb15a3489974cef6258e51a7aedf4d8b6295849c4a9639e2c4e7b47669464b080015a477;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33fff0861dadce62e8b7e1012a9fb872a925baa62b6ddd6855b7c34ef37e5637436eea8c30bc14e80dd5dd67d36205822cc49f9d9d7befa2236a56b8f99e7e7a0e4ab7dc4df9604f1a0c85eec257a7c2fc0f907b75e7a6edc1671f6138a3dd402035;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h582a024e9cafd24a262312679b888241581cf6bd5e8c91001bd0b0784c41c15c2a02434762323797cea1237e19c490f4c94166e5ea2f6bfccb49216a53d264b85ae86a4e960282fc8f0e095fad854d8f46818216179ad328b486064d16ba430a98c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24763f06dec25c4ebfbfc5736c044fd26824cd0cec8e204345ad91c8e185fe00e8bc057201e97afc8e503830529d600da661b2393e672865585dc0bc4e1361a31cea97fc156898ad82f007db28048f81b674658b2b715fa7907f058c03d9426d3f90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h766aa31d430e7cc5872fb5fefba1796a656a69d07e039e80fb8d38e0807b7e1defdc7df25fce8f217e15f86fb2e993de2c23c4fab17246f3e679295dc850646d2b27ccf1d943bd3e25e4c1e2ce73cece0343d8ec39b3980da591e6542954e4530cd2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf57efd5f97f14b5b2f2744d152b82e87613ad3391860c772c46a8b457773cdb07628c4f3344fdd95f07dca3a39f569eeef24a681ba34921247703b9f2f6f04e299d72702c1a52ff18bd624949ae55be931adf13847ff75f19d22a1836e249dfceeb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4f8b99685597eeb6e0c75f4c7c6eab5edb01444f794e288e9ca90cb1a1e5ad30c313a8f6afa19fc57a5a448d86b653a29ac717412264ca78f70cf6f0f27662dea75e595ca14a06e5f86013bd2b28019e548337e2c42ef3ac383f0ff7c3161c0e5db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cc3040a91f6d6b4d6c54c16b11fd719d350d547ffd9780ecc34e30a57ad62df43c5b5cf822bf473c1afe999dab6eb1e1c9cfb1ef5dd2b362c1a55843a64d77bc0c0610cfa6da6d9f9bb6cca1508ebdbe130f052cef1eb15e8f011e4676af7a26ca8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h542c929d41d97633d11eba523d734ef912d9347ad3250a6e66443984b3a873e47bb76c8909715f60976defc25b1476ac53acae4d8bd42462c50a92aa15ed5fb462ba1899029c99b10ed19d5c5cc10f8082533607263e77f15e547db2daaa51e7e873;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h843495ba4a601b01c02f235d8f4fab7e4583822af4e93e660708e240e52710aeaa39e5f1854715b3bdce0faee12bd57d97e831ebe3050189b091ee87f5b226337a8c40652cf3e2c6c6fdb10f8da038684176880923bd6d21500e2660301e6d0f534b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9846b36c40b4e0dced20500c6c3fd42cd222cbb6c4e38310f9bb9fceb48f14d3ec2878e607c586f39a40bace8edf760557184557b0c5a13707cefa6153656311968c6335314e0fecf20a4456f40ec5e780fd92f1c31316c3a6bcd07c3ac68286c58a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9440e688287aecd34444e2194ced8b1c59f49f9cdad6ced5ab74e8cec43e6c967e29f626b3585b25bd367d40ed2302d259647d293aff1afa8d06459de33430a25c7af4af509edd899172e195afcbd18cf4acd9cee04dec9515c5c1b471962a8ad7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8221592d961ac12d27649a3757435eebaad9b5eeae505c3b4e04615a35dd4f0d2999867e610bf8786f3cd054cec7104f38c36731252f25bb6ef56d6a0d9533e7dfb249699ea17f241993434be37768dcfd9d89693ffd525668b023ccbc0936e547b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87aebe1b471e769e9e4adcf5241ef437503e2e2d744769e610d1dfd0182b3df918cb326245da98d10eade2625de6871f231a8fb3d64c93689b4acaa541e64495599a191912488192b699041b5c00b0c2474d74fd0aa7f5c0d00652bdeb63721a3cdb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h392b2fdd162e2830b55d865441b6c91f5893624415e5c5aaf6d5354a6a80362b566d35d355bbb139dcb8c6569824f0fe5263d39bd5e6abb5e27943b3ab8fb5e97c88f11b4ac1f1bf21fa401c6ff06027c58de5e931f74d5860252a58db497b0e022;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f2c2dbc46092eff32427cfb3e9c2ba61598d5a8c65f85cbfc9c58e9472bbb9d03c51bc329f819dc78885145f3bacbf06bbdd2e7a4aac1277b18fbd034f1e22598fca3ff95369bc258488dc9a48ad2ca96e3c384a7533a18d0970412cca7deb696cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc75b42bd1a61089fd186b9661edd22f7743e951a1111e9d3cd6e5452e526d984a75928121b5117de819aed018b0c3d7afb997840f6f84b11ac447f19d2a25f2e0d72adf825d21a6c3c99c519aa7c4ca7ad4737196848b4fa2a49c38270334f38cfa7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6146750816eca8f10d7b39c57bb55a085fae7695a958f44525d411ffa0184a0a6e84c75f9e596c6bf9d33c3ae6473b095e0420e097bbe70654bbb9b0873cdf3bddce4ecc7106c9886c026b43000fa33fcad88ca9ff2f4036aa2073d03c24f826ba8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564a45f0e5bb3418e41b7ea5237bfaf0e44598c2776ed86569a34ae357e22d6758087b137e55c331df3241779105751a1274e9ce25712dd86877572e9d8ec521a2ee5e93d22f9260cacfc55464c5dab0c0428c53aaf8c1a2170dd2597bc67f90ce93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f198dc99084503e51641cab6df491dc564afd7de36911843381bd967dde6842a5f62835fcde957cb69427dbdc8d3ce498d4fda1fa9dfdb85bb8134df17da20ce4cc198cfc1d34cc0be2b0bb8376f95a5d3fe07dcb26131ed151f6329ca7f780a4d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6abaf66b14fb8aa864ca075c2fea58e063c956cebe0e5745a452aec9ef55bd4aba33d9633bc103c57f2e6a6c52db0887cd8e9869d35eaed6993825c3258dfa762d4e0e1f63280c7cd6c639885112a20a303e9a9ed634d7f4ee18986c9919099f0857;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17013b709ed4a79d03f696e702f10d8547c6b63bf0bceb0d5d41849a77156893e11e8a2943cade1ad7f3fa5540b7d70542be3179a78fc97b1a28c3a7b8b341e49e1b6642bdecb17df51f9efd44471d238d24266921169377e7d2d6677419d202591e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h157c3b2e438296aec5115f97fadd3f317dd5e2066a0555a18728a20ea5c80becb4a0432d315c5a7325d4a353bd8b0a024f43c12fd79e46df152b97949fe233331c5209036e6b54ff8cb70968f1d754f04f7234bf14af0ee7675b17994d5173f5b199;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha75d7bec5a89ae18a186b85874db9b238a5b254722aa9275122c0c0c3dc94e77b7d14b5c2bafa8396b998896c112a20437e816bf43d3afc4f68f4892d6acfb75714a202ea9edda1f5dd04330117fda546088def74786f54548552e2b537e1a31d0af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1637baa8ab160efe5901d7a7b5b8ce63d6d557912683514b1216d83fdbe020902db629583a9215d6e83d6e873e3d85fa0589d12c3cbe9c80499eb6234e276b21dd6f262e502078d08cc0c82888e455b0d86d6919f12c539e155bd0afdcaddc0d2a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57600268e1bb59c688911c570fe6d19c7f539f7344f78d62d497fc09b5231a587941ec1b505db2a165c7ca78e04e39d548299f0b9f16a11232450a9a3d3f58f4075d9825bab08b8bc3de8549a27de52c8c8875232a7b7db06bea2b47a1bfd6576f31;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc646f59063e0a87e62bca7675975b9075c4af9b73d09e805c6ea35b62f110f8788bb526496d88860602cd4ab8db7b500d87dfbfbb264260a0d85786303c104d9148b85b572a59618249f39f5e9c7a6c974a1438725bd33463cf23deb3675fa345223;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h894f435e94d9a79be1a8859529ec4c32d2563bc51af53324cd0a5bec85be966728022659cd268ec9c6da33bb5c6c8ca25626c279c8f59015cbf9c5adffbf36dc8893042458e8870c16242fff272e3065ee3af447b96367c186c0eb011e3e0dac3b30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aa870ea4fc44696b677f685b30a6c6c2ed12a05bd631d3c2c8c8092cbf5e5f2e7c63f354c085e745a3b874688f453d74bf948f2403aa96d29323405f265cd7cc203125ad4ed2785f7bc6a9778d5bbdbffcfcb29a1afcc2cda6cfc8aa7bb7fa82dc4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ec8a46391815f5bc71cc56b9c16c3cc4d29fb0e204cbd445ef04ef3492363ec3c11d898bcb7534489c62c713817b0593042cf07438742d79966cae507ead990eea39ae65c1ccbeb161926e42daba8e13c3610f26948a419a9bafbaf70af35c6024b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4097115da6d28541d94fdc50d38ec21160c3de5e5120dd030ba2364f232fcf0d40530910d2376aeb6e4f68d12c26aec38dfba2dd9589147b67a1a720f05071810d20172fdb2119093a701bd7f058e44220d88e26864fe74e5ce743db473a166e69f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65e721e156ffb4f10bc9dde0988332fdcc06c2b15c4a2f2b8c14facfc2333b509c668e7565e3c00e79d22cb66f1d6cc54606c4dbc212c8918bec5fe27bb569b3339c28eda62d005de6bedfd1fed42569c5585df8038fe95b5c70476751a026c4193f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ecc28a383e9cb2e0cd8c39a87650fd25e8f22bc1391c40604da60ab60c96be232888ae13bf5bfe6de587df83b47355c7226c9c2e68f7022b75f1500cfb5a88ad47b45dd9c36666790dfebd7f4b6a232052e85964c3ea313579421ca5b30e2c8a7e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d959db048441c5bdfce008271a48c55e10cc1c557ffda56aea6abe4934cd6f4a02cec989e2b3f1d24ceccb7c511c08afe918d2306933a02c192d441acc6eee72ff5ee7afeb56a578af37bbc29ce1aa02d43f32b4f2148099c16b84b8fdb55e65de5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h658ffa235f8e11bcaa89568acf34d09f3f1adabab796ad90289fe0e23dffcd2123ee2f6e6eaacbfb1421ee862986c0d71305eb502a5f231cd9c7afc0d08ba3f05ffa5b49788aea4493ac30e9a3e7aec6275889181fc844f50341067ac2dca36bfeb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h720408433a215d65036461e3d4cb6a8e6cebeb24892ad2989845da871a7b64c822614a4931baa1adeb37ea9e7485ee5ffb76af827e1d364a56b787efe14c1ed0b31bb3c5576e250a6d2a9aa020210803ff84d17ead3228be280e9d78b415154c61b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8c0ab79a2d76509725ac312fe60c327a31e47d3a1d9899d875febfc40c44eb2d8a4361e047b57370622019dae6b0fdf67525b30c5bd199a0983bdfc6ff1f3e64ad23a6d6b4d58ee133b254243c7ab6fc89a873c1c72ca10e0210241ebc6a2fd6010;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a409a740c03c5384e08c441466e0646560d7c57c68f0214694ea492cb75ce27ecfc3bc132bcab8ee97903394b1c188ff5481db34b4780eaa68e45752b1456355715c249de8f86e8ac90a77eb29ad45997e07cdb740861be5ac3165ecbd8db4d1c16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fdf62adfac814e41b5864de654eb67f2bb3f6f00968241073e36009bbac9f442d3c78562b00d40dd3f23fae4f5c2199b4048358ffb29925f4eab3abd1b0c6bf4bddf3888445df3507120577192136f22714911dee100530c814e1d0f8acf160eb49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6abf787e3d22c76e979ca0a1461fe34ba5b06832ad6935fdbf2466a462da7f50a33555a83b8a70a8f6a1a101badc159404e5a560b934a661fb523ac7c8171e393860f939b19ffbf0375578b89a63af79e2bd1185d38b1afbd15196cbcb8dcf2dace;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h206a6b07216516622f78bb861bcd653d885199f4cf96ebeeb1908a5ffd3da3fece9324dca0de8a3dcccbb74c48a590bec58f362838ce4ba53bb2c644a22b7724cc0cce2b72fcab101ed6678bdd0f5b4ad71f018f4b871f9aa3bc2afd98c75071f911;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18d78ec395c52a8d0facd9369278e9bd0c90b31ce35eee46d30e581dc66edcce5dc2e878f1097878052986b4137d76d0729e637f60817b08bbfe283335f11b134480108429eecb6b49d88c03550d827463ad94c2136395b3df9d5567b5e4d89f7363;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66264924259b5c2a0857cbcca575ebc704ce5319f8e938cb6f43a5e85d804822859126a14893dd12f1fa471f68fe03e6847fd1d58c74530d84a65d5cef26cf62568627d84cf5299fc3380871f97a60e75c8a63f418b10742e28bbdaa627a3cf2ef3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0a3ed1e00a6f073d20648664e73f6a70115e08f9f8fa77fa4afc9d75ad8fd954c4d88f01c7fc47cdd7851e03f4bff989e3a2bbf9b098dd05daf731d884b16bfa91e0d69889cf09b10fd3c49bc4f7a5cb6e3ceec5471907b3f7ebb0c2d9ac2e60f1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4aeef83a7357d4080809128d210fd51c54cdaa104e0d0382d7fbb01d97b2afc24fc2597ba508ebf2e1f2d429c50d2b722d24b5848941ee1fd8e6de872da4bd71bc25b9b4d4fb55c6b6ac24767acc0255fdc58e15519a5f29e6697e5d20fa761c148;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba82bc7774d0002b2d41679d36b287640e3b2b96ea992846de2b21060f20a20c122da6fdca7819519ad245accf2c9db3b368b26dfba4482c1c728b4217f1f1723ef495c47d6abdae4a1b166f31e3829c8a0648d681021c285bc4df898613f640b391;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab34d4cf42292fb8b68e0adaf1207d6030e9a104a98adeea3edb15be7470e4a2800ee44c9c121499953dfeb8045ce4be5d710e5e7e956bec58ac49f550d358d1d88bbbccf51218f67fc3c968096d1c4f84d3b15a3949863dbb90bbd6b7dfd238f92e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h345b2897ec1d62a17672d14e38b1fc3090fd502b8084be91842e4e7dd2d4fd4e564076c76a3cb737ab5fff6cc8fb5ff24ecd50bff1c1918eeedef39d4da8c1cfa3dbeb761cdb43974af42e4a5d3381fef51dc51afeecb45558bfcda7ed837fc4cb87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb47260f13c88adadf4b52fb7ff4da4694c2c530a6210b3fdd7516f365d7d301f6e9f48eb7b2d07040f5eb22b98b3f73779ca4ef7ca7e880cc135ad9d05e2b471da3c80a6023923fceb56914a15bfa487d139b10f0f72f74fef2122e5cf3b61625992;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d9ce3fa8874d766fe7c7a001b013566ea2f4c68829bbdfebc671724a0a3a65bc21f75a8648d2da98406b7f249a7d850af4d22efd03be77a9eb7fc9a5836cf3bba7065ebabe24f02a4734244d4cbb7148b3d87e18a9f70d81745c95d95309b9ac9b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf9ebf090f5fafb55bf7186e40d6f26e9118fe134fa4c84e0711b82e61e474f9891369040bffcd59d08be62e6485587184f0bbc88a007f7ccf0c82c4e9410d1269f892076970b9af235a3fd216a06f765a4ef695e5d50c3f41e6d54f34f635b68315;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e748ad15f2b3ed41ddf05d07c1acda2d30c5bc6d0e60a61e654a1897a763677100fa86c2c58ed525acabb617c4d51cce867822be6ff7999749044ad20fdd37a0fdad716daaada77426c3fb204e337ba1983b8ccc2ed02c7b2c0cda8dfeb7e46a1b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a89abf2065af7238ba4f14ff09b071759eaacc97b3cb64f2d6e82e546247b9570ba0019ed7a0cd3a3a168d752a3390f88dee634dc4e6b32c62ca6dcf062d354b6363b1d2abda53683b301cb69338ecddac2f188ac0a8115b19e6594b031ae1ffee5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d9a65a00bb741bf71f0fd0e681411841290fb98f41c8796aad46ede71486aacdfa2563b51fc2879b348f5c3aa69e1045ce19e8f303850e0eed5f49e5422152f10cc69c46e65af479185e2c3f36d5074db7a155ed1d6e36a016775de80d6a4f5cb18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a09f8693918ef92e3cf2b195f08d2d675c64a31ecfb2da7d2f01143f0d4741690c59bf0bcbdbd2c36bb60dbba4fe9436e505e0dad56a1014f80a8a2aea4eddc4fef9fd6fb8251b29282cb61ac4d8d94db29ebcb34b935d9f4733a48157c9dddc703;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae7a8c51e1078eeb132fc820db30ab649c9570374fbba3be3302848257a19babe475baac852ecfa00cd95b918154f2d3735496b6550ed2fd319d360458b07b477a5543c689b2d6145f43d13417d2c60db7e63136ee18ae841aa139dd243ccd406ec9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3b34c0038fcea78277cf86280b916ea1d8086b06359aba43e791da4c61db1fc10328872a8e73190f6a9ceb39ddeba167e7461ed1461fb9a8b0dab30620583c3844b2edb2ee0acccd4adfbd5221d690690d966efe3d36f33f0066b040eca0bb20be4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9738c36ef9125805f3aed27bf4698080d350af0c7beb5b71cbdd36588f75a5c2135d178ff0637bdd69fe8f813c8bb3f06aa609ed77be271a7b826b8c5aa373a09dbb12cb53fca58bdf42a6f0d8fe5721d3f7c88d37998116bc1d5a2437743966a676;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h697e7d0377530508cd3d6f41df49aabf4f3ff13e391d58322a09f863f34e297bc3f0c31710c158b780255d6e6153e10928776e08ac4e883e543e813269f9af48611d138246a47fdfec82a0b6cc71bbc91911367056e3184fd3d56f342acc3a78e87c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60a4ff9cd820250b907170800a2b9a7f24be626369ce13af7484f00f69d63e07df20552fba8f4cd5b3dd107af12eaeaec24692159de97dc9f9e1e193428d7e19f7b6b638441019a2e0da915804ceb888bd849c6323f056a4c113914703e6be837e61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cecaf753d590a9c21046d1de898e427b25a647e74d75a0a5259ba3d22d78cc92087ccaf90109af300100edbe9ed2f6dc7faed3e7e9b15db6659a3367d3fc90c1fe5bd6e6482c3beefc95f712230a868132521a8095370f284a0669aea74be1e3762;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb6196c3e1198599ecb178f81793663d3922b3f52874b69bd19c5490df94cc61aa109e4576fb533d6b9dae69e68fc9ddb028f654c352d88ed0459db4000d1008f24eb8b4299af21113a49842e591b252ae26f989f5d7d97139fdfc457ec9883008d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93328b1c932455197434ca4f8f7a9c92b059c36e1a178075c2a1cf2187bd96826a2843ed2eecd6e0e0499aa8057f8d42a43b4121be5831233d625cda6c5e5903548908cd02f5ef711090b00211a21e7e651d500ef651de22d9f8f9658b8f2ad9f4cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca74a218bc7a79623d3e3c78af70aa487c6e195823643dc8b11cd0ee996850c08c2dafb20892ed1b05bc1a85eff301a54494caa787a4160477fc9cd0365471e620127ad7eebdf94bdae39177c571127792e0f59add582de42c40a56277d33350e422;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2abe5df8eb14bc239b42ca20e4c930fd77cf12f6e44d2d1075d70495b3a2074d00861b41e70cd5d704dc814ad69bb2ada7e1912f43f7f45c4e8f8872548c1229accb1aaf7921b7aed20f30436ba4239de3c17cc9c62118b436b87d33178f1f68ba30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e808eeef523f062ce89c1f8f4d92fb5f18dd53ea20c40216be5a8b979a14b706c5a4029d2d3929b7714449a0003b888bb493e27a67dfa27a179e82396cfe84257f34d4ebbc7d9284eb76d82694b704d74e1065f771a41d162c49f6f36438008e30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb38bcf94972ec39cbbae66dfe171d58ccd35d624debe5b3c037bab3639e6798bb78641a8514f42203fffd556c0977cfd0df71f65e8652c2dd6dbe2de1d97d9c340b6188afe7fe64618f03e8221684ebb61eac4fc9b4744c6b8946fb1620e753343bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3e593912bdb6865cb616cd32d578c5f34a4b0fc1368456c49ebf46f5af1b595d14c3e3004e674a34dceb4e83d9392789c9f1387d045183e8bdff56ef29017124abeb4ce4553e50890c393662cc85d263113369b08ded21701c2881866670bd997c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4f1bd9d6004cc67636d6215ee3d4e3b29c802e7bc1047ea4cd6a936096ad80d7a6f176a2851f03481a7fd7af0cb92f427dd6bab8106de87e0a99d3945a7fd99d62b4f1cc27c8f5fd6bd83527f7515239a63d984f4a8340e0886349a20b4ab40f6a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha546cef18ec3a303c9cb3ff33ffbaf0fba454fa9a9d18e07377d3cf6cc53d33f84fa90862e191d85ddb37ad00803644ead14fbe6d14376e6677865c6d96458dbc5cb98dba1dadef55eeb2118959d25cf1aaaafafcc0f1e91d202b25d86e5f4a488c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1da2bd13464f494c62cd6678b9f474d05ee7e49fade128445a8b5e71ca446ba4cc7d279d958d2fb0773c70db9b80020d494b42850037707ea0145fa6451ebdbd07237df5c6a3bda56d89ea4191515a4e47a538973d3e36f17c50ac762ce464fb2b02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c2aac16bb3cabbe0ecf55fd7458f3ae7dbec934f437cbbfa7fdb333af604a36e8d3f4dd26b375a5d5108a0cad1860fc25434170aa7745818388a0aa2a62046bd3eed8b24ef126468ced95f90d35cd762084778ff2911ab7941d29006f9edccf169d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85395a1cb3655cafc1a5d70fc8fa1c7aa0d6ba902bf24e5401080a278ccfd35d6fee130308089a1021be19773a36cde4d8ff8164f2bae631a2387a63da58293b2c260895770df70ebbbd3f9e70f89992aa19de91ae78bc924f77d1364317b53c37dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3df88e1dba4513c497eb51bbbbf0598f152c2a445e3ef7f1c2542b63579bd3215b6c632ebb494899f239bb856b4736c54b6529de2bf11d14382c884cb5dc06046a1148dfa6f550f106c1e3c30daa4855a3a80ef620f28ec2a0ff16144bf454455f8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bd50788a489c7f595d4b79b2fff29d58dffbe4fa4c6789022ebf15559c53a109f3189ba3d5e1ddf9f36810493f313599e46221ed167085b2bb63b5f945ccad684147f05ecceb65d7d9293f65b7cccf059808a2328cce4db776ffa8a5f36ff1cba8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h468fab88d2d139bbbdd4c071d4920f14e97ab527076e6ff9d291c903d7514cb4fa986330cf8df2bd0b79d0256f2f0f481504cf34cd24c14cfbea99bfbdbcba550878f42fdb5d54bec331b1c35c987fa209300df1ab4155a713412ac284c77fd5a3c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcef35d2e218843ec0034da78a814f099c153e8b9e785c4aad4163c191aefd1bddd7b2ec83b8d8c6fc06bf3a701e7fef500c1072f80f3f1c22dc29daaa62ed770e276c9b61db10f8eb199aeffb839ce8cbcb67102059ebfc2069df12b04669cb52ca4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1574da4a434c4ad9225c2f19b27f94008a8c226a0c7409b5fa4c0d0fb1356944ea15b9dd809561fd0cb1b6833309529a721172201bc0126dcead08c835e40133857479bf197077b3ace51a8696ade644cacae50d8a4390651a473ef0fd1056b73b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec6b227cede3d2f97e6e7bf2d8b7d3674df27596187d51550dbcac4ec1b8a9923e43d13e89e7cf17497d0046d5b8ee724a8599db60947932f7cd8d9b5dfad71760ac1d0e4abc2847a8ecfc9061b5590c40550cfb10b1c8180269f3222da4fd23e832;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9d9257f68d4d105cd2a18ee10477bd974634e03b9b361c2b87a26457f9b60095dc81d7d7f40ce6f41b3aed0e22b6812560a9a5dca0e8a05e42d8dbc892df333cd2b2b23ca9e49dca19c25052b29dc69eda70772a01771e050c2dd79f34b8c4ff48a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h945182ca7c102352b4cd58cae0aa471673171ea1c6151b207f126f593304441eb7af1993b4e23005f6d2dbca5b4b3f67934dc9e7d0d64eebc714f9a2e425f761fe122b34ba6e9beb64fb87b22fee5664bd878a89000c03cbbc1067ac8178f0f2e602;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9345afbf65ee97a7452c56c9f8522161fe3230f2e785ecdfbe339145771938b678ac18076d3029ea650058bb4a20308f205e90fd00d9c27dc65267a8e172f257315ccf63531146de9f6b2e9edea6dd8f7fc81e06b8cf2836e61cfd69399d5b6a9212;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdaf65ee61f9dff758cd9b13d1a793052282ab1eeba0497c5f514ebd327515324d8d76415c51a808fe2d158c800a267f4958044570200961a17b70f57d26fb8f5c0e15fe61944c519e914f15257fede5d8cbf03d5bcc2801e7270cb3ec60c1f8f5dac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91e8dd11c70cc9c9ce91d809d945b5c4556dcaf77be770c61a46458813e80318af6f0a911c786992bd299616eb1bb115817e2e58a057bd8ed303ebd3611018c69624b9fd47cb14ccfd5192061b3e7b09ef645690f1c9d574e58aa4622851bde9a60d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81c37c9a6f0cd2eb0344380ca6f07913b1fc5e966eb7bfd93f84a2b97bb395ff2986b1856c39fb3e6acf6ac0ce9d4cbf33329e6dcc669b6da7adb70ff68b1dc59694f351ec2dab8c718a2a246ab07c398e1905d4ab512f60813682d197b70cb11081;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb439a89d722bacdd13f16595ad6dd764c0be5530b56bb5205eae230402ee895cc354ed3b6ccc38ce8c48023f50c8d6fe593d07afe5a05f31f31c510d5a20d94683ed5685e2a9ce99b9461dfe59c4674d0eac820b644a63ab83e99f56db6f7bd9277a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62965abc4a54260a330624ed9d76f3ca90bdacdc82cc5a4c54844c120c10e74ed259403cea5dd3dd46b11acf542bc3e21ba21c2e92d9c871858c9aba1e5c3208cb54b4647eedfb152bf1379d4cb16cf852aad53c37765c991be17ef91a7e1d65b134;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34c4f9e38646cb869a12d63c1c44e44749779bc8a62865b5b842a1c5d4fa5a3e0ab18e72b4303c65c3d76b423f84afd991a2d1d1de66d0149b0b6f467955fc3c4dfa26a225f11da5c901ae3e670093c2c0910b9035931443fc98d2f6e61b85ca79ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a827422dc3b517520002ba35014f7f7de780707066825e7826fb5ffaf3766ed6027908e84746d43bf0be2bbd763a5a6d0a8a8aaf45b1750e2324009e0abcf7d9acbf9a8b49b690e827b9e16243c322a6aaadc5c3c82a81517ef449fa6186f7fd34a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6a30ac2c2ba2c0d72454093f78230ba5fdcb15b213174b20452a99f96908fe96677a1d78c47b79862c3b15ea0236cd6fe97bb6d2ec0f3ff834c0c6c1e843fcf853b589845c7512032804026e1a9e77ff5bafd7dbdce52f7029748ab6580a313608a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf98a20f80b0ba839b89aa94071d03917eda4a832b12e72c0dacf06c90f973b614be27fab96b73130d905a32a12764e8f44d57fc933e4243d900f5599fd5470472529eb1a97cac09287b20df55e845f90556fb00f7b70807b9c019e505f78272f6773;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee7355e248d76b85040e21f8367f2724015568e2ea7ffc5a72f114102887280fef2cef686cd1db692a0dd68d048991a9185417975c195ee3b71b3a8aefddaf71a54719cedc6d7893811932e827a3c13efb92e8706fe85ae295d2c317dfe3f55f91e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1906d786b2be20105687bd9a4c3b8c19068402bcb7e14e0726f1f8bf56079e581c12d6cd0fda3a305c77076069ac7a42240f15b067075ae7b72cc043ed1fe6995a1f555547bf4e4e1356520a5e3e862c696b6918c4def9ad534352e8958ea6106a4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h105fa3454d4a8392cd99298124dbd026d73caceb6f97c819ef70e4dbfaf8e8841eac86ea5fcf90093458aca36722ba5af23bd8a37414add047dcfd6bc75db0ad0670ce472a8bb879b12e19aa713ec8f699dd2289d2eb4ccfdc8234c1aa3e7dd54556;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca8c5ee2d13c882d411a4ca3135d8eb67718f844147db092a37f21dddaba5bf47da3e51c72a128a4594dd800fdd486e396bba6341b5a6f953f1a4f2eace0e826fcd0354178ad569dcee59321ac47d1920fae7477e2ab3317d11fd3e25de4e23ce4df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h731f25c0b2554c3ed0a402f6800b4a7e43fd65f80037d7695c30f0fb0c48b084f6e39be0187da3119e65c0ac8ec96c787004c3e823efec06235073432d7c79cdf319ed3656080eb3729a94048c6234ae2a728e4f8e7170ed0f63e4faec931576376;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b0371d8b69f2fb1fcac55520d370beca9ad0f77a83dfbf2e2dde1c59f577ad73c9919aec3cd16b0f34fcee0d02a35045a4d764ebe231a853267ede8e4c48a710ed804352bafdce891adf436646a56fef2644f647ba91805eea97e33e8c36988b1b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha793b16a1d63842637d99093e56efb85e2390954ebffb29e075166853a3a493f3829a6f4872c1527e492233ea230a50ae66b454ec8e5c9a80934916b8180a384bb49f7465813e56c54178993eb77f4c3302efac2759e6102a3dc0eff0501502347d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacaba7df86a0d603bc332059d8c7c4ebf9c54ad23a0453f0d188400e99deda8ed8ed174959ccb1993202f1f05a6566af4e9fd88074e2f75d248bc4d7706a65172cb88997aa11cb1cfb78f0f086313af0cf7224e5fc2d0bfa063755e45694981a09a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ce286690cb26770ff8b68d7a8074c9b39d591f808bbe323d1869fa2cdb479456a17aeeed64c61e9ff30eef8d6497eced6f1339001c5dc56eb4ec80f0b953371fcc0821bede61fffb05ce7723ce55aee58c7054de063b86fbc3cd9f25269b751224;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8283a1c0d36a2166ef2077be66eca35e217bece0325f9db88ed06315bd10f56bd52beb552fcda21c593d2d44c8e17de4d1dbdf450c91ca9b638b30967f90ecfff11a41aeb8d0313f0eec26c626db862d5f5e1a94939ffc0da125f56bf69e5f6e54c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8caa564dcd6d49890083cbcdcaa0c4d66701666555284b35d4e0ae6f3f864e6febe11aa1742d56584d61714f2f8ac1bec89de61f366329e55d8ff467e3d254ae1511f64e4a4caac183c4ced350c5f733033fa428743e3e253f9991205ee37f817dd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95386db074f44edf513ded5eab78992f9b3262f5227c4f4b28dc2dbc18f451f37eb1a890102ef192b80762da09f11ef1b18e072e6ef56f283bdbe0a7310ebd734dd2c1a589668c37aeb6f0b8b5f235113e2f6ff5b8178680c335a44e4cb2457796c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdea0fd9f9e334b6550236024fdc6dc3688e7c63fb2a79492aee67ea957e82a0c781f83c291c0ef7d25929f2a69723e25d8a160978d1562e7e3c6b2fef16636ad5fb3aa0c674719c04be6014c914377a2cc1121f558e42dc4ef9a6703af31d616973;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26e5040167d10d9176b22e7e2fd815dd18df1d24010c8a6a456b5b1613db1927caf4d8d61ef760a7456a12aab8258f2a22da94c74d86c6c9b12fa936f99520a6c77cdb31d963ac4237f6f4ae5766af913a55ffb100bfeae30b768d49ede89eb0230e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46535794a5dab7637629798315e81a3924a989d3bb013782cfca7258a2e88c3b8cfb35634a75656567e514190f866cf23d6c8b888fc5f851fec07b5a87cd586e1ca30480ffd8728dbbf164242def1dd0d4b8c7306e0decf6b7118665a1aaad9022cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6358c7f08920b6c146d4ce1a12fbfc3f614ed74a7b817f2af2297482e200ed7a5f0c5da29b5e2cb91921bac1d2265264735d133bdf37fc26a72eb0ba4e2afbb5cacca3494c083d6361ffb3d6cc301969f3a69d460b9c616213ff39be4221f285647;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc697bc427cec0bd62e0fc4388741b7507267724c1e32ccd98abfc6fb4dd6037e057f92154b6efcf81d6f0d286300ffd49fdf563b94789202b268ee13051d823706a825df787f5063e3a58d48d174f47dd616782e64691b53d71fbb497fc04914a8bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he00aa8348ee4bf6957be09dc0950b21df79823ebab7c3c2ad29931c7ceb3b349fe243863c0a0a1c4ca0755759854719d12d64860136d77ecae3727ddf5d3d9c73d4c4059b2cced11289aaeb0b768d33f9561538b0abdad9a107ec0da942a02ca6332;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27412fe722e1b27de13e261d327a8a3fe57ab15c9d8128f10724df59a3cdab09e7f4d2c916dff9a76951b06de0cbf7df5c1506cc0942494fd971ad597ca118e3594dbe4dab65463665ae6991fb4b335d5a7d34349ef97ec08b5e5d42dfeda3d102a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h168b359dbdb876dee032aa5a6093aeef9ae759ec4ffec4226a0f411e17267c645f691cc6e0953e1bced0d8d90a2907a0278a63cb35b545ec4240d4d7c61ecdd3f2bf50f31ec47d8728aedd639a4a8377ad0d14fe300a64ae304c03d49a40ea01246c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63bb49e06cfcaaad6581a1f09b5c2f22795c65d5c3abe01f1fe8a30ce0eb910b01b741f71b86964ba49026e8d97ee5aa1c37cb1681ad1974c8778e57a50a8261a34c1314e66870e809d696b5465214b80133498cbdc16cfade3c632dbcd0fe50b753;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6422a68fff74f1f92a90204dde4385e02cddddca606b84b345b67a1fec19aa2b0e7a60913502625f218d1d1d7b1f7c435d2e0e7cfcf9a09da6689f80261ad7494d07442e0d7e923ecb0ba9d647ed53cc26e7c998404e555ca253f3ae0bb657c1dd11;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h817a4367ea658a50e994ba8130a5452812be11db8e6f85456b038594ea3f167af8029db589d71986646741a3a8b6b5e52046d9f578fe7386447108fef24cf2158c59b45c85c128ac6cdc300de71311388191fa8b394a83fb189c443cd24fd0f79893;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4271879919a9016e1b78085dea2eb2c26c4f26f1b26b3a1372ad04a5d0f64d7bd205968aeb66ffed387d8c4ff9a49385f54e93cc2725cd944bf326cb7bedfbdab57ad65cc1f61ad36d76a39f104ad3b343f004b459a0d78ea761729a6fd0be2b0580;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha29ef088df9d65885955b758c564835c06236da9235f9c254190bdf64755147cf7893fa2e5d36191e06b359366630113edc047bf0e28fe0b25d9df1480685422611d946de0f5b7cae6a1205970a60e5aab06473f2353d7413bed03526e23d2ef90e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6eadcbd5e17cd24145a7da2aa08121598adc24eb928b468137fb1c5a404f48b7505f5cf5eedd11eb51801a5b09a7b1ce45ecdcd7c61fcf220b0f5f9477a2da1a9304c780d949bc67cc68771094e1a871bf55aaf13eeb53951eced99a7ca3e2a376b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h316fd4373594acf7f10c81122a0db5a5f7ab61407ee6154de7dfab9e4063e57d240eb86b5f087bea9cbec756d45e894aded15d6b9d126250db8fd62490273890d8ea8be362b9c4272c1e9b5faea5edec4d48c7979abe2b462001820234a722b255be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc4c8b3910667360849cd781e23dab8f08db6398e4e0d40fd48989a50242a7d21fa8ec1159cb2545e291eec332d8e78666399c64ef3387db01522b5e22130f9fbb59c1bffc3e3a30d1081edbf97ab58d2504d89c4bbd5838eb868c5d80a0d9a8b812;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdca7c2a863f367042deb95ef084a197f562f8172c8e54139de4f24a140b91498ddd14ae5ed68827613f58bf39dd7391788b4a3ff5242d10cc017a6c838ffb0525aa4368d2e16fbcca9c687df4d41e2b6e27529e8cd5c351365726c97e7bc700723b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc08a6768d05c37c9b275e974cfc25bdb1b51c82655377870bb242ff6cbe373ce66a236836566345f8777a0d7cb3657ff9257a65639758ea0dfda2d59134c9676dc407f1994d3b603fc0827dbb297750731f11f3e0ce84d54e7539705346122497fcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84baeca084801f90f31ba5173a112d48d07c0e168e889939b012b129e9ddeb00df696d751ec7433f345a554eb95568e0c1d45f135a4f1176b35912d1aae2860972eaffcc538df3fc04f0f7ddd390645c35259b55ba325fe7431a724416e7422f0f19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3d136c800438f071f7f44917567ffea6019c1a6a97575558362d066a05d5586a3081f79afceb802fa3aa570597c2f79c849aa3da922fc8a5723abecbb90bf090cf875168a1ffdee2d8eb37e6a2bd9864de64292f4f10bb88739c2703e6ec99ec727;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd49fb8451d0cf311bc00d5b045049163cccb5d9eb608e0cee63db960e28517c4a5346e61ba115ef55a8f6d10085ef780c01a63a71db4119df551e22c41a75da18260fe4fb91888e1c43ad935ca224528ced78161eae9619ad860c5094f6d53c6b4e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a74bf50d421009ead29f10e8aebeacc7caa62a72064cf80a7cc8f22cdfa161632fb4e89b3626ea86f15cab497ed0b2267579974bd715391bc76cd6ac36d4fce57ecaa190b2193c2c6736fa75d38ee4cfac4851bf222326a829b337889680459c22a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ff11eb2792f10aa48cca0f6947a7bb32f59b953d86b7846a5ff0c7c209788188dea6a1c0398d910da6537104d05bb64ffe5b70c1c2bab4fd1bf5dd25cf395c21478d2e7164a12a3b16b2900e0ab1c280ceb5ed54ef6db8c49de8bd6da774f1c5763;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13ef6fda6fc0e6869cf94e3c3e8564d7193f65d460715dafe5758daffbeef30349e025fc3b9d521e47d4147e0beae5a87cea4c4e7884c609960ea73cdf20edecc215fe0673f2d2e4259e3a46e05b7836c32d5f46791349980921f43a701b54b5e98f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38eb082ca729bb612a9666634419b01d14cb699fca07c18a6b7196860d50e541df492d9e49ac7484b89f6766fc245f3947562c76a26ac80ea91a728c68e577a188f6679bd4f33d3524cc0b2661d55fa38493077247b409e99e3d7fd5ccdc95599f27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10f436f23c5ce526b5370d2d57f876a1bc1db85f6b584ecbfd3c83bce57dedd8a30f52f0ca25a6c003565bd78f8a5b72cbf62740f63dba91062fc9bf971ffb5c697f75fdcadebc2031e318ca8e52c39a7f16972fb930dc24a5e8f5bf1be4be24fd52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2588654a950aa5ed589ddcd25d503e5debc56f2f13cf766f745d3f53a3fb9e1ba083533bbe890da03128eab2e6ccd6cf91cded511b1a307e2bb0ff6cb8e44721985f6644f6386a0571f6c6f2831b72d7af45ee26a999a2107a97bd7cc925d8dacc8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22621428f6abb189bea9b5dd8f553bcb826cfcaa9c5361ce2ce443b58b69e122f8f89ff07dbca31fd0b11580b7ce83e8b6fd73017e4baa9434b7b46dd15fbc2ccf5f56db33fcaeeffe3574d3c19a6c35a5e06e3a6acb36d45993119be8491555f983;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ed1295a728eda6a5d6765388c64c77215e87ab5fd8a2c15d48d38b626c6af2bc92164bb0141c073c1eeddbafa20cf1679149b923648225ded9fce82666c396ff513fb07f4ffcfa50331e91dab53f07ea2360783c409101539b7fcd0825d3da40dba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81f7c168b0e25b4012cc3abf468dce82cca959fa1abe5b485f1271324f97b3024e671d62ba64bb7fb3329a92cc5a3d050ccf1eb7b01fe42cf343dab7d5f41e138a9138acd610f304d1a008b6388a6c4affb4c1b857a45b2a54a931d388c34e5baca6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d787bfcdfbf246f708240dd25b6dbd4a5c8f7187c53f6e1b96f77510b833476485d24de8730bfd1646e7c66a736e376872512b9bb3fa636b2a12b06561b6096d6b8c1f12e4a5f44c01fabbb0e3c5a46c30984b4c84e0aa710f1a6cc5bbe24cd6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6dd5f0beb587267078e4b1c7ede10f430d9bd863de0c1582a4f411310c973f86bb21eafb6572e3474945e289763ec414c16b287772a994cf4282f0488fde551eb71ab796852a8c7681e965f65ef1c0b5bd31c0dfa564a4755db8b5267a3b2e4039d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he987f7686c2001d0411e617e0a8b7b434112d806f5c9e9e5cb19ac6449ce4f6fbe05ad2cfa66a59085a17ef534ff9e4019a78aa631dcb50746720f1b74755ae18b3866f81cb05d140253de55a8a06e7cd516a925f750535bd118959b4e33292d57c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h745aed56983eb6dc6f73a79af52cedefecb8874a984ffb0c937785ace24880f47605b10b767ab8fbf191841d135626a91ed223347ad5d17c129e623ff0c419b55cfc0854b03fd2e6f9b1db0bf1c2d93429a3ef1bcfc82c6e0e739424dfdabe16f997;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b09ed62608b42f24b7f531d5b7fe99bf92797cc4fb896e5d9e6359a4c95007c22904d54fb3807462ce953a3461e15b2e2ba298126b492f49003b1ffa11ee7c88372db9c09ffdce9a07a5d17cc78199537f98b989f685ef83cf628069935af4171dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h218c56654f60f8bcc029e1b539877f25774f4d55524885969f78c3a613d0e06738af7c9c9c4f79536f761f92eab5ed0a1ef17b42117fb3965269ff0338c42245ba030ba6790538b2b5647105b28820724a87af5b2461ac28b812e0179d7271d40363;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc281a64ad26c9a99927f0f50ed3357d20ee0dafd0255b713b30170dd7307e491cb5029d3575c21b185ebb2c9ec9c5fe53e33003bcc555bd3f76e7f8c19d33edc2d819081c11beba10ba4da5f1efb5795db32736e497320481f984b74a67b23a90bce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd23d069fe95c031fed4146e54af66ae3b1a0776f5db49cc824c66df23cc68cd1001438c6042be3b0dd0436b25e457928b0abe2afcada33dec1ef1284c680f46c979c0ac4a7064cb129f54cdefdc0304d6828a25240eb082827c1df99bb2a9e870104;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc94fe7e6075d9d68a706ac0521bad7064768f678daf44721aeddbbba15e4847f0fa98daea29d85f7639e50ef53e37c7052189d74ce0a2a8b9637782f07a5e75cef5b5a6c431e521b66cebce9e46d6615f031bdc9e076212a09bfe153cb5bdf9b5e6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1146c8bafa038b5f43807ab42663f1cc5b0cc07729df61ee98572358568bb5d4d20bbe70f030a3a98c23588991d002369bde0f645d1938f9f784b24f6446bfe363f78337aef796dde3af80672848017dd504c6d01f7884df193f3f3bb447d6b1b6ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee2fd53c0ba1f0f4dc3c6d516bd9c41256bc7ab7314c07ca37c25be26d2538c6b5d108534387e7888540bfa81d65c87178629205861bf7c8e5a3ff56f5bc972140402f004a2beb511d65ad6172038f963bbab02a9be3e85a367fa9dbbd04548329bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20e721d064b1e047e99c2f921a0f68a8bcc004b482d3f816e695c4e776715f07ad973cf06ff50ba5154f182c6e05f80fdfec5d33a8273aa25406311cb44167c28ae39841c8c52ff3d892a227d3c2f47b27e98d7994a338a49a3b8ac39b5c6f5d38c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h690f3d0a813172a56c7afd5d67e1f721714a83cf361b7d72f2ecb403930109a00e4663a4a5ea889d337ef025e3cc2de77d55f60a734d6ab00d949a99a18d3c129e253f3777043f2362d57a5e0be26be80380a95b5f2acd4d6ba4d94d689df68c3dd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75012420edcb7a9344dcf46b2ac5329d971b211bf57f3e77efbd2976b0863fb3ffc54da248618ecf4032992eb43818cc7c9b8caacbc1581ce31bea10b200d1fbf837334a8c1ed258112c9d2502efd15c68e9f5d6364504aeab23897afd3aab061f63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h705ccec2425904d4b5ecaf7fab72afabc16a8673b522016114bf579274b2a9295b94e691df7930a34bc3a4b01c707162a78c3cd139c079069f53e4cc4a5de4e491ff9a0c0baadc9de0910603ff2f5da40ef650dd019f29dcf21cb5dcbd7305d1420f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac833c4c19aeee37363bb86f5587d2edaff760e85f8d441aa0ce324789af08d5cb6ec078f373348631798c25550c0e94499f746e1253fdc1bd6a3f59ef8e0914fcad0218aec47f637c0eca881305e7957a87ca59d27730af57b2e91fc15b9ad67dff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0b63ea64a2ff048bfa1a5553625e07a5d4a2331a2f85548cedf10134f1a376dd48794f71a13576cf112a02fc71e9f0af900ea5af8af543a7eaca93fe86a41381c6d5d082ef44487f230652a36319ed4d0e78ea616d975fce06b0f997e2976c0e9ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2743c28746c7c2374493005897a29572fbdc586cdaf9a676cade114244396fe4767cbfd717d48156efa9e941918a4bdf60c14b485841162928867e443f63fd96573af4509958cbaa324d386f7e0fe291d9ed9b47c733fdc9bb1340fce816a521d489;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33d282008edfc2c32ee847942e783d3df29d6f0cfb27bc184d408e86872c4b0438423d0c0c9e1116803c848e1bb9c01e81282114f74f4242560df2b9796b6e2aa0fe5ca3c6b89993435f4b86e34101847e120270fdd2a36d5edbff3826acfe12c093;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h126a1f5f4907900b5903ab6466beab2ec167fcc9233515fd49ff8e2deab3091a44044a52bcc524363ad8f5a63b0816dad17df93f0405735615a96ba067c92e55301016d9a93fb594b7c852f282684dff9f9319ecde6f6198b65f28eadfbe1946e1ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a3aed090b2cf3f534eb71eecb204de89dd46ad2c4bbf75c0159aec26ec4bc38837ec68d3c71f0038e519b741b09c42bedd3323dc13c29e953e4b0fe916d67b5c0bec20ab936bdd845d4b350502b5a57eeb73c908971dc561f69c717d85af9569f32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd77ba3dae2508fe598d5c68371fd475cf3f3ae30f514643c79a60c28682659bc56cbbdd52998defdf1c49d779322f26dca6a3b6ecbac66558872eaf3c25d861683ca7c0e0679daf0dacc251bbe3313323c068393d99237f3932ad929b0be212fa86e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0230bd8b73994df933f76fbff81daa84dd460b7ab374d46ac475fc4ef8cfd686c880f1565b643d50e242a7b352503220623939a6e127bbeb43c973e70f42a4e5927bcfcc4cb43ac4e0d0905b9a6b17c7b23ca9c0baf2522117ba35426039e56e65a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8da8cdba8060c6872355a79819f62d9dbe3d7a6b369dd4e0793d604e899bf1daf1e7096ee07f3e76e68e96af59e3610f7314f1758f622d28f2f409e8727130ed4e230204c5ead38950af59102a525ef37906e6ec156b976a5ada37532a5e8845e8aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fa45532448a8035aa317a4c61914f00066184e80497ad03ba96fff1a227e9f1d5de765f091a3f773525da2112258b361b250fb5fd167127214641fbfb2516aa72f65de8371960602698851d5f2323253c7bf73dcd3669cac9cc9d5ef36189105fbc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7c110b2098a7668bc36ddb180ccc312e9bb54160da9d0b7bfb8fa4dde9dc9245574deea4696f89fe6fdc9460dbddd9693af1d79391a31da5cad2b6b0ba22168fd71cb9151629748e7d23fa45b1dee97d7f110ea65e7be12b225d940f98a50e468d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cfa0e55b4eebcc1e98ceb0d07d7de5a8b7f17391c6e9b03bba4265efa393aac063014fcb0a7f2748fd6b1a009e94a7527fba02d42b5389eb0f6d0486984458d6582fcbca687bdf09d181e003f1ea0cba96ace939f19e25b002b34e2f55835671e33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2f7cef23da6193efdcadecea47dc05e95d526014f4b031f0e1cc98b1da7443c4b2bfc4344488bf0f6322ec21d5820815be3c674a34caffbb0d8db01e593405db973a0832e7ff29756e1f979d9fcc23e9c1cf913dd918ffd1db738d9b3c432e4a0d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a6b80c6214c827b9d4561648c61f163ff8131e5a431a6fbc4d04f8d9ca6ff58694fda072fd716d11ebd624da70a318291a9faec8b4e7290e627b2976024de166db4237f3bf2b66157add1abef4825b5742085a5a2daa98c7b172c9a6e0e5a0c1f35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93ba6d1cc3e52abd028e9001d9bb0d827ad2cc19f7b997a8006d53c246bf95a7beba23f1b0f0985a92ee0e45f2377e2d58f9a992831d4c218ea2eaadf3bbe47fe544d3c70bdf3356b5ea93eb11719c43c38804009e9f24a30ab091b5e018d89b5c2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6776ca0c332f4b483c3d59b6b3251252936afa7e2a0d3035da3bd0088b9c2d7c5dc8b9af90b333aeff81015c4bfe1ea2cd0a965aae9365f1d94d681f62d323c759353b61495270bc8e951839df40cd40345d9ec95b740a23ded4d7b5fcc73631e6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7441ff2068c903f9eb5748706d52ec24d6fbcfedbf138783bbc08f5dad03410b6be82929c877899809786cc39b8802d085dca394e1c1d4c1fdec70479b5ce8e2f54edc0744e5416f613c390431e1cce6f10b27568e09a8e4e2dffd117ba498bdb8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66ec78353ee56fa029b5c7b8fc41fafc6822242bf4689a8765d45e93a654ae7e2ee6b63768a1bef0ccccf0cc6c49f29e1d9545d25dc2d4fdcd5966c1735d9d4e00679d07606bbbe7598c70fc0616f8b2bfcd5905820dfd60e7f212d0c091cf8c013c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f602e79e44f85e47d94f1c00232460c24bde72965379567c1233c2f1b0e886e1594a20ca25c010324274d5c70b5f5a970845e27c9c21c5902c615fe7b0e31962b012a0accbb847372805256e67dcef422483cd901638a8dd17514f10dfbe75f99c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89e9d2efd34b738c63dfbc8b492eee6ea19377fb696b720b1d58291a39f2ae819e398964cb8bf1e40c89507cdc7f0b9250f906ccbc87f6d2803d671507622cdeb0c729b5131fb147c926d1963d95d19f3e6c3c80a316e66c063e0b561299661ae28b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28915177b475fecae76f28d0a1926eece9f4dd7a1f603e077081038a4734ff6ffc4e0bd79149e69dedc50bced6ed88ff99090f38f98ec655ac9742d9fa82ab0818aec2ee4a8d64f1ccbfe9aec026cf30151dbba7a7e2a1e72935ee964dd8cb258422;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e04cd0c603dc10f4852f89c936ed4f22c1f93a70da3ea9fd3f2899b2ead073bf310c79d3fb2a9c76dc21c9f10ceef05425d7c5d2b54a9597834587d7f45f27b8a598a0464ea814b1f2c575a2212a2e4139fe45b42b773abe75ee5faecfad25297d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ffd1fb7c72377f7d51287f1e10aa22c498f48857c634b59d88f879640b7c240e64dd6312b23893d8519073c114aea6389ba7416a5295e9f6e31e7f244c58b6945ef1a91303a6144e0ba434f082453f1872e3b209953da4da0f7c1f7001e52173b4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34db651e9614e702bc666b1fffa29cee057dc7539c2c1ed48ce1aa460f372f1c3abc207b70a0ffed3c41f643dc7d5fbf2a89029b11269d06c01e5fc8e4874534776779481cbe5e47e63598f07d4cf93ab0cb8d882985828c5ce8254668321a5897fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bccd2a6f844942d77f68c5938d0602e2007054d547e31efa89df2d4f03115af6058ddbcdbc1a992f3ee38b717c6415b7532589abb3ee852364876028ad088c12ea3053001492e4313cecfb69ad19567aeb56536cb32fd79f230d0efb81a3e6d3393;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb598a47080290d3d6c064bbbea7d339eac2a7714d3a13c4bf1c2573f081ea5855aa0d0abed9ac733b9f01f863bffd5f95ea96eb8382e8baef69b4bb4fce0130ab2c97345b63fd13acf9f6dd001085bf9e6740b43f1ca5f462425ee91c4352bf2103f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd719c87773afa826e2a3f932538391ca07e00020593dc1b7c4d18c418e1aafc3ca422ec508dfa0f96a47eea16a28c42e137a7d235105f159a2424e38ad71815a5cae683c4ad8c3fc2e9f5e23e3b5c902d54f0103ab721551ad5b9339771da814952e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1750094804d1d524603d0d838bac57a55653079ee636703f6fd7fe84204d35a4b07c3f2c6265a01b65e36ed79b5f4fb2ae4ea3f2fa2b41e5dc476e3a30be013ab9f22eacfe9475010e573f2d4edb91352f22f53aef7d17e53996956da22b73ac9e60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35db8595658d2b7ffdb6e458346efafcef656cef1494bb921aafcf809a11c2b2668a1cee92c11916d7be121998df281356d3c4d293db19e26554902540d50e18bb181cba36aa1730a6eb7d18ff063eea71f57cc9d57cef6cd59482e3f0b9d031be2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d9d6c94a713975effbcb79fc4cecb9015e0b28f6e51c23b51ac012297694a58422f106bfd10133d75c94d40dfd694b7a40e25a36b4e417e894c893f085f880d75f2e70f17727a7c9fbe9da8fb9ade47afcc7fc471de4bfd55d83cd41b6a2b8fa138;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1506632135538783270af5eaebbab4cf3edb7c0b74619a0589bb709b710d9ec7ec3634ba82967b00edd1f6063919a2df573c62c8f1eb203e86017d7455c9fcc3e8aa482c9429578ea0fbdbac516b8fd4bd6793aa03c89ceccafd948285494e7b0e26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfbf2b5ac79841f55125034eb079b6c0a13286e32433994d19d99d143316dce380cad3d3a0e7e6cae6d7fe94cc94a430f53260a403f00ddc316d03747575e6d3f6f1929fa96f978ae4002f8bf98ff963ad830bf35f0917c53507fb1071a4c7a64160;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d2d3d7b9e30f2ea4a2e9fe3541baa1f1defeba0e64af41f1b0f6414b503560903f7f4edfa1e08964fba5024f24fe4078a5522c46104c5b09ec8030c2c1924f95140e28e59f6c8846bd135c7dfcab04e2ac94265afdf38edc31a46112d3649393302;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46cf8891434469eae2494bc1a470d59a48f4daf13217915e598d36e8e3711de980f7fd0c0caf886222207ff159c3ad509b52e7ff8371d313d34952a8c5e0bfc7cc5aa23e34a1e8a9ee5bf8c03487771b83991e7c7f58272de8efd4f483f8764a9737;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha46f1c5e8f1d99bb61bed32bae26f865b4e6c79cd45560705e4ee05c26c1aa426ec6c995c33ee619fad8ce780adf403e24c0a097e2e153b1f14927352260d904c0e51a76ebbb9e88a71e89611b7e2993f0f1409e674ab57db764092702ef581ac628;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15846bf60b43625fe6ae4ec5bfb6e4533a69242aaf5a49f113451ddaf4fbedc6d17e3700ef923e52dc0d360c2a8a212d15dd83e30d551ca760c0a84bc473b128798589f6140c81a8149744f7416698f804bfbf40bea562f1126fb64c785491d47bd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h901ec6451b0d2c4bc9b3287cc715f875f8e884fe041868c5078c8fbcb0a6ad5b7b749be74becfafb2111edc88c747eb0a2c7ad337d6ca6dea7415c4e2a38eb9fa54284d6ae1f92214864bfc744aef6b3f5f0e8a9568d80922e3ab755604058880458;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfed6b536073f55dae2348f6b1d3bffd8eb353f897ea9d8a91640c086176406c0d921b18fd6d6623bd085be6ce808087ebdc4f1c16e805b6797201d364c42ce2baab1f7b3e79d59b9f27a0a093be253aa1af1fed0707fc7056116e773dafe798747;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b5ea747e0aa90ccf63f1c3076b8274cae110668332dbddf299d455d9428232a56451a24b654daf7f325cb7d9b6cd25c3cdd7793bbf8fc76299679e1395177e9b8e022eb1afa7a0892b3ee26a8c0e3afca22b40c0881ee971f3f831cf5ecb373919d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25fe72b70499355c5d73d22dec871037dfb23ba97f177c0678f6ba6a9b575b8b5f5820338a63a6ad3198672023a3a44b009d11b321b493b738cb6fb1fae64d2493f2162750a71bf7defd28c7def1191dafd3ef5996df8c9dbf0290929d0c0e615c4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d5296649456fe9104bc84a9db6aa60f37784abbd90f5b0482816d15d8138b5d8f8fba62b1a7837c970752f6680398c562a5444ff7323bf56baae6095e22477aa045eaf80558ab4732bbf803126978e7034e3a0303ab2ad10c68b41762bcf0a08b84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebbab6c428c60d8d9d52d9ede0a09bb79ea55eed57d6496b83e6f035b2e3975cf623b4a26f3a4d7b96a516da8be48a332a74151a52146e87ff7fd114e4ea9c71748686a01c74d159f556b10b635963df131e6e416a8e0d9b4003025f4a959c9548a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36a1be2474099c1c9e6258a19970aee6823a9e749dfe2e5893fbfb48901127d5fda9fe3e1a82b53c9b34cea63a5e14dd878443602c8f953484133ea24747388771e32c627fef31b546b8d0bfac834b7c856ec3b6b1afc33f4b0ad82b8cba7d31b1c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b41b9c326f4e2af6c7013f0dad8084bc31c95c98dcde86c25b2010a1be429cbd1cbe0db9e64e7aed801fa401854a5df23abc17ad9b1ec6a7e2b1118b28fa26bd29312d7c1ba994d7a1634621124df0befb92ffbceeb47c77475973540a11aa361f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1bad6e8e8c6af27fd86efffc8f3d120cd00bc4e48d5693e92c5b9a21b045fa6d5b6689e400fce0eefec2a030535b8a05738a7be69754db9c48559f91f2aa22be7de47170a1020c6b212e068644d350707df2648de370b81f9d3cfa9bf9509c71e20;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb279bb87e7c1fbe601ee7e863befd710d7d89f3184bf9a1315d724f67cb26436bd996a8a348b6e970dc6071927c8c7b36b005efc9456386d04b035ef4574740f17210b4b74b3895243103294aef361b7cd5eb9ac91699682b9e495012807446619;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdc6a0f9c970b5b620ff9c57e1aab3b13dec965037ae1a9d87d1589e1c8550be69c5c8644ad2c4bcc882b1ddc7201a481b4f5c68553fcf4d1d51cea0b6e7f98f0263c38d3bb9caedceea79f7213285954ad0818d3819d09e778596b75e717d2a53ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283b4d9499d3f74fa8bea522a40c9a219f00b03ff21983706708e6300bcdae77b7eab7efcfac5c7032d6ba7dfc0177657f3c4053986a8677e889df89cff09788a7f3ad2de133af21ffd2716b2bfc5aada056a6d0863b52dbf25b9e4b1108006e97e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7129b9588e704d47a5f5c39f54dc91978bac5e1b8542ab8bd59f210214ff3fc82dde35826276568841dd37f1e79c163f3c22135106af0538c01726ae5096da9f40b835166be53c2577c2307477a14ac48ede4b7726f234205901ac103df350e5e4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d47bc5b468298c3abc90a02ee418fbc220c809c0ff9da4c2e9ed049d491d32146267eb6bba3b85147fb9e2d44b6b541de276c7bcf74b1c55ad23b82b275c08652b6209236f54528788e11a651df49ab2716e19d6ddf4a7042214ccd26e6685f3a11;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71861159bb481ffd1136d44ab8c43bbb124758eb633b65a083b4a597f86ff7d9223810d2bee7071ea57cc226a394cf114da545f8a8443ad0f18f0f8cd784dbd8f7e675e24f11f73a2325d4d724674bf628cabf3fbe5dd16cc7e58a70358aa6a358d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81dd582e95392f0b262aacfc5a0bc1e9664f8dc06c2b74f6dbe49ede1c90eb8295ccb217dcb5ba5c07c767654a1391aaf990e804e37022a9e4a25b863d6f399f0c1c41e99802ccdec7ab2fa455f3b7995331d9237f2363e90a80f987262f8475aff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf6a8a385877e8452c40aa825815649aaecbaf37672c162d72496292d9fcaed3b60a727c4a4b99bf8b21318bca1397001625b1fa03d33e34f7df42c7646bc72ca6f0f981f882d18f8ca63d5d9b75f5a7cea5bbea5e63b5406a99520099eac8e49f24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17cf6cdc7a31de879db5901d6c5f3a903d860d51523fa885b682b0c493e95c3147a58edc94fc3f89eb9a9a9cd5c325ebd252e468b6d84836882019707c45c96f9d128d3ef2c176520f7c552339ff8ec0db714095d9624edef13d8ddf095af1a5876;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe0b256d07c804ae14cc44d2660922b7b582efd217538b0e745a73ca1f6ad3f10ecfe4ac3ed170aa742f858365c690dbcca33eba45aba6a533dc858c89296dca48919295b8f67c46277ff4042a6e1badca3f940c4bf9265b61573b3527a69d6b387c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeec14da91f12af4939274e58e1bb5b0d7f7bc9a9df49e8998b40229230f4e6f8da4e2ae554adc9cae0c1d4cc203198849ba5479751565e48fcd9d493b242d6d018db68be1d0a2aadd1315bae6882ce1878d3d7fd56831217294b0e02ad9d12e1821;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd41dcf8db5d54aed0b96c3ce0005b4b302259f656e2628ef7632f4570c51e3940d966b4dcc8024c023f5954a1a75fdafa3e35f963d661d43e27bd1a7df1558b838ea9586c8a159480a4c679f555c50efda335d86489dca800def4b5db8ce13169a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbc3f5d4362bc6903b0385df5afafd6cd30d52f3cc7006720624465f502763af1f3f1c06bad3fa6a05b0cd04ca9566c5cfcb8c48ba72fc408880e560342cf2af07b59b0ec3703b7d773ede5f81380131bcf14726fe7cdccea6ff98886e1fdfe07ea8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h819b35f8676f9105404ecb0f9bac0c7195050c66ea7a83a779d3ee8af9a825b4f7f64bd135c2bf99d32bd4a17b041d7ad78983873210c49f777d5a6d9fa2498dcbe371640392f918cd35d7a71741dd05504ab0eb95589e9870ec81782ebf660ec679;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31bfc441796eead0ef424d0820d8d0d5a0af6aa7f1151e35835e110bcbe0d89f3eb756c22d36e5a31e77797f147b8dd2905294440262de8318e789d89bbd1a96acc6d186c1d48ef31d3d4c8d0854414b22523e4b41b594a9558388eca0981159d5de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3054aa7d5d230159af7452e275df233b7ba54b2b57b7ec481520c573861ec722f9f2fb6d3ddcfd9bed9495abc9e086d08975e4a71d11de777cae98e544c8d0b9096fdf39c85f610c1bf6ea57a69d0a210f2a44f9dd03274ec4240c8d71c2c97ef1a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88b622fde6f7e9674e256433980daf62fa9fe16c9b702e86d16401a176ab8ad6ce6f878bf4ac6ffcc9971416d3d2da2aae715c90a78392bf5ed587f3bacedc035224fe75389697dc4586257e0af130afffbebad6d3102bf0362f5d831d88b1a4b964;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d952061e10479204d5b7f3fdf4feadc35fdcf8363744128af6c54c45c5334109badd1213b14dfe6bfefea8ae2a2d135ede36c41c0a0417b40499f43ff4ec134f1180fde801e990a384a5912b25ac019b9cf343492acb314a1d672b7327426950024;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8034d9921b10acb2ba792735961f7618fb1c7562e92c274fc9c33439e55c87889bc685ca0687c267c5caa7042217e959f5cecfcedf1ab99ddfaa7bb3e30b1db85b673c3bf257cb914bad085c4854496e7dd3f95b87db413bec1526127f2f01115084;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h625f7b9238810c690ab213ff45ebf3c34c3d58011117b13eaac11f03c4ac3b59189d468446825a0a08b457e2786b66f99b786969f2884ade2dad0b648de7b0e4ce59ae2cfcb8a0ad2857c326eb5767faa08be258ee70c89801d8c93dc0d41ca5617a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35077077e4cbae912658385f82c3034df004f61f5ca394e1100ce0f916babab43aad888814d274384785ee843f6c531171747bc5702eaa929b200d100638daa25bbf725bfe3099e140d5c62008ffb3ad1f3759eccdf1afcfcbff15831eb002fce8e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2125c1e157fe337944e29c4bc6e0aaa38e8202bf306c3223c4237bc2ca84f8da75280dac40e54e00a282084275f67e788bee5d57e5f9b1434c5ba0dd997e0f5b1cc7398c149198081a44788d634cdfbe88d871447a098613203f455c8101625a872e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28a943e1f90f1fa1116768ca8ff0749c04e08c99725b4dd533e1f8df17a0b69f1cefd62853ba526a9bb0da5775b4cff4238cebf415ed67511970656e7a2ec3991bfecc682d80eebd00e58d1ba9c1936b0924cfc02edca4d78ee9fc85bbcf7bf25659;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32a5bb570e6047e80891a3ba5f13def1a49ff9dd80fbff2032bbbdc81714015cda08bb5d40cde1689352bd7b6983de4bd31d450cb23e0842af13b4edd42096d4ec86b36ff7743be4c509b8676d7d2edbf25a8ed6f220c0c8b398b3a29e3960f65501;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcba1b1f4297ec324b39bab65544e2e4cc39ffad97de68cb78350f38a8eb1f517ee51a20df62f36e73e95da760c1492a19c234f4f625a14062e68306b699c79c20808b483c7722219680468a4e3bbf38729399c0e3df08e12c3fe5336d2bc23235ef1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf438a588e01e49711e0603b9ff7974d10b468d7090afe40e25e8cec072fb643e4e230a8a7f0bbb091af4cb3be6dabf84a2342d71ac097e765d7a32cb9a4933abb449d0bf7ea16ebb35f46203a3edc42aee09eec75ef6285375781bf33b96228d47f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he33fcb26e7afc077bd0666e6f17bc6f806511bb0877f5ea1c82d4afcec51023c590cf318f0b63705bdf8b5f9eae404c222924d52fc330306ee83371e7c24a42ff422a9bdaccd98da6639489e38912c0c33df329c78327d481bbeb4e3c9a2848df6b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81e2b32eed35a8020642176b8c88adb56691e0b3250b962e76d4b1026a625c94df17127952ddc68de6ae81739d0d0502cdb40300b53fcb64d24f88b6f2fbecba2dfad83c4e0ee3850cde7d579fd0579616d6decccf3c565aa8ff99269f691a229f65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haaf69a68665bcb52ea5cb728480d2a2509c259e81018e46aebdea9bb8b564d44e8d698bc81a5295c71c3f882f25db2421382c525ee5a122633ca90e43bada8cce8ad2ba1a0eb25bba3f170e25e6f2f4e44c76e9d2ff5b8d981d6d8126d07e85e129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7beda9433c91215da9163613d54a4d2114df63df327205df69fe0baf9af5b34b24dcd1145d5f251bf4edf7dd0004743c79e614f4b815f9d584353a98df11edebfbbd341c64e1f384103d5d2e014b344f616f30f84b5b6d4af41c1bec0af8b516ee90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44924685a54d93f1ec5b2759750e733938b573361e36641de398a0e06522e71aa825d0089afca1963a1fbf15c911f7e8b7bf9277df4de3645847e940f59e1e8b3c71b3b207da6f0adb3cbf1acb73fe00a6acbbbad6246e1977e95997ba6bbfcf2210;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8035e39a9760c68d71b6ec9fbc7a657095c706406ac2858f713307f05998e6f66565ad777c2a30b0b7073bf46db7819041dc1200482e7e85c3db5e8c700b106ee4b78f4d3ce8150e4e61f44726fb1afeea79832f23aa63813b82fd54c2ec807bfa68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h512c04bea71e7d763ee02869157adeda009061305dcb8eebf8bdf1834263db81b7980404f37bb2b28e55578d6177c7d151df1eeb0632da1abd2a1fc8ef64640df0aaaa03724cb6da1b2e1a27f8f0ea8af2aa0418253425075c5ed8fe7f5dd794963e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he26b312c931ddc7a2941e87bc5fe58086062469d72abbd83b127a598030f24859a97acd0d3705e05a7217a7ef82d987c511c0b408c80e719f60a8ed66897b1dc477749ed24423613069073b0a2aa6f5087f8c7228a28c4c1e6f682019f0ee49ec473;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88fd57fbfd6bf55fb05f1f5c65ff669e73bbbdfa34804ea54993d5f18a149059affbc552a801e173d3e30e8c2cec478d670913b2a5f63a4dcd11810194833697b6348562d1d250cd7295a48e7d12c1f98502f8e82a261c20779d5bfe80751f1c958d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17958b33f5bed208017fa4515e4916dfb106b86e9ccb301b27d19949c728664c7da48fb8bb9fdfd89be284c7e2d8737f80797d0904b2a7a9212049d7297568f2d798a3d302ce13296042ee0426d4c5de22b7add51e8a46501bafaf9c653cd88046e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10b2be65db4d072a1e672391a324fca44f31fc55486edba02f6195d68b3c4849b522af9d1c38882760e8a77fed177eb37027a3eb2ee4e26d3730fc4647af1e9b6e0aaa2082c7c955afbca5672f17429264a7b64690556e122851ee15f17b19b5b642;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67ad54e3584d5649e2770fa10e3cadda514d85e339c54089300b8b6efbaee47ce19f9e2256afb687c02c0e13b181d48cab0b26578264aa6ee5fc902f8570719ec9f7d1a08715bf193adeea7cbaba3e6c963515cb61eb88e5d15d0c7b5544e6aebf78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10c8775cac920a85f54add43c6a68cbf18d25176f31da20d0c57eb39c7dc07c74b20d5676ed7b92101338ffd7bc4655030ff2e89310b7881fb0f3f5d193308bf9de97007ecbfb020fd81a98edb46e0f65fc4bfea3e514f7eec794a757643440d9c43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c7ab9a0837561c89a026bd14c82dd171c572eaffc34cb33cc41a20dff78cc3ba10f199eaf32afb2308a1a2e0a98c30aba4ef2102f185d5677888838cd77cdecc597be788216ee5982c607e97b1e66127e36e6a88e1de384466512d45cc1e34136f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36b389f67d03ff95062d9aba3922d54308e916ae54425d8d859a0941a60b6be33104d13a25033c68a6add45a6a6ec845286e002cde81ee8da342bb75535a506dad405c00d883fb7c09671087875f33926af33272dbb8bbe8fb28ed7e43a57c6f4e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b04b12eb459d201269ea03f6c4736fa633308f83ddf72cb2cfc500127d6befb1694ebdd6d812148de917bc6b79ec9441cef17fefa0cb2023c7d91fd570aa2b307addd185139232ffa1ccd57b00921be3a7d94a5d70cdc8cae6269a2aa9defccf559;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41b4d035fb4ba003b181b7b91cb06930e64affd9569e4aa8d60d76564b2ee3c1eb87e1fd00bacaf508262e06005fcef57f16ec7cf008d22a386ccaddbefc4a1cdd6aa0fd586363edde94d457b580be1135ada3885ae610badcd5f7efc4901579b566;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19de04accc00c44e99a859350153cf48bf7327dbf02a42744ce5ab1f062ae2a28ad4a2d074ee0805c021e539e6ecbb7539d7a890b209ddbaf8e7d3bd30b4b3bc1bbe2cdce50b4c304c1bf48721725f222e2ac7b1ed1c02ad2de0f86d4d45ec9b2a5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92562de3a3a45548fe388119e8c9ff1f54f393385364b35ad170be6896f78e161e1bd36e93883b6f7f2d6f12e81d32e13687f6be23c6c3b4bb1b341d27c76b6536e310addddd8a6dfa938bb41db3fb86576043d8c1db6a1ddb491a4067fe69f69147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdaa5da508c3f65b1d906bf84ba119a429e09bb37caab51c8aa02bf3c1bba7949919b58cd209d49a0a06a43808aaefed76274cf810a964a1ba552b1ddaaccbab1f0ad61631f86843d7ac00f0f6c800c5da51ab7175e4c36ac724c59a013627c0aa7c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1249305764ee85389edf37b7abe700d52b348f7e27dd19ddf630bca2e76b5bcfd28b78d0389ed17d09e63d27a97cdaaf1f54682ec999ef6aaf76fa731de8fa626e11b5eec0ffcce55c905f6ad28252abd992b7c34f71b6f2da925b891b6ce90f3832;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b98a92e01be251f78e4d5b93db80b79d8229236e43df6e56a826a45e3fd0696b7513beb56ec5f5a9c6a4d1967c891dc53e133a86ed62c8d6ace0ee9f98be65ee7c1664fcf61827055bf1ec8838773aaab720139a00147dd527cb53484131618f7ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e51b467a8e03962c76e8e48af2e281827c0a382ac7ab69ef4102b57610b436cf607947ee4bffd5e616a81b9d277b88e334e8a5fad7c5ded5c11ffe0cb741568423583dac0ba1115eebd49eeaadc14c36aee9863faad4c0e84c66c302fa8d2eeb4bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd61aff2dd3da6eb4eaa6ae1dd3c3b0036289af970a224ae6df659314b06564d9d004821f6f43df27d20d5b272760f29d59eb0930351f88983a353b98eff24336849ed4313a8a0f594552a0e04a2e544eb5aa5d416870e491148565b8d02c5186bab3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5214d6f0a8d3fd22af1fd5b69767fd48c98688be2b66124e93c2f30d0844c0acd0703f9722dfa478abfcec04b9d5b0f5c7b34bdd90ca3d5cf7af3ddbfba92551c040a6fd41092e8ff39ecea4eedb3bdaa98eb5b87940c6cead78ce04d019ae4fcfe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h869d00a578ef5e3d02246c340e2210f5f4c6d5265aabff3d158c57498c6619d0dfc78df1e1be5d6a9d82e0354cca93379b6e0b7b67ba4f0c0c6df32283c6b547a7ce44dd9d870631bae755ae315f806f4256968579768f4a37443da32fed26cde8f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3292b8b1aad390ad7d3dc256da403262c51347d3d66b59f55d205c9ba096de63e887500f4afe627cdc5786c69cddc654e48e82fa8b0ead4a670e1ac698d7077691281b7b10a9e98147ec8265a2a74e2ca2e03da76331faf876600b728f4d0f3c9e65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cce4104f5a2c0a277fda25fb3f0acc755b7b933c2a05b1e4e8861aace31d9ae89c302b096c2adda43027298e4bdf459843e148283d7dda5f3609e87bdff33e0e3377bfcfe14415d03560be9e2f07721f18adebde8e8d67b6f4891150a3ff0e024e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cd44ddc613954db525d98a1cf7ad3f7c0f37229609dcbf191ff8c7f8de021f6f1e2f9642597c889f49c946f5e29904bae8272c6b314fe94bde651b682c23fce34cece5705d2cb2e3b30c960928178d5753a24c564f4ac4863abcbae55f3d7b49e0c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25438a9946b5da56b5ad8dedc5c4e6116853f3a03dd61e19359f4a4ee9001fd1a69eee58788165603d62ae8bcef8870d127861763791941cfe2e46b5a930d35966d97a045f465543abd53285d000d89a8b38523ce58b8b1433508959edddf7af5aa2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19d1322e6e53bf9d2867992be76e21e715975610aa9acac0b04c8c93fc3fba805b3b329d8813788353d08c42cf827c64ea3a187f907df4ff02d70ce676b667a28d464e8c552875d74c733750de4e1a2ac03f8ed4c747bbf0c210e2b2542f224d96ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf5138b9ad7161d13256e850ae9d3e03145ef982b8c3816af607dcc15dbaf243e29c8aee994d91421bcb69f9bb310f3755dd4d5c1fb6b6130b0659dc5df8e82bd709275f105fc319607e36e68221108c74432895a85a3154f5aa06e93734b959fea7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd8237fccd6eab1487f23fd0037ce6214a022fd85f6d8cac505216072bf7f867df52f775bbcec8ba19f6bfa6c7afe318bee55bded9968147045b6c1342b636df892fd52532d1b2eda509be790b2e72ddd2d6ee920b62f9df7a6164df78a7a8e412a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4bd0efe324bafae96c08fb1d50d4bcc45c8d845f9207edf33fa51ba520f648175e9c8983394baa33717527de663afa1d189ff5ac7e2a86e2bb5af034c41946d4c577af49263cbe2eabaf75bdc89764157f947c176c0ec2e402233aca32d7675052c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8b09c6624bb2a6a97f807cf82848a4a7651fa784f26a19ead14a1a3e895547c3984f92ba48b43b6134bc85d252f5cd89f8ec35d84f28d4261bd4d7a5f7a46ca34bf7cb0b2db85cc3d88fdf340d15aac0e8427d53019354c8e8f451a7c1a32824bff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he41a76b4b0e9b6ba722a83dd0ac814796b079e5396f8ba0dc3866cf707ce26c499b2b58342e7f89bf0217abefceb362f4243c46e69600f4efff40553a074ba7c0fac551fb84c01ea16681f4f0c9fdb913454b29c59cd9eae8e1f6ce1845a275494b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78768987ea24bfa6c33a5cf5185f31d69ebbb8ea82285f6fca7326b6ac689369dba23312989c16fd80841b8671f44b19f2d6102dc339090437f61d6d8cbc97d8f334fc0783711d160cce2d0337d19e5865fadbe85243560fe7ef2a4288306bc5902f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52eda6d4c2ad4917912e445216c5b6f93edc15114ec2d413035cc2f824465c6bc55d004ac8a9ba17a5c918ceda9a8d4b524bf0139c4d9c8ab6b26b47c12c14549a96bd8b8d7548611e7bc678110ea35ff5ad07d66cff38b13d380b7172bc725206;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha91af31130ae9d4b7c9518623a97a37307ccc02b9ae7827d8168b9fa0e8841577bb38a9ab47109996db7dedebe2d17fa5dfc3630070fb5b24e078ea4b059d11f4402f6aafda8c6fdf380ac7b61653dc403b089bba21625ea1471f5566a1f9474d8c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cae74f6fb23b9acbe30a4716743ecd113824fcc1891f40345b66986b50189b9855090ca5e3188926805772c894ab54ce7cfb95002c90f22d5b503db0c339cd2fba26f16b9d324c8072f823386f1ba91d7f69e90aea2774be801ce2fad7865f755cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aa02b3d1300d15d5b0353abbb3abaac8f3d40a06a8de79bf032ce9ea2e03ae4a292a3ed6783863d939757afe8985dc7321a1382b625efb889de39cd485289f20ac29451509b7d4dcaf718f9449232717957697fd55e118d9b987efcc66be0a73e5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf38ac0e56a955a994fa375aea529169119d18a3aea45c8ae9619dac34c2458ba934b90f4dc022a72a0bd5e53745eecf975463ae92cb9305f444baca987f16302dcfcd7b5994e02d5acee95783ee64df9e78bb981bdcb6c05c08b520f2e289cca52a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3276b5aaead37690bf47cd986b2b325b2912d5cd65944a57c647cbe5485ac4bd29cee072b05baca1f340c10d4a6185ec8122ee2ab67e9e0a35b2d291d6ba60e8b8a40da46f2e0ff73cd751df11a70abd25ac9f7eaac3ee66c2ad87519ef5f16ce11d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he06b80e70e6e1830ae3af45626b97b88844e18b7d5d627b86e04749d7034c554ce312b8ddc8bcf29ebad1af6ebf725590bd1bb130dde5a74d8408d7829e560019df37d949547e63fd302af8a991f245d690ca456c0075ba7e10eaa7ee06050f0d0c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2a2be81f93c51e0f39366f6a8e797fb8d36dc60560e5d527fee3050a1ace5f9b03c1369612856ed12065cd58a3029a6dba4bf747bcef2466670a08a4bda711352f3e5d3faf913a89b3285e361565fb0135eb6fad0b4e84ad7faa46966e36860be5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfb1daf56259e7f6b07b6a1c4f9ccf0fac27a5cfb9920f3af4220ff3237dc5f982134351fefb4f6fd162f7e403bc97e64fdf22edaf3d2054e9447a589027bdf2db8eb441e11931034768decf11fb4ed818feb31bfaafac24d22e62b3c0721fec6cbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2bfb5d9d933b1896989a60f4bb01ed46932919c377caef3636a50da3ae9093ea35e2e6062275214cc94a6d80d4223976382296e144b4a3f730cd5896426834fc3b12515802ae665b30d6f184cb2f8cbd95c48657a7c0ff26a99648745ba77f10dcd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb15e1383ee698666e0c35835e98cc450182323365a813c26cba08a447f6caa1c52c3169191185c3f4bc6980fbd290c45873928d9c3381830e0b220673cd6cb07528b4a94180a2423c80ac49c157e9cbdd4acb6a3b25d766d625ffd85cee61529de0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb07cd49071d954d96ac6b2e65ed647feb7fb7fb52e0ef9e162014ca0495eec599a86d997bfc2417311da5e9a94cc5879b59ed317313573728363f82dc94775baafce1d1963526442d73729ce3919bfe8cb403ed46f20afb965044a4a6e27309ab2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha06676a63c6257a612e434284526e9cb384c05734e9598926b9c51de356fc2b22de31e4c16f483302adf25c128b0b17de1a9009a5dc7ffaf64d393fd9fcd5d835d53bb23c2b0eaa9438a2fb259d64fd4e1cd17670740fa65472dcd22abd7a8379f93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h451a90e83c048249ce258dfce506c961cd6e80e2d1d61b04df376ff320ca70be97a3840a06544e1ddb5cfd4b7f6e333dc3111f50dd137eff08d5da7710ebdd8aeaedc9e5f93eab6796568e5f5c830e0cfaaa953f36958f53de9aa3874954274bbd00;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a062b5e0329dc461fc7e759dc21fd775db34d0d251fd04ff4c48fa0fa6e8647d9d5ace844e7b7cfa019b86c02bf0bc15a023458fe21877357edac7671b2ac1fc69f3df0156dfe397118c374134c9c5ec9fa19979a5d3f0b42c992a93080c1455f66;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1f7183c85e854e64f0831cdfe507a910a473c52b61ec9ae2b7eef319765686622e090156a013e0d62f54d9383e886b42caeec59d652f94a8a70c05f5101e51808b0c6d29e32e7faf83185388c5fe1a8d8a9b27d6580bfa3de417638dd62435fcf3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3e2d82260595792c5dbf3b8601013493b911239b7c96360f6b3ecc7d33df00742ca2d4427e3332e9b6e19cf942188d2070d32f590aefb293c8aa70baf6bfc1d2b97ba2debd4433a4daf8b86ac6dbab2eff6a207d90b850d85812d942aadf33c00b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6777181a4df992cab75363a6fd9818e9df6b3f34f0dc56bb162e668b5b152d8c187849a277bfb8cda259c19932395b1f585a8f6554aca5fd2667ccce58b88a16e6a92956f5416cb2b20f6ded83c3dcd3c3c22aaef2142ccc1ab5d899c30139fcd4ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dd0eca22c94b4b890023ea092879bf801ccc96d0822b23fe73d6318dcd87bbcd92d757ad1360a399b60b5344ba48a9a49bfbffd01465248a602ca3f681d4958c84e32fd137949840f406d9c2eeb1263aff7e0b4ff367bf3dda523b39ca0a59690dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55d41365bfafaa4e478b051a395776cc485a3f3a6d4b4d108403ca154d30721b6bace69bf090202daf433425066e8ad61145ae93f53e299cfdf419b3da8e95a1ced304e302b2ea9bf853fe9954d47541fb55a98ea9be4e372660c487fdac45404bfb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b429e7814bb2b77782703da35c0b6d9e9f1333f6c3c08eab4c1a189b65f4e06edd64809e3c6714d5c419c4ae2215f6ba690e39c7f43b0d97a0e13218920058f7aafae1292b86b582a1b47c60b34303c782a5007230f183adaf88bf409d80e8ae14a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3096b79cf7337a402cd246cb76f18c002e15cb0a72ac42185bb85db0d95dd87ce56cb63d4c2875baab274dda64d7376fd3f3b2b7b767507d42bbbed48465ab89d55abff11b89f86abfe9d290a344d3884e4d02b4a012493b4f0ae890d09ef48a881e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56a84a0393d280f0bc581fe6e3ef738ce11f9f83bc339a7c04a93358c943f41d7cf9cf30de061689df1eb4b59421923130432a081b82b05cd19d73a0ed3509239e5b64931929db32bde89741a8a05b063cab232e8132f8cf1f36da76561f62129568;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7335d34c0da49b99a9ed3d3ea644df800c589ac579ab22a8799a568adcb390b26a7d44f2329c5b57dd3aaea90e8dddfcbdbad94997eb8c70c597ccda9eb33e8a166b17b67b791e5eea01c421e51e6b77e15964c3db1178f8f2230f09d78af66b6336;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2de47e3e6cf3d7b5313ed914414f580faa4ff850f535aac965f042946f4afa053178dcaa73a2332614d0c43caebc9733393d7d62c46c623e25b80548cf1b739eb5b1e4a5aacb2532a18ae2cb8b7d8e6d9389969ba46b7d1b7a5f9fcd2d530305ceb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4e8574ae94219bc2cd617b7a280a4a02d05a81fc2c94f320c40a722956d56269d9d9951ea7ed85c79515a40ec1a98554746c7120630db2ddf8dcc5a26c3b2c753926d4d22f4d2469b14405e8a61ca3224808ad3e99e368eeb9565e429068722723b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28efeb650e7355e53d2a4673082a2a0da791bf5b4e0622b258e3a5cc9ecce2a471fe57f7fb1f8c5c8bc37ff5ce02108964b1bab8de1c6d797a235a343265c2205b3ed5a0cd2338190252d8646c9add87be0d8023c10e037f815e698e68a846bd4d6c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fcee84f7df1f266c2ca076b6bdebb53f0b96aaae0f43538c77d4159d78e63a725ecb794e5a58f331d1b5aa0b7febeae950c0c427cc479866d631248586e8e492497c6bdf7b1c8a9f5dd0ca292be5430328152932b77442b48bb294634a361bc9c06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc725c09d7c9357b68592e47a0fa43b71b5eefe4411df5de34689a91f22f8faa7fda309e275e69f74bcc02e2abe39626e1ab78575518810ada4b03cbfe15cd0a1a829d21651ddb104d6e17d18e45b783be45c27f6aab14a6b89497766f715f61eabd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52759e76b661e8adf18df49b569b2f24aa8a30e2489bfe283088b93fe874694d1b2d93dff105c71ced12b9369a601b1d219f45e8be24b0b4dd1f10cf37983e61b8056d36b6ff95834726a1d4d50bfb90d22fe881b66ebc629f34e0ed8c9bb71201e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h760e53f50bfd7b8c0c2c72521d94a872f5c8b72f41db3c6c3aca4f502a76fa6bbc3fbbe4444c565573881d2133ec4c282caf2cdccd9e0e63d4125736b9af96ae1c4d20c670ead9c8fd618977e1b6a70c1a2a8f954f0361a0e23c15c16784c6b593fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf99046563a1df4f32cd347248a49248ffe799c24164cbebf74ffaede9597b2e6504aff07ded1658dcc1453641925e21207b9b5452a66068107e89fadd2375b671649dc3c803dd804a7a72cfed13ab25f0aee8933f4e7f868be934e5e31389293875;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h914434a93109f4c318d5c028e24dac5ab9865eef87532b8bc9e5d8c8ace5f3851d6cdf0c81b3f880989b8cb7adab523ec08586962e79fbeb0480c17853099f2956d6bf9dfcadbf15cfa5cfb9f9c287a7c6b899eefa3f47e0340506ddf0a401176939;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h646ccc3b06f6379a9c5033c0a4f86312962226f2915c9c88404c73a4efb61f9301e211dc57afbaf41a53fc41bff1988450fdfd057b080b515b582803773918f7d25d8ea06256d5f46d6ad22a825087d043d94dccc73ce2ee1de57835fa6abcdfd82b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54e2a2dbc996af8534405f879d6d32674357c2ee7531f2aad24cedff5f863415a1264e53509c8d4ad31e36d82ec9fee33d7a7e814d052a8b50cbe8cd63b6ef4e8e713f2820a8775cf6bc11aaff6e8e39a650c40e13d39c34657f1a04b962d38219cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ebe39c0308692477b0dbe576c02b1054bc73ac84c22b91391fdaa7a28221f9269f79a039f235a133ce441fb521af239ff489070562db80ee5b50009dcd604aceb5c4f9c19ec1850d39a9f076cef088a7a4ec810e59091b385ba53d8bbdcff51aec3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2ca7db504f81784414479d33858bfc14dc5ebca605d3eafee4d72870236b211a26dc4afc93c41a4ae51618e2c016fc2382d2c2656c17b1768b4eff9693424abae2e4d493f1bda547f72017095cc4ff4bb1bfd57c45f345adc70a731f79b3ebd8dfb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ce971895bd04005b9e0d972aa7eb468bf94dcfb3493c6d2a184c681f1ec7f769709bc5082884f96acc76c05d843275bdc16b5b7107d03ce226b14a51a434e9ef65ccac9c7376f1d74826aed77360cf8f91839803c1f7e2b96a680e0be482ff10fb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe3e84420940d3396e25470ae1877b20d4d1d02302a698650f4af502400b2e1ced4981c7a143f92cace693d64c7c84a05ebdff31836e04945fdb601b939dcde92b0a1ebab3bd00fd2008f0aaa75b3a2fe93e299088cf44aec8c3fdb5df7ad47a373e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ce6d45e69170f7edaaa04e0ab3b6b86cc70fa57a146d7738f4a3a481457336500e0046e8b593644f46b14e2730d3c0e453b5234a9bb11330d675162bacf4ea705bb5e10367c23fc935f562fd22a73f48683533ee4fd87a965c99077c81c60bb4c13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab53e64e6acea5f8fa5e116cf638e5ff28af9fc1211e3b5fd8143421237de4aec13fb91727d03f2c8bf15dfe589bd1e0c8b2d2c053a0261335ff3b4254e2aff4de269ca60d01c66c1e25c428b725c9055b6217811eb4cbdf6e3c989fde354997078;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa0d4f98d1e1612f0601258036fe320824f3e0cc19beada42da428584ca09fef8030fd3c1d81438e43d193cffee1903907f69350fc700e6ef6624ede6e6dcebaf9705bc30c4ea609928a261907cc1c02df30cdd57bde9a67278a30b4274dcbce37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39e95fb01891373c6760fc5cbbb1232acb0f7139cba0925ca9020068a3bf0e4534ed67598e87074585dcb1b9871758626d01277727afae4d8dcfce7793b6346d995243c60564a6c6852cbf577560fdc351756c3a139fda9177f46757e0b68318417f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73b37198ff24f048a0e84d34aebc3bc8f9947b8389061d45ebd0bce274bc9a8c7d6467da937aac463af601b0b9b4a8b60a1f0decf865f377e39a2141e5a4521ee6777222271936ed0203d7de252df56bb13b2312181a6902e80b778414cdf094cbf5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a959f9f6d15b076a1a5a9e23d32f0b66a7ef134f9b5f9862c2178880cabed9a0fdcd0e4b988d52dd98445d7d9d9ef4cd57dc76eb056d309078e325b6c6e8101efb4f24267099cad08b77d34139c4bf37667249fe708114844e96c2291659278f17e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75ad2ea7759a697f2bb0fbabbb2d5d4050eee6157527ec468614c2eb486163362f3cda6b3a497996633fdb9015823996df9d840b404bfa81d4584b0615341acb18de0b2c5e33063d0540a0c7d13f29cdb4c9b1ac3174906f76d47627070872821199;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf95a13c3655c6d8c00db71756f10dee20cd0c6deac0d50ac9f6cbefe16de9c2ff6e7b249f5b227fdfd21d2adc98595212a4e14f10818ef7b3ce26c48e45206cc0e48908811d1b80e002f840f6b674022255d546a7857a31ced9463e96c4eb813718d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heafed94a914d1e2ae24c0bec53fc91d17cadd707372313dd61f1fa79fd759ef215c77004b465a9186af404da3ac944150d88b767846b2e218d2d00325db9759a8d0be12b9e0290c01fbebcbea47952cd0b25d084c00dce5942ec646507fdfacc93dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4a2adabcf72783fe45a0b85b4c6bbda087c43498b0bab38fb8b6e8047cc297016956ef1be2a618480000138e5dc167cf093b0efceb119e86b66fb521f19571cacc20e6ad9075cec1447dce416b58ef6f93daa89ca55f4d9259084396fab5f7dfc45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd02a91fe6ae23acfa2c84be998dfd5bef2fce1152c9e8961e5c584cc8f28ac4766ccd28bd2b815232f0775543f80a21c7195164eead67ccd7c244b9b7793227d55163942876f0d971d86293b69bd3e5380ecd320132c6baa5580cdad5074d1f3df7b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68efc26424c9733e5f6c1251348bc25b9779ca215580c9b39681d475e5d69dbbcd705abb2818408e4bbadea859ac2942e591f3f6ce4d197c315615d8ea0942267012419b2c30af0540c276cb5b7a2f696d23a5329314df1ea1d218d33ca788134af5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec341ab087d02890f5bc70745f864366065760236c9bffeb23f0b8608f030e983bd3a85ae03dee4139c98f180284cbbf494dfa54497b7d2f07485373104e14de55cb399c8577c095bc64d0043938c88efbcede43f0bf7d874c6976284e8a178fc698;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e81b36340bfdfa3fd43d4ad1af4da88d1190c903d1ade10d7ad40a4eb14a9ef2c6bd217c8b1510d4087388626561e17e0217f6514439fe570b4e164ef1106700252f7ef6fafe5c61e1c834d44cbcb6cefcd9f242c879d1fc26dddcb9dcb33367f8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b4fb937c6ed334e5e155fd47fc80502a7231a02d8daa53904ce188b3fe0cbc7995117dbf216bbd684f4959f6357f580d9617080d8559847f87910873fabc3599b41077823e6e9bf090baad9d482058f976a6a30b45b952585bb911f82c162039759;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7d8763fb44085f358b32bb01886f612a8cb418477b4893daf7af8d36479976c8f8baeb4be9b45d8664533b959950e501993e582abe07b3da14d8785606343fe380a2da7cd9a4a0d6f4c682c27afec6e175e1b9f45e683170d1d2198c5e1df9091d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa0f971eb12ab4a7aa0dc0bef10354aa35f94cbca0665a02a720098082af74e404ddbfc4443e1fd8ff069da9d7f74302649e7d931f8909c3d3b5a763fb38583e60f50328502ebe963726b5e1686ac9bf43cd88f91c58143968bba3944bae42c176;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc151a04b0c99f332696578c1a2ae420f99f2b34acaecd7f3e39814ffeb1429d5b964a5c57d5d23ba668826803498dee5c63b131465e9e66e039f4598b0a69784471208d760047ba244c1eb9d2443a1db577dbdbda924d8f38c21ccec4ad61224913a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80a610bcd3b663e7d6de3a7ead78add21882c10695804350e0a2248f75d7475e07d1a4feca2e2cb1e71e5d2c2a9d69ade05b50b6f2d56b7790be7d3a471ec0d2897ce5015f0475b2b6e8037654294b2301a5d078ac45cbd6c1c8654a7fb9a8f66d26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dae7b524b0b940a38c6f38c065e36e00d2224ceefbb5e3e5a721dfcaa5220c65899623a6cff29c7fbff617fc719c85077f82959fcb8c06308d44bdb8ae741c0fd9050c9872d6a88bb50ac3a227ca4c3457d2596fefde5e6d5f8414f72f0b194804;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ce99ff365fecb227021b625597608ead1611625aa937d69e346561d7f00ad35309e13594ed96dd13ae40750021ff5f9a89fa3e0a56a61c0c6c937bcc93a0a55ec8344226d222d74936e5c22b57836f0ab2679e0d51d052c73a4acd0dc9df1ad01f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea136330133e3d54a08235eb2025cf948c90008253c4d3a6d886b9cd89dbd4e29068a87d3acb7650c9d063b6cb1adf00b1014f0051cab6b768fe2ea03cc18b0c032e7989dff08e3c6809a028f0a3733373906c29f183a833c5ca8fa9095275349b61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffd42dcafb9c9e65575f6b8429ba8e544dda7977397e56eb8daacb57b5f6e69f2ccb513467946c086b1dea6ec13c9c4f9f49e6b6b565e9fa724a9371696165d90494493a9b14a6ed980308261e8807d92818ac20f6f18cc4b19b79ea3cc270e208fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c99e48caabcc8e7debe82a7aadd66b171ac6b7bcda148cb8b9881f0500a7de5f2fa02d9e2ab66a0852273db0eac2760fbe76e62eab2dd5e384b4a8de5e3a7464efef705dc200b0e3938fe440edaa7c2dd0ad6eef68c9c8de6c64e93f0aa08ebcf98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha44fb5991070009b749c2d66c952a07ef0cc267581fe24578afbd0ccf8644f1cd788d07341ebf298363fae2490f7e1a1ef917606359d70ffb806e73cd8d9a60290491657671dbfb4bce7b6f6b561544f2198ce6e6028461e31ecd0edf4ef13ba8407;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8388f2536e6210dc78990cf2bfe350c9d78c164f03afab1cc4e8eae5bde5b2a2c8f84b84f217ab5a5093d1d811199fe8bd7d3cc4ff786cb1ab96795177ad8bd56a5d480d10a29f8f29a917ca202e82766fba5f9de1a53a112a8dd9a0393a30aa1f4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha93b04f36a86d7932e404d06ebc535674d4138255f427139ffd9f8b92eec19f37998fa38bcb452ab7133be5f52ba34c94d85167a3ab4bae3a661deb43ab59f292e4390a3d49c83f0c72aa12a89bcd15279746b3cb18a1463523ad020647e1672aecd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6db72ae846299892796ab66d1aad6adb558532d5fff1879adca7e5cc2aa81a6a6b653d903302da9dba91bd309cc5634fdb0ca22d02d7dae858097c02699a3746e51bb9fcf234b32ab29ce07262ddf9265fca1b9f8cccc0219ce69c16dbbc66103da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfe10cf232fd41d651c00a11d3e5b5636dd072dfcf57751134201337c9cef140a4fd25ee8e27455887e183ba380912228131cd0a19ce3395a80317e2447ef7bfd62c0b1b48e81a7a3d137b5bd2abcc99f064627a8ae91bdf921dff326f9adfff25fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60a5f8d1c35a7bc6c399f13688b21a706c20f5d48a23d23443ee1bba25d3c73e9c2ce676eb3154affa3f2c9bece83aa8d84e03367fabb8c3eae2697e38cd7a6896acf11af7f21f244f0d1ae9a1be21f721bdd14ff306b5018d53d1aaed3b6982008e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7be88c96d09c287000f26a2c903d7a47a7662380ef76c5beae25bec59bc28280927c44f363b316aca0129d586f86bffd18957aabdbc70925918ebd697515b50ed49ce3734e7e961dba7d1aa907d3e104b4c3248a8cc3ae0828ce1ccbdf7c1eccde28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h941f19d25438839630edc32fff64bc76ce675a64f44844a56d9e3cb4d10c2f4f26315726a42b887f482ede6269db8a6e7d5824e56ffa72383d0621c4136f50009b0818b56b589af13f8e4789df092f4d2eec73107a429102aea584002d506c5efa43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97f6618076f23e2bafe2aa5591b840a64b0aafc0940b5edd224628f02c68a31b5f466514ab07172f3a4729d3861caba49894333e2694f278e6586da62347cda096ea59c49d88b3efb333eedf66dff0e5682446822b9ccc5ea88a999f41cdebbb1769;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a33abbf9c9f4ed57da7ba89f80cf5e97de6122f3c5628e3e555a9278e99402cccddc7f27130e07dad551f8d1ca2b4467387d8f3527735f864b2e1a0a8130cdd015cbfd9709ddbc06b94da1fd52f6d0b720495e7f7a61a40009b0ab7ba54d3ad0e55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1be0b21028f254de5349282bf087c48618e2809e205eab235b48159140fb64708572e9cee30282c8629bbeef55239be818cfbc211d56388c4caea6d766bc4f92b2ccb564a831aea6a33950f12c5f47ff3b92c91b629ddc7e1c2fb65622d7d4c6a89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8960782fc41c6422f3574ae1d2f23cc9e4be16774188956d0ae3cda320298557189666ec53b5aebd7be0890fc68ecaef1cfd717bcad69d3b0db7487573a680bfb6e7198a36dda7b1aa4051dbb92956eabb5bfddb32c3a783e41a089646955fe82463;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47bb186eb7d0da821782658686bbf87d14e40ce6b311957944a86367c7c9b4cf2d593723f340b68a6cc7e23f436810f3cd9f69ccab0b72802888584ba87b7fc7da4cdb11c77f118690371b6cab998d3027636ac274e63f615d6b3801e4b08dcb6d76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h842989f960740bccc603b92631f2c31ae8f7ab4a885c113decb2b9dcc97291fee6117aec37a84d2ff039d4ec9375f160aa4b3eafcf89c8ea19e7495c829ccea3eec5367290b254b982c715ba5ec15659ef058512a1a923d5f9f48ef654b4d2b9ad92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b47ee4f367e940670db87459c168968f43e56f47c2729dc165c0bf4654610b5b740420b717698e4ca519cc3cf55417d5af9783717aaace8adbb735932ed9d6eb805cc49d8c0f76075c9f38b8176f5db4bba4efd81c7449419b7c60130c4c846de0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha56c0f4b385201237620569f5787413767a9e99c770d115f3e175be9e6953ec998cb04702dde677ef83cd76e5b728d7bb2722bdf06bef1ace6516bea6767a91112e49ed2c97783ed0cf71320257ee8aa7897c6d120a490684d11d218867888e639e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8859965e119db39b93c2c01ef1370c0f7faed51524fd0f760beb251c42ff8ed0612655daf563a7392c441ba72d6a361027c645e5778f67f5f5f3aa921e90d1dbfe227c4a9b2f356e3be94da98286e72cb4467b2bd2a327717d7e237afdd82e9d642;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha82ace6790dd5c1bf90216a028693eb0d68960d0829d3bd68edb31cc630bd59e6cf95b46eb77a858a6a379016cdfaef68c477cea61a98352ebf5a72fec366182b28ce07cd41e6aa26eef050b16ca9eff298af194d8e291f7db58a9781ed3bf180724;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h179c945f20b0e1fb2d8d20c5be346e6d34862b92585ba0be30f279a9abc529e63b4fafcc0ff7bcae1f4f819e5b17a6a70a3479ddb4cd00a2495b5934835393d41dd96133f0b1402b9f6718c211ad9e0f239e07ffa4da0b441d6cdc1cb79a00184a93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0aa142bea5202deea9a079596f775e11c3bde95b87b0a1241d13bfee4eeb885073fd8fa76891ba229dcb9b88382fdb00a2da0417dfa1d8acc738c19f097ef62341239d21c75d59e33922843192c158d471f96297b363661f265be67e148e7108fec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1398a8c073caddcb454ecd8076b4425f1f8b9d64ffbd194a29d2a05d3c6b6f4e8c9d6c7467edf983afc4e6b5bdc05c6029590794f3f700b2a165aa36d06ed87378ac11231ae6010226e6896ba6ed0d348248b2780fb5cac733233022f28af53283;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7a98f57faaa2f63ea8b28c198f7ed367310a06a989273f35eb543187a95e998936fb48892ecc0767b93a30164b667d7dfb3adc2a633e4e3a5d7118949aeff27e9b6a23890e4bf84aa81bed937b6343c66216914ea6bb2de111e743fc87863959426;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4907f896b89d4483f506b49ab3e5babec28b9b907c855a58a12203f15d53e09c5f3909bf0a03445ba7b9e7616d95947d21fa71bede804107976d23fb0204507b70cdb99938066391324ff14ee04774fdf87f52bdbb032e041570cec7e040801a5340;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1e0f54f03085f7222f85fbee2b4953870e759dc7a1783f5f1cd4845927610deaaa4581e29b9d805ba656b08c11467d276dfb7cfd01defde2faeebafbf1d10fd6af4a1e90a4a6bd1cc874248c6c5f81c2e9ecaf6aaffdb5480b134cdf1f13923b172;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9abaae1074f2675f431c8ac96689bcde9bf308aaa5c7d42a7593df8b1b11f1344685e4fcfe6501d484c243c614555cd1912a2d35b546f9858e3c74be27dbda0e4451b9b9fd754414a1d3d82ca5d0a6aa89ad999c6e51311f0d068fdeadc30702e13f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he23629677dc83c29f33febe107e49aca1dca4086a6f9978563c8ab6a132f78033a2cb041190ec34dcbb70e0f670e7db300b8cb1a51c60665c1f6b54d70107851f57892c73f070751d79a1f324eaa91c044fca326e3556d95544ad25f3b62f6154246;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd07dd4aff853d07b4e63169a3caa200b654bbe737373493c38cd452317d1836cee85b0fa22b6ea9041a9bef99b68385517fd21c61a0e9588264809e99b474419a4df2e07ba794d06e8050637ae99c4e0ba1d938601e35d70924ce219928336b9d5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99988de12515766835ce49c72bc1a99fc22cf66e7aba74ce752687e63d28425956b9e2d54bfe56a23b1bc3aa356515676a96eface6fb8d3647e235d3ddc6c418bb37ce3a67d88149e22b9e7cd401b7455866a5169bf3db9530560847613b1f69c248;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f6f8d3fe45ddc879d31503d0fc1abb3ca187d588dc16fc3d698f479b10f11707bfb3a8fc6f0eef963098c77ae7a6c1472952306405f9250d5b288c3b50379e015656cfaada817ff3e69bb3cde7315c4a7f1c8dcfd06a71adef3b8ff00bd50ebd325;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd51ddd04040565610a94771871df73ce30b0c9e4e28191a4fe219181df4744ba781de3dfcf4c7d293e40862b4da6be59f10e67a75f9d369e52b9a0e37809cb9e9858041b84dd9ea29d78b0399171030bde2e8ff991e25adf8095f6be4daa9c6e4f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29938f630c9d7b1b25eee2aeb1f57d0171dd4380c1beefd83d46afed0fc160d6772e229f971615051ab2da319b0f913151888dd562011b41dfd941864625d94d22a377d62194a1d7995e4b6c82c6d2d61d136dd9be3f8c2b1425d1f9e8c03b93d3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfccc43abf585be1084f2c6bf64319f33d51f5c0f5dca24bb0c5930f944e5d4965b4f2fb3035d2b357615deb9f8fddfaa9a9f208826943d1b80ba514b6a1d68e7e458df965a065090d8afeee7cf08fed5dbd2ca28d8e30b57d9b697de8d53a7c80143;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29b32ce4398bb937db326439beac0a0f1d242bae98a9396b9a131724c08f881ebf9a93f4bb2fb1ffb24401fd554252623e4d4e4c5340521d1e14d59bcca46b9f090eb732652bd209cef87fa2912f802321bb0819b9862fddb59a650d0f90d273a5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4680739654e95d77a8a4dbc803875ec1186c0f9bde59032e29f1a4df37d1635babe467a8ad04af964f61f4578dca549e42d26199f0de1998164e9cdfa8e9e26e17b952bd3c14d6f46d14fd7af15b3ad74ff36fbb1605d3d1dc843e58f4bbc3110fd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7292804d47755be2fa7beb101246d37b0225496114a1ae03fe7cae4df6b02bc0649d39fc640f600f079c94cd25d28123d6b0347a014bc460747e1cfcc91ed5d584751aa09aa09392f5845e184b87b227936046e75431373abd38748825f67724cdf4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb230344e2c63d337c3e72b934c65aaca3f6115286d0bf894f5cd7e3cf820b21ad0cc9221887e4dd8e286df1972ceb8c560b3d76f5e120cf512848f94f1d854eff58dadcb1e95099bdbe0040ba9953571e4b5fb09ba5b4e5bce274516ca47fdcb117;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f3ac672aa161cdcd7663b976d322c15402c83e190fc47a0da1b1fd80e19f6bb84487c5fd05b4fce00f39e698d5e971e6eeb5d9038ae9a066b586dc112018433964f4fcbb3ef443bdb912b20d6a75c495d0290feb5424fe73b220472ada02c562586;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h287a5ae33f3219fd9e3075831331a24202c123d4949061f88b91701c9cb9ea76844c9f0a4119fd6767d102383d2e08a442a2b0b2b1ec49cfd394561b2424ef40a0f4d27b4867badfce4a3ad26dfb90b2e231a79f4996ecf684fa8db08e007ef964b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h187f1d945fafc459d07cd8759506ea819541c77bf41c8afff3198f5cb909b3c739a40f044aed10370071b069b6fdc52e2b18c21ca732c1da954880065a843b8f68264de7b74ee1d3de979bdc634dac55149cd1119182e9330954e30474962bcb77f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8d40cf711d729390e9f1ba1a763c45e594ea86579e7f43638028c2843cccbae0978d6796a8fbe9bd43a50e7fa087b50c1607aaefbd8164fa755c348531fd5f2dc3b30f8704566537edd93c0397c7ef217e826d22c4d501f60b0074e828c3e1e6222;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76889a47420867f4e1cd525563ade0f6e72afaddbbfdf699281382dd96332cfe1e84b1c6cfcfa3f70976a8eb59c5f3e0f9fbb7318ce2e58d9d535fa9ddec6f89fc45480fb584f3335eda5451a35ec48cfc144c1a550513421e9f8f553db685cc8842;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h249bc5786ce34d98eedcb0f08d029ce9ee71b7f9e93e3a4172e7ae1469acbb6e47ffcb10a888fb557ef217d9d9c01995df9b6ddddae15393a5b3da68cb39b61f953d862b4677415904bb409e201da34ca9e9d29e237597af51422422d11fb3f769a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1971006fe5859e0c2ac8f09bfd899b7fac7650e57b573eaccc2734c8ea50170dd997abd0ba442f09e8955c100ff3d8649818ef1a4918130bbb872f133dc36df981782b3e1be05d5ceba94acbc5804e3fa6c77df518f99610e487f319e436023b54f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h339aca65a1e54ce642ab2bc42c86528f0a7dc42a8c1fa76da84ecdedc56a35f82c8abb0244e42f08a2874203a4fb609e4f81cb9274c79321eb49638aa356f59062c8be80d98c5fe74c57e741be41a9980866d4e2c5c7117dd48f2ceab27e8f5cc9ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1f23dec931251a98eb2391968572fce40821c7b93a9005a4b21fe8031cb3d1146eacd9bc8d874c5deeb166c0b53060824fd86ef30dfdae21f80cd8e5deeceecb4a90d94fbd7d8cc3366b791a405676d6c55add53a4093807c921696e080e279734e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd6d3cc8a9976e5df0359c5fd6b64765053ea0778b77654b7b3fdc76b8dabdf19ce6c4783d7a68ff32b840d8b898ad1b80a11945957f59d0f6e72c79efaec37e096017d8a215d19cf7caa0176068e8cdbab6472aa029819c0fdfb8393005d101dca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he69d6f86c85246bc65329a8654d8138a6b473355d75b76a1c46e30c59645bd643f6e69e1e92f3fda67cd6971074f6952c75b6e5bb9b58b10d084472c2987cfd7392be24cf76b2cb000355b5843ff3085322ebc39fce4b8341ef122b635f74d701a8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68f66832a32a6331c27228aca6c7a26ff2ae3eca3781e14b51806b04e7a1e9d6b2ef499c2b97b00eb7bbd7f0cce42f30e70d1d1ec4c33b4e5a0b22b732966c87f399653e4a6e07743d4719f52c05d69c10230f9557e0d0ec056385adbff06e5b703c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf33126f402113244970512d7f1c7613fd2e1c69ad630e0862d41cba14283b6fe0403b4a3d5bc493802e39930b92cc35435a1886f573c9e5674cc8b656ab01adc1a5dfaef8e0e56161dd2f020410234c9dc2282c0107f78e4688bdcf2db8b03ab1831;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5407a3a88da1c6b6d84fca7760fac89c26e087783d3c46b230ad942ba36215a8ea49129abb838256c455ad0c2669502bf1c6f5a6674242428b5f40bee84abda50f4f8ee47c59a0f874aef62deafde961c3596d5850c00dae0618bd07121584a1f18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5686813d9b708089aca5fc2959f1346f3c52517cb95673e6acfa8090a53a91bc1b489d8c51509ea8ee3d1725b47ae56fb529e53d15948125f9dc3bd20e0e919cf92d38a296a02c56f78610f73f1200ce86312e4b3bd9d529fb02634318ec9cc0adf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6d3445f1360cb3380c94012431e808bd6d11899bc4fb3c6d43814430c1240a7b1dc6252083ee23517b68c18693b7cdcfa5c8cd2c8f28d5c7c4b26b5d4ca63593452a85e22e254612e3235d02002756f4e011debbdc815e301f83e53895a7e0b3c9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dd29ca6760a9df9ec8bfc2713a5707513f5f0c71263d6e044a558c6ea447d585edbd055ddf5f1aa6604a6c518fae72aab900e35f045d8379d49f8fd0505a731ee97e0eb478ec23836de7e4132bc6da95c5a42f11a9060118d81042233cee2b0a9c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d1bc24b51624cd92e363d928021daec0a447304dfc8c890d8b461d98b63d5ec15d60076fcb3d9d14d99a0be5be2c3037ccfaaf2c0d8ff3b3b641def4d94658e0f7e62f95e8f895f86d497a53565a866aa29689c7a7919bb7a3b25093a9b1b65f1d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2db58f8fd2a95925213c5bef150a0091db8913a3d0588de6779ecd20e8fc01f47cff47f9930e3b6715f8c8a5600d7b6fdfcd4073e1128045b66fb8c0aa75f568caaac942cec48ea4996f1cd9d384cb117b20c5eca7b4561dbfa07849d120f9350fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7637da97a2560e142f81398ec8f9cf940e2bfefefcbc4edece2a83e57a566812cfd789fc058972e952e60616530f8dd02920b54313e91efe3bd0d924b81cf1b758405b424ec27242c9127b4b8c2109894ca7645ab5c666c0926c446ac1d063f123fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28751a180c5107957e71a84578141d140a5966f027817c1e78cf1c4537b6e8f2634d3b233e6266902988fc7cfca4a32d6dad7bf2cfe21d5bef487655c9e93ca0c59fa9402b49d78d4c6c2f70b36f1c3cf95feac00b9440e755899416418b01a6198d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebbea980c496fe7e556329c08474a882190bf546a1fdc82288d4bf5e65cf647e85228c01a85afc98d95447fb7eb6f5723d19b07cdca951c12d06a663f7f760d4ed7b5602db41ef26f3d4458f6c11c41f6d133c8ae181c824ebb32d4e331bc7b48515;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1825c1ca82f194146b212fc122099cefba60f2db1a127c5bf3fc585f7a3409326b49766f933a20d8ec046cb96e877ee1df873b00e6866ea781c72d20ab2517c7017d0020f4d350112ecf4d75671d2e36a3ed84f123882f56540419c0b6602b5776d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb844d9151fb87b8f0837c83c8e5b99969f7432baccdf871308a9461f353261d4ea3f16c10cb8eecfef45f92d845f44b6d2eaa94179d955c003da4218c653ae195985c4366418724d04653d39c00b0834a3e2623b7676611bca37534673e5fb51b92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2bf72c84277f7c1594f057a603ab4d0fb4324353024d6d7cf598d94d902c09f3a6904ede9b185175c1697e8d3543bdc669d67ea8d6a55ef8fe5d241f8ed117e56b7e30a3a130f900d1f8de7366f0399d6a6279a572d7251c0df5c52b4e7219f3a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5caa64a0a9e61d1c78b6615ee645f13e4ce64139b15365f42274f4604fb6ab91abac8b84d1cd4a315a39f981152cbecddf8fefa0cc3339bb65ac9065b4c1dc05b3751d2852126a90eeea8a1701be95f2605cc9132e1bb2ba648127a9329fedc33f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9c5432bc7cdca706605e421cd719006e47fd4ec61cdbe55365a217c00992dd2f19c60269157ef7eaccc2696b1fcad255cb1e486fb525d8eda78ffb6f15ba873839d3cd45a7a0ece08159721970a4bbeb5564eb183e4abd83c1ee6919c612946e2c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha856dde104882a0f858c727e192b3e6e7034df67bca114db4ce225f0237bffb3cd77ae7d1dc46a6552e3466b0a63a3827e832d10c2d4f2b511516d9bef57f43a010ae37c046559610af2c681136768d6c8679407e796596a3ad602d1aea9d3637404;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26adb52e40b7262ff80fb36c297117cecdd775b531291670234ecc715a6ee6dc8e575586df47ea64e6a8a170a79f25970674de28bac39d0f81f9af81245ff356c019b346b7be12dd288d19bdf2258969a412d146324f853c53ff06ea9d4c98e515fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5e12dc13caaeaa52b01709bfe0b503c5f1f667ef78e7cf528f6998ebb9480caa53ca8d8ba24ee3a144b195e80165d5f921bd505cec5c25826d16e9be9ef979c7cfff388e91ce8bc61b0912c0e921d9622e622607d904e486e2535e38b41c14ac73a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e27f49877de4b08cde651f0e4ec3bcc7e5aeee83c743263a60a215d41ed6de48f2cbc39277b8e675f51a456c55ef026082283c8b6725b108860e5fce6fd48e638ced99b0483b3c50b9fbd438a39233bb2697596df77e1cfc5f74667482f12d0e25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe48efdc6db552516a566b30a3243069a25bc06aa953fa98552e039584ab4841097735f53d4a854573320e6b9ecee57eb17032c1de90ec722b342a9dbf9498205daf8b96e07b545aa00a3de42758a79f81e9610e6a76905f2b33225d857d42a75230;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7d5b5ce7ba211681fd11a48e587d126c0faec5c5434b434b79de7832aa03bdda23993af4314f3aa6a0edfe9d29c783cd38ba3fcaf3dfb3e618616908dce0a7647d077e5dc17af6a6912bd3a845d95a93384b7fff5315fbdce87657dfca9a336a66a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0f20f9fd89d01b620aefa5ee43c683a1ec5c5aa8253f859ab778023a91a279b08dd58710eb451ac273e15dafdb53d36893d8fa985c03b32b032ee9dd79cbadaad024596d137ef1542dcf4039ac942c0cbe110f90e7341aba7813c924a5208bde0b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1267ca15f5b186be26979ce83f1242b9f53f9578294942f85d65b2b0eb2f7332bcc9f7cd5b32dcba290b5e2f1aaae7b9e472d514bf2c9bdac3c0f0b8a32ae1978886821a6e6ab6976583e34f8a753c906b360986ec0d4cf873db62c9cfdd95a8f095;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6a2aeb2be38ace5d97a3760deb78032fac5b3b07b1725651d9f4d557b7b716f175f95beed119823674897343a45e45e8c576348521b883ba390913f6b35443463f65af8a422c04a584596eceba060a85ec3e6f657b99d4ebf68b7de399f229167;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27ea1b2e713e0018c559a61fcae5429362a7cf3f84d2182d4c5e0852d323d617ab6a2e0bebae9465bb02b1de1c6c83c3c308f862251ac7e522fb593196dc1e950ee0b40f60514806c995833b90d5ef719ef048d8994a579a229f92a6157a1965bea3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ecdffcdeb7c40d519cf5e85dcbc4eedcde64ec43f7d17e80f89cb42e0989a22e9dc64c65f5c188c9a6d1f2e6271bc9d301da1eb5522fe858281ef5b1c10ec1a4e1e94ab1bd68f8b0252bffb29a08a342cc51f24dc22ae738515f03f353780f36cbc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h797f3c37fc08e40071d796513912b427f4be5587329f5838b46c7bdf1ec1d65b7964679712ed9027292c115c70271bc3865d03f356dc6d23a2e7457eb73f9500600220ec75dc18a3648c3152438b290ad7c46543156368c6c2014c5e959eacc2b9b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3937b64f3fb5a3b6d8cc47e2557f605f5632d66d8818b008e0ef42acd63cdf5d364c5e7f7b5b389afc82ef3d800990a6e7c2a08f0d025fca8ae165317ac5fb5aef527748ff8535f45b92682b792e14a0c28518b675441e1422237437a941d98ab762;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33c63e8fa8dd206fdb5e4dd626fe902f1dc45244de30fa7cc10e75116feebdcdb4744da75adb33fcc09060baf748f0a7006ac6f869408950b13cb4b474c490098320420ef431c1559d8fa86966fe78724691d77ff5b4a4c6873f671335f5b2adbf98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h433d2e5cbe8bb22a7b2c287bc5753d9b7decc1aacfde6f10ac3ded1e7e8f6025500a94e5a6ba45a60e99be901414953dc4e6a09d638830d670f2a02115ce44649f941c5781d647e0a7859f94c326bd039a5a217b1c42803ab8197a0b15bc4d233f97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb11f51c8df046f9058b1f8a71f3666f83244149ac2b8d1114d1795cd7fe2ce897c68d00266e0839e3ecd0b2ec989b58ef552d520e38a1778491217260a38098cb8cc1059415542aae1a85ac10d7d2fd5be79cd99a6cee56891af181c43aef3ba4704;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a50dd12e1d8410940bd4888900133354503fa99096c61c06b05edd40792105ac68f15bd8b2ee8918c2ef69e406ebcb665f5d9d9b2c47b4d53ccef0a3070789d0689288bb019653e81bf8bc1ccafc8b5729e87704f494201f230f4ea9aad406c2355;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a45712e59cba11bf7262bb346f065f44afab72b3108b28c12c4642d4d14731335d202f7561ed30816a020f9652763dc9d0835c94a53462f5578cda872915ec60b85ac23fe95af44e00f6b758059eb885bfb5177d9250bdd04d9b2bf99bcd3c0d07c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc67543641ba314b16d142545b20271131197c1b311bea242fe1edfa25f2f973d176427cbe4bd151a27bcb0a0d1d0573c1c9e63fb5d0a93c243df41743e254ac9e5a3a1d9c0e4c31763853458d9472b8caf5048425355b32f4f2346bebdde152a947;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddf441d50f739d95bc3bedabcf9457ac6dc42d4b25f7350242311a8bf2d822e21cbc876b1e0efc4a71aea497eba9f2ddfdbdbc80f7f5a9662b470d8be606875f2ddd905fbb9812a07b8667e1cfe51336942a05a26eeb9fa0f3b35e0ad4daa1c1888d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h994d938726a1c56973d2347a7c03ad52ebe9cc15513d9299b4e16092e08fab8df7c39a9aa2590293c26fad7c8ddaf5d4863ed372d83da6c92e4312fc370c73744165465687d157f66d6dadd8faf2e76c6d3ec72bd256862a7938039fac28fcf2b125;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23cf13df3a37a9fb38922ff1c3080175739257eecd9b291d2d65cca68c7cb83f8927e3392c1f3c5379fc5bf328b9a52595338a6691b292857152b9f6fa1fb4596ae03e44e8f538779c45293de73692df6d7414d3d40be2d24478b1022a70227aeec9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3d92c593da8e94a6259663faf43e18810ee5e0c9af60ce6160e5f6d1a6d37fe26763d39f2e852002b383a9accd9d91c426d988e1c00a3bc0fa7a78f2c9041321fe1f86dd4e6bee6321f5c32ee2d6e8bb8dfd91d3b3c342c701fb6c2f8cebe584614;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd850ce5fab9e16946f8f4b7c39cb2f4d4a03e71b29f3c7b171dafa41942547e551988b38e52993d4d8f78dd6fdcd839a8d479c23f69e6a955246acedb245a3371093e35fffecdd63016e497cf351eaa21e6705a84aaa98b5de3f8c60e3bca4338753;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9c5c54917de39feee6ab3f06ebf2c022c5b5cf581f3a4d2b2dbaba842b60fde84e27ff689b5902f3969d1c36a3710d861a1469edbfa9023558c116fe6b8d0115c7c962773270abf4ae54198ceae247ffe048ab9b8784799424de412ba2b9a8caf19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb73951b5721c9ae6302b5f3a6cb187e6eb91d314367528d94529c41790d016cae171409cb4208380f0ae7f83951e053585480a4e4b9461dc2d48171fb5d1342c8d253849298bda12afa17e6b34f263b42b4816863e6b8c80a94bbed0d82fe35e092e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7eb7149924376383d5103272d7f86d1a4532ec735ce8acee3e7fe6565e43c71d5a80577db8d4d0811909e2974d79175ac74e229fe8362c23dec42fc5b1233340787a3e62d4e04a53d192397f2de2f707fb218fec59689de09e51f1dfc3a2f13ff48b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e739ad3ab5c2ed6256c999f9329fbb4aa79b37c016f1c6b90a7282624a90fcef422264262e7d43a9641c6b0cfb69f2ed25f267dec848f536c21a2224cdd95e6faf0559062b44b9130477b71c1c66d815e75b18125b803abd2aef42b20b785127f92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb929e27ba86d37b915dcc96a8a4b04bc349f4ec7efdae38135f259b1361edf93183bbb9a1705afde0a3be5c1403359314d30dc79280e681f22563c4c41311f32ba4326f52f5731ca564679373fd5b97c028f89b59a3fccbe407fc9e3fd76279ebce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haba2dd18e86bee7ad5afc2d14edd0afd986a98ffd92973c8b1ab3ca5ac319b428ab7e8157fec60940533a10fd6351826514c42e3b3c9675d5d8ac3b3f1cec86f955764efabcd2910653188b957f294a74fa3907ea0abb77a0e8274d5fe69313a9d52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haab59cac042e84b2967a419d500875a985afb743229c7e2528a9e5e7263c89935df9ea4eb44041116dc9392159fa11fa3365c23015389dfb6397008228b76e1c167179184e01f76fc2c342e2a32f83ed66481cd990486d90590456dbf373e1d1229a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4789a9b7f9524c8a0447aa656264f5b72c14a9722d1af4925c66613ba755219a397ade320d2e54ab939fe9cf66f19f9863ee459fa9de149ac4713cfec80d84c3b44103a99b71e84a154f7e0fc3b7604f79a7bb3c8e98ba07112aeb61746a5c52299;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6d408d0411672d7191c8e5e12822af2ea833522bce6ebd78345731bc73d439b560879b606a6e541b05edc7eabcd7540861a6be6ced4ede6e9790d2f1ddef1f1c34f7ac5c0df00c2ec3f7d9a15d5fce6bf3bc2081d90e560f9f7d47dee2f76040b2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a06236cdb098826ec307d8d59d11c4adfdff7437af8a13666a7db515bb09246887c6256869651735b0b477af9f25d89ac9f658d726181f6ffcd89e81b1f99871c2ffb872af5eef9e366f5fb7c855cc36a4d49b9f3d3acd4e748c69ee504864a34e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h277052778a208bcd189c8081554561619f0e5587061785c763828b03d823bcdf89abbfcd52ab2545a5dee98881fe967ae203c07763a105771b5f44db7024d5513c75a9763e32e7a4a1211e5d6f1253905ee1f1635061d24cda5cc5199561463a9c97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe05db81b6814ea88d0c56a145255de2d422ac4cf09f22b91795659622aa480f92b5475dffc670b3d1bdc8b9e35be7c950084f11831f0dc46757d258071f0a2024fedaa528901572a6e091fe8ff20003f71e59e30f450a305f325e50dbb080db5385;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1bb51f363d06290bd376e4b7a95ab874ec02d412929f77940ca9a27b69ae00ad125b723b3aad52cb71d861f55acc1a252417a5aac972d4b944738dc5a3dbcd77e4fb8f88e4914368fbc2c0eaf4bffe21970590e1922abe3ac1e8a520f736080427a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93ca7d7a5f5a94932bc8e2a5a417c82b22d1754432688ed7047c7c1660a9a18c183e4f6d0b823317f3bba0d70a344cab99b58dd2c9178f751939c271cfe76c3d24f6415c1b4f8921ea707c17a3f84414a9685c130d083dcf23b374ff380322a6a69f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h750bd9c77c1722fecdb924d477405eae455787444f95751583e4c6f9db94c20e155f0618537e05deaf8545c714c661b5cf49848e5ce902d95fc810337911085b7776224eeafe4b427abc6c0fb0b4e1e3fa7dfc6d1e3f2c1c50ecf8661491f0be94ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52d03859f05cc1277011a66edef8682b9b7184fc9a4846b44c9e40dd487c7c8b99319b2f4d43bc9b320e2789f515d9e1fc9417160369b7df02258a3e5e3120bf83512d91e77c37d6c3910976b0c77402f6ce39b57a42f8ea21907df47bec06ed79f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2151a4bb18ec5a18947c639772eebcb65ccba6cebd48f0adf937e06cea18ad542b2e5a7748b9d8ee1da7503d02629bbf3a399e1057bbe826999d082020fd5d3969ff6af4062d6d84ae40318e0589871cbf15685d65417728b0966050b270f15fc36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88114f8d60ea73329c8671e638d6f17dcf5a41d2d25aef730ad111a3200126697c69f261dd3f256fd1c8e46871afc7d930a1463b7276b5d2f3a5ad3526c2eb95273a3f2f0392d3e3459f6aacf131ca64fe8517bc32afe731f6535d6bb45edf5cfdec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h762afea59f01cab7fb07193140d786a29b9251149081f5297d61fd0b0d4041b7c91e51f8f49a01e6cf6e5d9f83ce23ee086ce4758b79d75250fa81d4e7a61998001cf41d68b08444e8fa6446abc3b685e83752465c2722e247e0549a34b7dee18857;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9f63614b5a38b42d5d59975582b8a270c59a91973e5faf516912fb60e54808d9d210bac2e2a516a5ab31f95adf177114612774bbffdaf5f2b2d0a754d92dc3ffa214403a5d9a76da3d7e3a5f91ed52478580edf7c63ca506d67dfd73d24013d0b8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96c7b6d9e09e601f9955b72eff5ad7a5b526cf259a25b7576219c7b5cba259b9c4b81a6a7e39c2ac263ec2c597ea7d25e4b77c32862a6d42ff666b237f7a2a0cd2ffa54f0cb2cc958f9a39a3c5548050841f6424407eec51e2116ea6aacfce12df02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14ed794edaaa921a54e3429ab1d465e7ea0a4e88b0894375a2995579b919b87661aa9c4b104436c4d0f134f53270dc669f8203d347d338e048a900ca7ffd76a1b7c7910bb4931b884a84d6a1a60c90a69f90125642ab16fcd366b80e9db71c9d12fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa10657ebbb69a82bf3117d913ae2a75823dee588e20ac15e17b64044c4bcaeac077dc018cb015c191a229bdf8fcf10fd7215638bf5b6d574a6846674ef5e2311a1c127a2e12ee32ef356f8c96e2669c329793683969f07d3823a6f91a4b10a0ce41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h397be9e0e9180191675ec2b308ff1014c5a6b51f6085e751b643ac5bb620f81d9275cb06db6990f39ab63e8ba33998b1472d14cf13b0db6b57893c5fd6fdcc0753683c472bff49122196cd1188160fcc718a98e9d3e92c61477d1180804855b21a9f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h844091bba59aea996c0a515219a70c57028d7f288609456c4fd141fbec40f2591ca06bc10362537f5aff0af42b338ab5f12d4a7a0f2620393e44949bf22f7d742125770b1df1f0d0ab27fdbf02de9a6cc73124cdc49d7d050078dd863a584b0eafd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e12e32c7bb28de5fac14d9e4ec023adf95161b001fca24066eb6341cee69ff027841165f5d4156106813a0dfa80f9a9ad2aa2d0fc46a209e5389ed39aed3183c1e4846abc12bdf79d833184149a0260e4c839b5a97c6d2b92ba316121481bd1ffc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a135d0fd219052fa94b3520b63b63ce2d2a2b8c6f62d81e61d21912381beb405f1da6c7f6b992f8603d78572b4d82393f633409f98368388037d706f26deeb0ea8c894020199e46206a66854fb802f0cddce2dbec9b0d32e6336cbcfd031326118;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdab09b4075b05eb83a030fb1e353803e0446edce210dae2698f565536ec541a7ddcad693063620d3f4f80da93aade4e814b83897bdbf0a17ef9779eca20edf8dc80e81a2b8270ee5ee8ac2a9124d94e4784deb7c5107dbf7dc60a005b918b0a74dd6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3955cd52b2ef6d80e7d724fdbde147f5c322ce1768360579a5bce0c58788823c3333bcb99f21508057d9f68f696938b2ef64acd43e2817f9eb446e8f0eeb4e3f2ac2bc9ef0f65dece96c3bb62458447d32132a716a4c4996fd715fee2e7d160fa54f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dd9bf428b380104ac99145bac791f760d19211c71c172f3e274db888d1751f1f5e727224bba2ff32e4f79fbd11062f6a0887195f5c3ad0036c578b8e66089e17c87c0d3172c37f8a69702dbd308fa1a5cd8696b50af77e23c7f546a92b14400b3c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9f3ed19ab7fcb19dff0d840479c254fdef7d65842eb9f3b46d289ab902be3b2426080c10b3ad0a2171c0b0afe4730fc1b297c99f7d17ff7942bfc2141940d5feedd758589fb6db8dd22b59d45712e6f0dfa2880fe94c9b7fc2c8b9c80c99af01831;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha82ebc7dbe879795abfcbd6be6a2f8180b34bc9bb991aec418f46ff06d03bdabeee7f32cdcd87a4869cff307711c63a89ef30a3df5b67c825ded31854e5e63d55a1ff16fe3300eedcde881ae788b53dcd3e0017d525f9fd14a1071b66bd6f71f0b92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h877018a61ab90633e8ce59683d478f622a7ce2770e9a0880eba9a3a3946541c5aac3beebca4c918ec38ed830a17bad3f78b78283569accd71acf67abdd8b997ed126c8b0989407dd5d2340d31f62acc21dbbe5210dbb4b09ea4d935e682e5da984b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha038d6e56f1103b97383e9d2dee337ea97b18ae5a45af3d2e1a136daa9ea9380551a0bad2bfa928fbff968d6f8677752969f5a200971bf9184c2cc27ace46b09e195a23e2a6e983391f988590c79087c601556f1bf5d3e0ff87238197f4be58e2e7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4b7af11bf485bd88febd71477acb803b758b0d89c04fffbfa27e8475965ae7a62cd6d560be02d2189dc348bd43f3ea82039257104518c25ba0e575a9b115cd44a629c2a52a31d7bda99830070a2253216dcff76995a9d9f279769816074a613f597;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h537f19a26a5b7847dec20389b4acaf1971e9e63d02c24a772d79c22362329bd0ee5284f0dea5576cc884c1410caf88ac33e7b219a832cd2542135e3565b2ee91938e1d339d2fabb6f83ea2a25c3ca5e5d42c3b7957d8b23484b53ccd7ee328d9c1f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93692d5ecafdfecd93e48d90fa971b66061a463972ce6bc3bc85277d8abe5b8ae960b05d003cf3c466a541d8ec660afc0014b498387cd15ae2075537ba5066182e07030ea04a48eac822f8afb8eb07e2f967a72dd1fc23fd7aeaca706d8bc4dec079;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880a153202f1a8f90f3c3cba7443adbc58ef28703dc3e7f491a1051652d6f76951c9854cafdf0ffd8560eb0cc14846e0f8664df3d4bebe25a2c694a7437cae54fd50c7a0cf4afc71d19e086a27fb0bbee59f5dffc83f8d4113666771d1d56ed936f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a20d3df6ce4a6ed893eac26e28d3f5a2b25b79251047e5de932d80c04953cd6ce9a6e2ec4342511d4e4f7c60869c8d580c3805349a7816602d71d362643f7ece3b3c3d6e04f5ca125bf43ec1e3604d78d8ef18b0be26aa4a88bb8083d1351419b7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he96487c1fef83df9e4e48e4525c8041d2f0f98c37b9dc9095b676d5d76de71cf134b747b40835f0c46a3305927ce5dae0e40eeaa9b113ea0ecf60e11075223871725a273687c87e304fde3ae163a266cf1478f39e84bead3f8a9e55c5eb1881d0b64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd6e2e90673175e146a4c69a5a86e631a3c979fa955688819a20cbd4ed28d7e49641af8b95c38ff83db898a7a3cefae165681f52ec1ca11175d90b0a7bbdb171293c417cc18c5ed1510188033c9f44e35ac40fc6418e9e09a813a648026a438f59c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he866730bf4ac322beee71ab4ca302aa1fc9de9864ade0cf5010c1d63a1bb4e89ef6a01a25a9a78f64cff8612f71d1e32f56079056b06b0f5591decffaa9077c6581ff32d1593152230de47e06933b8aa9e58661352df542e2b7a68cf69219dd9f855;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3a0f52633ad412a0c1fd2d86efeda0dcdfd5fc67d41046ddaa6215bc10c534b2fe9c586b1c1aeca6b538fee1f2de7ce3810892450f96e0e700f97fc1ca54270fdba2cf9ac05a647e3ea53c0a10b1ae216349729594833c510a005f8bf7c80e49c15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc697a2c69ac2c01e120ffc5fa8cb71c5e54a8447d65498e3e80cb004b3c51675dcdedc2a78fe4a32467797ea3521705f06dbb8272b8253a8c464e1f062a6188bf6d63f7169b5b46d56591c8c0ae15698a47983a812eee67c77df1e7d89d91e1dde89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8912c6b7232690ba294131f7080e881b1e083b721cfe59acd0c79dde4accd43082c471f7e3ec9943d95c4e0b249dcb1912165328f68ce7ffdcdbfa61b4a94dc8ff3ec7dab3f648e46387702ab7f54b70b8806ff97a56f2ac15cb782f4e59054fdac5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he478c15c2b44e152a5a9ab85b9765724ec9c564954d3da84c6d08ab450e0b7d94cbcd814cdce854d1f2b5f92103b459e8fb333815bfd478c6b19884ab592b08f890d477dbb9555338e63a111ea4fffddfb75a167236a9f6559c0ee448bc8a1e17612;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h291df69a72eada78ddc7347ffab428fa3751f929f6e3a5d36771d501093000f46614c960778581ce3fe9c63b096eaa4fb6a58b697fe1d0516c3d287476d6774c45fe881acfc569ea6fa7adaba44c77f32a9ec157095d77307d84b64447431f48078b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1d846b5bdae91dac02d857b60c8ba2b9f519aa54a747f86bcd40134fd26f433897531182a8e48818ab610c619db26dce3d33ab2dacc726d8285893f08a699403d9883584f8ff45e2ffe2b41293028fd3a543d4acefc4b03a2775376b5f4c8a340c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h434687fb29f975b87cba38302333ea1d3cfd2ffba8df6d573c6ddfc16b7226567c0ccbf60de68c172db7915aa6470377f32d7ba8f189d0f9952b4efac2ff5d68120b21b221a0ca6efdcd113c0bc9e2139a7ec61254b09e7c32210bfd35ec437922c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dbbb895f468a3041961b5b406165a813d88bde665cb16718278bec2676959a63547ebeb38c1704a27f0a87320a791ba23be09f2f1a841458f62f8db9735eca30efb6600046e000d34e40e125b81e9485f22b97dfd80893f4e9ecd5a9e62ffd86606;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h506170980a78ebcd5a4886de6db77cbe4ecd4bf03cea356a1b04f53430d113775fbaebe8aa1779e9d6e7e5adc10ce1f1280b0479f96912ae6ec16f3d15979faebedab6f1fd6d30ac1844d3066c7b55785fa252421eeb5401bd2ec791de5c600cede1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1415765f8081236c04fbbbe7fb12e4d08c8aa1fe9d5f6270bf916dc31cfc05926da73f9fc1e80238c8abbe7b4f6f37dd81d4df810312d09c91668f7767912bab99b29f8f268b6462aecbf4361dff40da0b907f04ac57aa52d3676db39e476b72fa1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9efe28f2bbc1195922c98ebf72824b368437273b84c1caaa9de4d2960313bb3cb1a57c8f34c50b63ded516bd65d2b5c7846e5ccd7e7859ffce98fa026048633641da60b6c5de47a2035c0bcd89f9272a7917bb809d844da41a26b091a0501ff8382f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a6649c66353c5f038caa26b5b2841ae986ae3bff4b0c80fe902701aa43bd13ae0681b3df7e8c6e601bafd7b0a76b1569d0cbeafe2814cf215c10ce106bc7b69c3f62bc9aa50754011cd21c85478bf078a7b675fd9a68e9686da3b6a698eb5eab75f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6747c4c5dfc379509a95fa25905189db0ce6908fd849212918afe10bd814eea1d158d34367033463ee5c4a7d9419187f804e4d73ece013c54c3d37c0b97a660c156f3c2e4788eeffb30199bf12f90395cd1dbd4f950e6e3afcfb4828c3ccfbe99de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf78de2df1ba08bf845221517a16412e9d9c7b81af8b22299314dbf872007b5bbf02c56525f4e94d63e0f8bb2325eab5ed11aff344aeb4753b0de41e8215c99ec8589ac6dda4cd333e2a92c92338dbe1553bf9720c4ed011a7e72dff74cde1b8fc9fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3f2869321d1c430c42652917a488267391a8321dd37debe7189768f87dac93ec9b97b10ef722e2dc368429d63b94d117833ae18fb346c93f05daa2d1a236ef17fc6dcc51c3002770670acf9433ebf9809cac26cc936125a48a36542fe7531e9094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc77289424959d229358a52080ee2288c2a7a0a82ef93c299e38bab755684f20c9d19f6a2c10aa91d2d57b158915a61f19c7f66ff1fbb06a98194332726be74aa9c1b7c1bd5e4958a7df7fef54fef0f27462cb5623e0a9e3bd7246a24d5155d693a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h426a81a35e754bda0e040cb7f198d1d5b1093980a040ac0fb564224435b6248b295104d2480a9f925794c8d89f7a74409ec304b58259cb8497bd19d41355214e7b542e224db4a0fec74ae73354dde3ce7c6d5b1232afc4533c86d575023c7e8466e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86d6dcd329e56bcb86b7e1969fdeaa71d748f06fa8684f27547ce13771356ce89680c3fa0b5a2e584d27442a3c3d29f3b2cde59db270ac6cf6cbb58776a5435ea5461c2bc11a5d8ee3cf57ca8b539d2ee00fa1649f0100b0ab001f0164d860b1ec0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36a91ba242f2d6e486247e817e60545ed3df31fe866e63f3e0a98441cd8ffec3c919cd9c0a4852947dfdbf4412a4d52756ce82b68c942c5728690c90905da02866e9dc824e6eaa9112cf5c9cccdcd552a604ea5fec54c89c44c775ca7976859571ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h872cafc0a1462eb1abe5b8949461f80ef23904492141e571f12c1d224325ef74bd67ae378fde9ecb5aa8ac50a75238718ea8d8ba372080805820fcc881a8f945d8b4c3fbe6e34fdf58931a4fb49a768e47fbf55fbdd1d6c36161819ae3fb0e462f86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc7c61de939a16ca08a60a2409f1d11f16324f9dfb99c2e6748a68e280e94b37ef7dfc6ae3088e24c3c98cdde459f32fa156e27e2a62c9596dbd7a1023e4f1bd186dc57abf8d3c41ec1882aefc11b8dc20ab41cb099627441b82f162a6c6687ca2b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd826519265a2c73d34cd21157f0565cf2ff0591e6db254cfd9ebe8c1cf7884f549da2129038c1785a9edf50113c2d492ed2cc77c5ad154aebfe8b9845a315631085d365530a3bbb0b642728fcc8928cf127522eb80368a517e6fec47b52ac27a3ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7ca283e9127b5133354885d81a08c7050ef3be065bf5dafb3ee5ab632d8285c82261dab2a8b582b4a36700550ae2b9d382efb2baab5fd8c21ec174c9655ad103d6dbe8cddad944d029b68fec0123124316aee7a6cf43151292acc2ff3a953da172;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec4660ef26a7376845a987e9f2dc84db3b0dc12197ca4950aba63052c7afb454494c89a2dced4499c5f739aebcba4f378c5e801977c7e33a94ec36f77d5e3c8c96ea69c6fe589d8545345b72eeef1477d8839281afb55eda9eb120b5c103b88d61ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4317c51e58c9e85f30d147ea91061fe97610a6876a71f354bc87e47d87c364c26582b3a69c39259aca53fbdd66da70499c7f9069c474c32cf795cf5a6849fdb5e023b55ad84947721ad78e50bcd81b15134a59436f2d9bb014c7dedae0f86d4ebc87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45797c424a784489fe76fb6b674472c4b6e8d19f6aad5350a8058519e30091ba36955b3cbfed3d3f6855b084a780664a13361329bd92ca66772a3bc9c59118a316f5e7fb68b9a530fa338fcf73fe0eb2e6c0bedbcab4069ba744167d21f4e7e6e476;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5fd6592551ace08c433a1a11e18bee92e68da249a57946d5eafca97af2ca4f7fdff3ea94350d8c174a9b3316bebc09516706c1cda5a4ef2ee210e597ad3442e020af0756bf1dcc7c09391fec6de3663245a8e881ed36ba4861021c4f28f002406fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20df5605a36b1d0ea67e5a9b091a58a11345ce90da7bf3a3d42a0b2b93aa21578a7fb79951499f6c9ab87ee06ce6dc5d00190196553387afeb23e55b69fb4f962208ff92c49a3dbbf1da96d18710dea9cd80bd88ffec201e7dc8ccd6034926848c72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3197d54cb3359df94be1f35725438705655a96f93c290b4fda67c0018b8f1e106a2ed542e75547ece0ebe0e71efc9c59bf1ae8469966c892fda455fd8b4ed7bf88b87cfbacaf044fc96ed58695859db0d2e0c2f2ccc105f0aa1c19a23ac8dcf67bb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3b35c08a81e5461afff0b927aa3eeb84eb8a0eeffd4e51d78d829ea175977f666c4ecf343123e2c23729eb4eba2eaadcafd68eb67ea5bc9f62c6b1e31dc7d09d5ca5c2ca7b3294b05c658de4b5b938126f7effafbe18b7c37b1da0ab58509001710;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19e264128e69943fcfa7160971fcfab38491328c70495dbdb29277f448461f7beee4e4ffbb594ceca343959777d2fa160e1e3e16a25f55f752102310b074997f5a4065a568f6d90dccbf485da3a98b0382d7e2afe5f4c0ac5f36077e959d5d5361f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1849a67dee327ebdab47ad657dea4846e438a16e5cb3d01df89ed70a243ef0b42ed226f07ea7e764553b13c412c5c362f278aead8c0003efa7a3dc3042191dcdaed18f7b63dbc86e7e8bc2b7aa754d9ef68d9a4d3fb3f6460dafa6eafef7a1ab9cee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0775c2933714faf1407e3f8e73705a3d2303da2b652d6909c6725258ba78632a8bb9488975c0ea9888b26aaeb6755e529dd6a42adf0bc1e6254b0e381564389cda01ad738633c1e5a939138845b825003bf49efea8438b933d6960b622409d0c133;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a15f26f15cf47c16e15d13bc602e823608dc7647e32bf20840c846994571f04f873a1184f0fd70157907839e5b3bfe7e37cddc760c6336e4febda349ab11da46b6654dec9651587ddb6f6e1007b28749a5c2e3a237b48a03584c70d0ef03844e66;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69cc0e6058f2dd73338c159b611824933f314a7d522f8c5c261fb434c764c3c8e62b18cb319cf3446cef9301600210218d9e26f54d348edc7eee74710c21780227ec5770618234a6f3cb97ad6590834ed8e1149d9a671f21a6142a9aa5c0b73983aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42ce120445c62fbe691955df5a786d278de5a6ad040fafc2b6e88b1edb3f78939618539c1031ff2c3dda4040c7cc5442bf88945274f18b6afae2f956aae6bb0945f87fe4ccca1834f1ec48121c036b1ac7b4eb5c52085321561f6249ced5e1785ce9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bfe8a6ef59a68426aadf4d07a3ea674cdc31a909536d39e8464d0db21ce6224877806fcacb28bbfa178078d60ea7f9e214cd82f421f1afc03bd92dc107c5ec690a997af77257e9c0421f3ec2d8cd4e8d9809f42f43cacbc0ed45036e043454c2d8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ae53ee5ca8858874c0618f774afdebf0106a2ad1da813f7c3d3e548752cea296a6c90aa32e8cdab9fee04069599574184d237cc7ad28aa775689c70ede16fdff88426e7ff667042c4ff720c3476e6121a735bf72e53aa0f05126686f35c061b66e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a4681a881192549ff2370cef04e16dbcddf8d4ddcc37eae56e912f8b66152f01e7ded14e6afc6fdca8b9892286566e18d783499f057e2941c912d050969e1f55bc64462d9023d66471cbca7c8999545a8a56b0043c0f23334ccfc958174dc621429;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f7884ea882f49f403cd146616b6e355c74dfcde8420ff3f1d35d37711bdbc6fd6136a6bef2756dadff01dc3066f398c8f0dcc3ca726bcf4cbc7d1f9edd2557cfea8a5bc979466eae9519287a3d7dcadcf8e9fa7fac1da80dc90038b9c231f05ce21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf580130b7895b467cd44264e8b9edf93057ed263121c15a1795a06027a37a2e898ac028f407bb9746f126e3323b8dd22f469bfa98e8d7a2f7d77072ca66d758a03fe4adafb4333f3a61e2f88b321c11c7818c26e2d2872e88645d02d384585b144b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf27e25dd821cab35070f62df90b656005764f78130077ba6bd01a01b8df840966610d456eee1363af582325dd77534425652ca7837105ed43511986f503880b5af7bba8d25e9f07ecc6eb5d374501cfdca261934b44b3ee6eb44ca56cf1dd5002877;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h544eed86b0449dde1c0807ed363af17bad5df2aa6735c322f21acfd85c8c6916f4b7cdcf649cad96680249b1c2335dcbb84f71f0fbb62d1d28d15164ba58bacba9e23b3e9511e876093cb9744faf6f036e19f9f520e4d072d67d82cff66b0dd55639;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf22683513f342a7ba113b164c4908ccdba74af7766e3437320d23373ce7dce278afba6477d0b36ec7e8cd442fb39cb4d8678d0cfd83ecd8381126fb56ed117744c9cc7094734f71fba4630227b2a9d3feea2f7482ce80fb28e6b5f358f79e9e612f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c54e629b7cada54a7b195365f98b4d8d9e7590bcc888908cb51c42cca5dc35608e6646eac5f8043a7760f6a450cb95d7e64aea9fbfabe50d29e4f85c38f5727cecf9eb08239c3edfb633629fc67dca9b26f8f9a5f7ff75d761f83d4983f4891ea96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc05361f020ff6b3f8a4a571e13e0aead6814c5b422df6b4ede00d7dd1603463db102378420ff85c1bcc388a2c529aace8c1cdb3e4561da0f7b094d07a70174df7a0e464a975a7fad00372495f68d75d395ca8ef5ab4edfada548f58c0b1ca50ad0ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe277f549f9103d90c0874d337a3070e6188a2e9e69bfd4a35e8ad8240709d6bfffb69cf0e2935f261ccdd550b9021471411628cefb1e1cd7a3c98c8a6baedd218da3b0b500b96c0fee942b029b8df0e2bf24490665893192a1b9274c0e4b16a058f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7e4353b4ad4abb16f5ebb1113ea008eda225e505e253c9273c97638273e041d3fa0f24a2a2a66a44f498c01e2b9631890ddadf34a7180e59c60909fcdca59468a6ba16208c9a126cc5f527ea47b741c67f92762b65629b1c07ca467a9c149547d10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4c98cc89228e60e892848ad7e074d7566de01a8546dd200fe87144361f4d22a541d416725b013a3ce454fb59c8830d47e7254c4106bbb673765696fd53662286900533a74425f8a216fe7777a167d94ad2a2a5603f9ae213157e8129b350dc4c0a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h975e410d9331ac0bd93a4e64ea3f4e393687ab2f243d7bb0dc7dc53ed0195ded8c744a3a91e68205a4b779e6b4a5e2808d30482c01e31157bb99999ddee65ebd867b3525a50199b926cffbaf2bf3064688810d44c576ac50f417363e7bf3d4cad47d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19b9f5d25bd30e4f9c273d6307b274492e98dcf85fc0a5fdfdd2a8e7a336a0e6c4a2a56edf409a096f24e90aea9777ceff2e8ed10db07ec47cdc31934814f3a80e4696dbab4dd940d5ab34613de2437f1b3a7114c95bfabea4af4d1a85c2945fabe2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5139bb6acf11f6e809fe56676cda8bf8fd319fec4ea6be62acba93a64596c7fd57a83d61d3aa1b2da00679704c007866c40ebd0d35dd3b80383614a69ad7ed21d4db017ef73ad28681fa04dbb7a67fbfd10149214489e0993b9c870be05ed14b50b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe8d016b9ea3ad1eed864d793b678259bec06f55e60c84303ee7e6448772b3333829914a0a2479d51274674694c4fc76026400ddf0a7679e4c08d86be79a1bdf149c26cf075b830ba29361c4545cf916c7409f6d860e8722c6aa5ec6aa188b09a2ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67c0d800e149ea8af95e3501723e816208899ca4a2492ac974348f2c3429d422bfd0d960e0f69f59692c130bba0c80bd5a9a95feff5ede076eaa6eeb89b59f7822c71ca34d598bd2426bce1df99164cc49b062969c580d9c70986b9c24ac4337dad9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1541b441eb49e0cc1d5aa8f96b462e0f627bd324b52d2f0be25e02fcdbc49f877fd581c80c7d1d362dc5706ee189976538475fd8960e3e0ffb2a93c1c2c6fc069c0500de0510170a174f0c49bacf52557a643152c281582770a2f27bd37ceb94f0e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b62a32e5565a949da7e4ef559fa5a4b56b9e547d47ae064bca8d30a29c69eee22d31cbceba388a49584491eb28e0cf7340ba387f68c62d92dc6cf88bf16796d3819bda6e80d5e509dd8286a8cb636b9142e2ddbeee30dcce579f46a0829a5fed88f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd495c34e901a0d2296968c9287efadcf77e45c95f956c2b601358b1d883efa6588d24609332c93e24e54611e7e5fbea3520defb68dbe723e138e5b6cdf7e746f9f00e06a458d56559d968811b7b96edb4e9a215a95629af1b831e27c1da490fa42ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e82ce60acd5c8e6445e73ee0fa6757e7fee20fb0251b9105c9b2b6310ade12def0185db6c2f563f9b1d1551ca98268f58bbfea929cb2a3c83999966f3a20def6784cbd2755acb4e921869a6927fcb4ae5cc13426095e24508b1ef75dbc8d0a3c89d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93801c0c98df9b2c167edfcc4cf26a4c29952f7573dc1dc9ff3750deed000371c4549b86219399cd68e39dc200c63c102658333e7a7463d873dafa7d929f65981c25a77ab07dae9b6f52a38bcd1a94599b666c305af71fbfabc156578a8a5ada3da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2891cec9462556e7baeb69364c8ed825fceef92fbedd75cefd8fdcb7a3163610a6cf624119abf414f257a8617b2767d932d1311c186dce8b63b9969735e23d33b9c03e6c3d9075180af7fdd283098ea48881f49f33640ebd14144b347aa4a588d72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a1059140b9314f9b19dd755179eec87093e1a798cdea1e53fb12606668e0b5c39fd83ddd406ad778021b5c46f36da9b3a336e09d8bb52a71dd1e0ccb2d07787b8fd809255528f42a347d39ff09fd18f7b679beac0767c704950c475efeccd852b17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h879b588c803760c9bcf7583f66739a24d25b1545f1f77a24a04059c41262d2619652fda54feec17e20713669f7b69003bc4b15d6fcda2916b84c48cbb850981cbdbc2246c2860759e9a20bae5557fc36187de99d833a9f2514759dda8cba21fcebd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1d089a0e01d78ec5469a74d285416c54bba746d84133286261b98873d8a97180a21917854b66c73da2fdac6bc8e58812210a1ce839d0f41ef92a87743ff3f1478b588fedc4ae3482f0af9e0ed91c83799aa0bf0411dcf44dd8f3b17d11dac72ccb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3db323b9fd8706e460f50df29632760e76c062ad8a6a9dd984c6202eac626de36a55290663801fc2e2aeff860e2335691d72117e711d5eacaea6d89d97d8534c1640f4b253ae6685737301d7e8ad82c62ba222d115338f875a5e6bb7a0dbd30de3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a67747daf5e7d28c97144f674a778ca7e690cda05855800d46fc5591911170f98e02ed339fdd1364a55325a90623ec8cb99dedcc07e226a1ce15ef1f4c8d221fce993ca5eb209f5a8661a493ba3db1b98fed9394c420491c5e03db3e4b6db8e3df3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ff6f40992d2fe3af46e11d37c8166234ed5a2a1236fe87516f99eba905a7358720304b2e39c954915e8e62e59487bd342b2fe349e0108b92232fc2d50f848dd9d9d2facaeb9ea10b358aba13dcc2325af5f4e611dff1a1f2379bb278ee86bb4417e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2d847edd1f6bf558f6196072972e6065a9bf0905395ecbb6adddde42505113a960de56a075cc60240888bba7b2f6d6c89ef471411a8ca4c37b51d4a6ff6b333c9880e1597722650c016d72bf2176593c3b28174abb25a2c782c2e1b0fc07fb66989;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h206833cf78b0b3e132d9385e44232f99527c1eb271124d53e618d7ccefb72c9e4868a9a6e7e75db9b06c3aacaffe5926890253fc8b9e8c2ee3ce939c06dabe764b72215d537edf002d926bb233307cead145f261395faa52d0f89410ae4544e9df6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2f371af23b672039f90cf40ecc802c04a310fede373f39fe779ddc1c6b4b29ce4b100cd4f2cf36a33b11a5546e9887aecacf061c438b36f0ef1044907c44dec90208026bc80f3c7a59a8d45af3e862363838dff3f6d41a0c5dad8958b6eaaeacb65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd6ed8db89b1b1211a8a973bb45483e5fbaec53d2d6fc948a1cbcee16507bbfc3e378dfc28e021c8edde8ddf612cf4910439c9be21ec640a7caa1bcec9f922a1b8d606acddd7b01c426ce5810c70f32ccd4b6885bdffad390a3f2b9f6ac95027389f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd340691ebed2f2fa5cb1da4431980d5c4e70abbc984ff0b1945a3525b3086c34db115f6b045f547f42f7fb95cf06133c7d0f8846197871f47d9f64021d60e7e0796180fcb2752faacde3e5c3b492a30418e988b9312ad394dad8dff6b1f646c38b58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h651eb7ac14479be258da972e2b8b29abd2a5e7fde24c127ff371be8cb184bafe9124fd77a0755495fc74853f2c9502cbca6695ef2864d56eeb748bbb38fa73ff80460f1f5a98cf8677d29793576fa2dc5b2a0290caa9c0246a4779e2d1b3da790b27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec859e2e4c6b1323d78532a65d4d3902e87050ff7dd27fea0a0cc9054b149e9fc2eec4cb370d37a0463e9b89866d1e390163e8f6996dd500fe739ba28adef202856ae29a7eed8a72da4c7c535faa77928d06ec17ba8935e8eaaa490aa17f40322596;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dd13bf8f4a21026e633188b3a4f90c94e5a0b4d9076232bf849200df8d4b4f62b2de7ec50756b1f82f443207a19a5aea8c0c5ea12e071f4c1c910ae3f1f7c7f7d5f7797ad3fd769b5b461cb5d6d5dd3af550abdadbcfd4102c15c4c5a6d55509000;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd859ffe0035b2618529e61ee558d0c733034cc333fb6266aa35e058fd3cedaac5edc662cb0a8721833b3003c8ef95ea906ab63107f36a22023d685434b9d9e6f2fbfd7c5cb1e54faf14671fc017d0d3af9ba3de9f5e0daeccddad9a602b63397798c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h920b8129f5221acd7f87f5771c917540a4f3d5ac4b2bb84bf044510a8ad0f5924146d9faa644c71cac80fcfa1e74950838990053af57a15ea6b9335c628aa85064bf77b316372dd2ee09b459761153e589f54f876ca5fd2bdd4cbcdc2275be3e8c2f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdedac2387d573ca13108fb49f719ce1a9c288adf3d13e83593978975e4f8eab596a1d55592f1edd017a1262b019212e0ede4f7a1296b659d0fbdbe4be54d95e8ee86d9e7e62ab6628a3e3a257ab6a86754e6288d72142608a0a17cc3601e576d4533;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9d1d2e1b0458dfae0ed9d480dba466f86e3b9b49367edf627ed4e5cd34df8760e01dd8f3e58776ef4ce27493ea9becefb8ab0e2c3d203b34a7bdacec9482ebea06437b6145285d94854139dd0014a33680aca82aa717dbf349a4e86dc04da8ed957;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a21e613647c976ba8806195ca55b9a32f3f1fd143d6b78b1b9c3025c1524399c550d37d49e78a3c84121f432b495aba72fbc630aa2f17cb7cac35fe2d9f682f14fc72360aa612ca0ae459488c3c908a93b22312837104356f4c9ddaebfb7e4d5b96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b7b890b4a8f331b395e57df535b5d235d816f19a34c4987a28436c1fc08ec962711539fad7a78069be6f62841099d210c5d504b6941e62e03ed334533eda65cde1c82aae3a6b81fdaeb0bbd8e0963fec5b1b6a925730f9337af125809b8ae3b14b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb51747318ceb8d0c593ee167797b5dea6ed495d95ec299532cdd21640cfeff32dc97b9f38588b21991b913895bd2dc96fc1a2a8780297c095f7693df4ad18ccd81372dc1ef51e886e418d176135de48e1a426853f017cb3f7bed539b20296182cb6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34ead37955250e29e9c56a3e414aac2e98fd77b3fb3bd7c3c5460e83aedc50343adfc3aa9591e91cead05d8e9bc66c3bc86cce5e7b00814bb0354334f2f6e92278c2171129418e08a17fce14237dbeb320d13a9ce894d20b240bdeb66a3964370fcc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h666052c58081d948bd8a821bcf06ff3b9eec2bf3988074e49b1767ce04773ba697fc6e808843790e505821c868eaf2b1d53eabd7b5f84fe8a8918d8450d0f78d817e33349a1b3dad23601428813f7179be18b1fc4a6933b123c154df35866a87db45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24b9c52e7824d8376737eb0f1a2d0199c4c6ed4999de69175a319ca2cfd80757c570439c1070bd914da42dae8a2c1b7dc69d14718b49a04306cfe8d846b1e60bba0db557a426ea55249994ab49015b8c48cbc63dac7c0c26ef6060deee788cdda214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b7107d8eb0c627fd22eee4ef3b62bacb2f449653fda1d7e01c15b29f797ff09d389378b72aa49f4dc3e931e676833a59696a9653f6bac713eaa500f7e25fa8c77d505a881059f32896151ba06d0e670b376d8dd9e140c6fb6066fed56dd750e8f6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3063be1c5567238d4d157aaaa5ae6a5a913985ee04f957caf9a888cfe7412e841ac3990653262edc8bc641c57b8ce9696ac272b6f8f1be21a0b5fa918f38ca76bb60e71fb44f2f97d672502ac2ada34467f80edab2dab0ab2373a30ccad0bf7380;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha25bbc798c0ce452d3c93e63b0db8bf5c6aa823a4295bcad44d246e0764a9f690eb63cf4296c3c4fd169fd2a241fcdac724169095b5abbb14bf2b8eccd0154e532eeb70edac527cfe32a57706311c0bf2302b468946af6ddd678b5b2224af31dadbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h342924bf39edd4d42dc0d84603881d21c33fa43080ad6478be5cf7c39d887242e2c6ccf46cfeb057c7c8ae640e467e27a7c864883fd69cc2ba031a841af66b805c4fd7d2416e3b1d613654ebafc5065914e82d1f6960ad43480b54550cd8efd251e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha02728e84ca551d759d0e0220a914e0c75028f762300cdb5871e74b654403c2e5cb465357fcbf7f725bfc6d2454c2cad40ea74fd33c2fb8d9449082ad5dfa61544b7ed172563b9c40e8cff5a2dfb8a12ada0816464cc18f9ab10d2ece82add6d33fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfde87c215cc044d1d4e3409abc4cc449e5fce4ab07509d32f0adf30d1e9ddff4061b71aeccda779d6960a9a85bca69af3257760cf9921f1801dde1a3a7c6633aeb7e1ba86b4940f197bac9f7be87cdaba8de96f12cb7374755267c05955803c4ed57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf35b28e17c909e22b3a40fd423d539c8ce9b8d1edf6d486c82238476690ec808eb1ad167e23979c22172ef34271a7986047bc45b0d64b427a962bfe30e8a65c48501f6a6d3ddc37482fae72b4cbd930cc8a7536ee87b7d20bf46f7e873eb3cfc44f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb028dd71254444cca014bda72ae9d381bf9d8c7dfb90e7d0278d813981a646b5e05e9d151d63b94837ab69751f80c043681b991e541b96b08d239d0060b8e02be2c129d6ae42c9e25050429c07acaf59a3fc6191de002bc00b1e4ada31e02dc4e462;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80b0d966f2784405d6e4805fb3fdaf0f5b2c5ef8fe0f3748e7877c42eebc583f8fcba1e4ac47b15cc042ea2a0eef55213fe54e66b8f3c6309b60480ae344f0be58219409abd1c58ad72f167157c1fe5c4d701a804b032e6dea58b32daf0d5d1b7538;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8eebabbcb1a3b80360eef210261d8ca46a61385e467a57b8bd35c31972142dbdd2f1bab2ce5d6c95d9a4c43c6d90c56c4340cf94eb02ef8d7bd1acf391ee398e9e8bc3bb5b785fc7ad7ed503d8a40f8e12ed54508f5eea3c5f76b2dc98c84ddb9dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h371b60c7f8e05a0083e5efa2cb3a65f7b0a71ea4308de179810cb9a625e39ef6089c5ab17bb253392e4f5b00ad95379cb3df25de5415e0b2e884486feff19b48fb79d8574dd59233d6850b4907d0817206dfa6124ec4693f444fe1dc36ffdeffeb89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb812efcf88012af507f9cc07cc4873d588bad304b1faef64ea5a15893b695bb08068a8b2c2ca5c9d1820398c8e410596f01521d2eb0801152a083ef81c42f1bf3cc3d730f29223bdce11365fe7b35baed38340325d618857a7d73cfff6cd92af707d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aafc6d88237aa05837ea22348166fc562d1cd6de353d6a1957f1dbf070eb380352d0d1a4f361060d8e7d19332fba2202e4b16954cc077697155abc7d7d5b73178b06d6007f56e8a5bb46654498b96ad0efa3457b2927f01fcb4153301e20b80bfc9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b1180566c9392e18921d27d60110a14d9fbce632ac5271bc43b892ce2cee158f46cf929a639ef2a20a5f5f9e9dee716529923fccd25080f7caa88d4ff1e0054ba7652b4f1857bfe7c5f11bb78185614b35597de89d59c3bc086093a97f6fb829666;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he13f1ea2a3e69cb43104d5c1166bc2c8e5c9a94280853c40a6a6e8691c075d62ddf75f2831b551ffe75524ffed79301f8e0851e7647dab414133e8d9117af241d4d61def52482f8ebfcd4fd4c25eb2751f741d28fffec3de09a3e818238228d3b902;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a6270417ba1e04a4ee7a02a2b0183d1c5c3f73e9169e967ac9a72caa93372bd9b9955ada6c80b2d8dd4c286fbb0d571c69e052e1e405b8cd1d865ae69a52b3c083e2d2620a615c66a9386c6c4ad217ff7d92fc72a19340fecff04956846f74499e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h701b7a8bb3b7d23c56e52a3be4a6beb548348ad04b3a96ad278224e06310909378cbe80dd4d0f976f1ebdf6f40ccbb684e9c0e28e28df2239598400ca393b8557fb5837fa552fee35cecf708bac00c42d0f14291b7e8f9f3db2099fc0dcb888c419f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h971eb614460c1414b9c25b17372d150a6d47b8d744b27e5a07b0be4a5ac9c9cbcb52b415fe9ffd0a1c3fcb2ffbfd7ee5689b18f1790c204696d17feb8479a6a9f49638c677dc0f6a0feed71afc0ff9767b4ff7a4ce2cf148cadee5cfa8b91a201d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2225435f836ada103284259ff9b1238e05d2a60fd87d0f463735d663ba7dd1ac840078d1b65bf28aa7f04bb018f8b1d2eea04b06bd3b76a6433d96dd70505de2547331e717c1342095e184bdbdbfaaf80ae4366ac73363ba7193f7402b6236c98013;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76ca42b3a88f7c5514691898c525b0806f3f0e4a77add82c7d946bdcd7399a0729486107e33cf4fd21223fd5ac419f1a2a4b563ee7d638c822f9542f80ae69ef3506d3feff984ad98d304db06879d5daa938a204bae09e65c201af3f5ab30327dfb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2cdaf57b0bbc6e2891312a91b5deb3f8f1443b335555ad128316191cc4a8d1ffbb7d05bb85efecc05ad9479fbbb9907360916d1fbc70bb5f80c74318191cf03c8a72b0c1c8e4893462ca42e84d91f1c4e9b8a759ba4e0fcfe063d0396ea55f468198;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a49be7ad52def542707f8e14c23d9e808400b696af0b64cbdada19399999d61094e6a80d56173636ff8d7095443d6a8b3b8d2d034f7d447a931893289605e0cdf7def1c71493b779c5e475faafbbffb3a3bc09ef17f404083a68c12e10495906c1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30cf7c80beb6563ccd272b5f687d45f6668ff0167eb96ecf06a59b3b2d7d3c0f050471d2c3e01977394c9092ada7318d0df687b7bae85e708853060498809a5c91c2551f90a7023472efe7114c1e1b711f720e8f072351eb23a04d123af11890291b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26d55a8313a34c735384ad7fb7dc86a5517a7b3f51405e14853dfc7cf59113b730125c83671c81bd89a02d8b963af2e8884d8fba16a90cf169ad8cca93777f2beb4dfcf004baa8a6e8bf3cb4781fbc1b09b5dcd411cd3f0237c841759d8b30502d78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h183f0f2e1b31c59663483a716d0b35366b3cbce3d538a1c2b6ae9085943bd0129cd3ee6f812b91bdc9c55c5379d4e6e139a293765db31397d26a6ac27f69f00703e9f709d0f1ae103996151e88016d81af9245cea1095613815d559cbbb43c2ace5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84a0ec85323745105c95c0cca06f84c9e58d103f6a32050fd0c775b58c3b414afc7c891bf02fd38e5d218b3b49fe3624517cb7ce26ad08cd904259ca19d4daaabcd743f332de28f1514e3dad4793337b5a78aa415054b8cef06362beb306beca36c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d14395cb4df9c3870ef8c9352a638e7d2611d84e0a43c0ed2d3df3b8af4a956c90ac33d3b5e5f8b422c9f1abe31d3c4404ac7908104aa91688f6fd4e6facb3fb5fe733b6136e133f0683428208d7fa5e799c94d2b64409e2a771587e06be4caf80a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36ba038c061e7e8ef4703dd505354d15196cf0712f270f713778ef2b2274d87f6b582a9c16db023293f3982f481e590af6cefe7c0b83dff55146147e4c7295665b95770d4688b74e3d91f3a3499003e380ee65dce2d12f82267391eb2b46c7fb4080;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf41d96b4d07573979ab7ebef3455258572ca376a7fc409e9a6ba85b01df0c6432c00b6c641126e38696493b6039d26b6a746ac61044b4245a724bec08866f65e684f06c15e4f75936913f597368d439930b61ffeded3546fabc4196f6b5209b7202b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba9d90383dc58bb3d7452ab44e411b0824353cef2a61accf5846ea57972f126a63b0a4418de9a81ff8e9e658a3d9a8241a374e271de7c652328864be544889cca315f50ca915b9c165ee31a6efd33a504afcf5f77413e82968723d4435c7cd337301;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb175f02c2980656bac914d764752c540c535a80bbd65d83822dd44a19ab72e5a22458778853dade13d3d8d5fa557d872ab256fa638ad6a45694af0d185c60d1b8ea3d5adf06d52a72c0914e44ac123e5034a086be411e4e41cf8c231881cc95e49a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73a9be699a114c17c09719163b96f2de63cdc4251bdeb174877b7e5d519004a4c6a46367accccdabfef6c517c2579e953198e860e7ae0a9b5c663f9181a1e3e26a0d4679d146d7b27e0e1dc0f7754a7a565a1ef60870426195462129ee25ff0a6c97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b547bb953ed35242ab21705d72276524d29f3353b4b2c718b6de78b6b64305e2b62ae842456512d0818cd8d1f689fdf356a8f307d823d2ce4861bb5755bb6f6b6fab55b8386910927bfb7d9f367aaebed0e646d9e3e4bed039c32ba002dfb05615;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab739ea357dde52019ad9899eceef9df3338195ae68b1c84184f1b77cf46a008a45df178b3c096645d1793b047af788d8c6256281a29395faa7df63a6a79f30c53bccde5479c1cb3a09b600def2b7e5f175657203b682e86d08518ab7d98a7824af4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94cc8f1cd0e7d3b0e1b42d0827b305e7a103e74db068aa398dfa49824afa4ab178c7cdb934d7950552214ceb673ad5ecdb3714c15fe4b24fdc36bf9eebeb642076cb38117016deef57e207e1a9b0ce61be1530abb8eef90b9dfd4dbe0d2dfedbdeee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1bd83c7c535afb68c516efa0adc96588a9170ab33e91b0966303e501fc856c700d48b0ed8d9f5cfb74ca99d285cc213f96b15c28484eeb5f976a3e8d8ee510ad2b2ec6475ce7a569bdaf081428d24fe9cfee27b559d520e5aa235800551b0151be8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3077f32746b9c6d4f6c5be982c8f80fdd8210b695ba5b4076d72bc3c74c14d582ed14472d9713b66bc397e790ee655b48620c85d7370d1fb2744c08b2b1f47cc01f759b81823dd68314858d90e3dec9d465d19b280ebd7d919a4f5fc15885404127b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65d701672f288e63dc7c99d823973784d646eb442634f7b7dc07e306ccabd0ce6d20ab9c5d999c0264a24e3edc82cc64d17ca40f96b8d45737285a6db49757915bcb6fd873c05ee7ee3dd2abd01f005af5c85f2f139552737b8ea12fff427c148ed5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43e44ba36e20d81067cfb924970f22e47ad290505dccbf399f945c7aeda7f7ace52d48cdbabe14b57f83d5f74bb817db6b063a8298857a8320a7d0792f3bd5f5bfa37ba30545c7d05b8d7049328f2a4fa4a5174dd9fbe0d0eadc1d2536cd6c2eb552;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf95cc62f02d423f958e6f50ffcbe18f4c236fce9fb337b10b3b7150fbbdc876862762dea88dd0f9ab9e798bc7de3e5fde9158189b69742dbcf4ca60f66ccd1d686778c7a2861bf3b5278f4fbb67f8f5d55d0caa87dabb1a1e26bba2fe42235b4e7ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5e1a1bba6cb224c73120c34ac4facf747721ada35fca5ee63effb1b72f4e570990fb87cbb7159de7e6feae0ae6878a5b191d1fd09e242e18e2f8b8b764a68a1040f30704d55821f02226b6e0dece61816f92bf35b8e1c90daf481345c1fa18d70a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28628a2878b37fe86d01f46d2c4c5520886f7972b02733b7d6e2ee06b7f51da775eb5212fe59ffe2171e0acfc5039ee102859b8c91b5b95b4bfe11478a18e9274631a94954fa2e3078ee519bdb80ab518aecf872e90835626a2d34daed8462a3d15c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10e01e4e41a7f88355e229513956e15dc48de3e164494ea8bc2eb655ee1066812b41007cefee3d61401418509baf3423bd310ddad8e3465ed0a4aaee391140305005b377dc626273eb8d1f6b63a0503e65c97f7b49022e0dfb3fd658f3ea6c796440;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf42a926e8fd8d77ce9eb16ff710c65075dd7f72272fa29999a4703ab09d27fca6ee0b6116a343c51ecc6273a60797c888df3ce23bde7298465c50df6e76893b8a9cfe13bb68fd197b6c9193866b8985950db0920768c60ab5caef0ee88253610da99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda908f7194801552dfdba598d549e9e28cc2576b6354d400a53c3f8db484c64d868b3c4ee4628734484e501fdc14b925d4343103bdf7fe716316b4d7fff31273473df92e768f63dfb1ea8e023ec00f4d873b83412f84928d637f31e3c3a0f3b258d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7768f5a5616870b0742ca2f1ed05929fdff836fa7fa64c52982d166c528a550a972a349f62b60220ac0b5cf17e68245a94cc69d535a8649afaaa3087f8440607fe2f008f7f5c40e70d40a44595557ce068265251415cfc58f72ff1aee7e29f982e8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5437e682e0c45c6e529239907fe7a1bcebf519f880bffeccbffb0b985264dbdd881986492a9008be0dfe2bb8e2be3ff2fc40594af48136abc8f9346dc58eef29153894b8409765d2e16e759b50394fcc1ffc97266ecd85f0f90e8631cb16b9047009;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h821500a5e681eb0eac3b42bcf43a02698bff816b74238247cb078a9f1e3f068afb11fbbc53d61a0701d203bfac8fadcb08baa700680d246531e19e25986190c1487f240a55a3447e66eeb870e8fdb86e642ac63e362ba4f300cbfec4418cc72cc046;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0d332d24e159221f9f6cbeff22befb47f9e96aca2acbe682d279a61bbfe403fb8516a77184cb3c0def314fe7828b4d2600989b75f25fd5208a44ec5edd01aa7d90a5f08034b48258539ffe0017d8d8d92d47a45e6c4779fcccb32fe515c348fd669;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f937e06a25a04d24ebdd5903cabfed1cdfcd56c660e0aa8213900e659aac9d06233265e3938d7e579f7e5436bb6992ccadcc55bca6b8f87652b0d80fa6240152a42f2710b8978912759300e380b295e278c531a8aa588e6c73a83d09383999742a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1902985f4c6401b0dd46639841417d0f83c57779737f2fad0fe00739772f071e6ce3f74985d1f369098858205cdd7d2c0ab0d01b5bd2e659eb793619aef81ed12ea0d61191a3ac7a46de21623655d5e5737c25bbc576c572f225a82408d2ac572bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55bb8b6d4fc7e2a648053d5df8546fb1f8dc6ae51b303962e92e00c06267fa90b0541de48c6f6b74123cb5caf8816ee4440e19fb14c9dbf83f80345b0d39a5502d26a1e063ff1adb0f470fe56ebb66f90ad0d12500a58bdc2440a1d22e04dd2b1ad7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hadff148731c41d7c350bc9d76cf13bf2ae606bc4e8d69a11764db3ffda3d2bc41db6eace45dca6a394d9482d94e47b95a36519c189f555bee749d8616242a9b547351a025e7e378c5cf9aeaaa35a7af9b822ea9dbe28ab04f5c08b51f8dc8829d682;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfb25d8ca8548eda0fec6481657427cbce2e4a1683ab1d48b0a808b9a2e72f8fcf22805228c817b2c9e13b9f58178bf1e3aae4abc556319df2d12e7a379d0cee9852c86f6dcb060a653803b4d86e6e0a57660008261587e66699b5de8f6d8b1de7b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9afc522e300bf7cdb0487b001105b5a55ad375860a7cc9c6519b55e058eacba2e61d075e9d00ffeeda81437eb939446f6e4ca2fe7df89d16e60f227b67644acf8d5d664166707f568cd5f54dfe7aa04d93837af8a6a2fbe7a10bd4d12310247a3e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c54fabff43e3958d68acfab03a0a7c00df74d3df4667612191c89a7478f897f5bd0dfd78759c7dc303ba621aa5af22113d0dde777ec8854fc275556e4b00fe695cd8dd41473c1fd4a1bcb943f2967cf9a0fa93ba703f0781b8798df53a4db6706da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h632fd3939024c8e424eccbe2fbb156b69638ac21312281948962cd11be3dddb4d6dc51757d0082620d0caed47f39e3b7a46c5d555efc353f3795fd210248f995a89c584e701f54e6125b17c50f7abf5a54cb61e5ac173c4f164d1d4873d68ca481d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h554f774d3fca16952a292ab675756bf5376a6d87fc9454fd9cb73719d11350e18802abac5ed0158e95dd5a74459e60285b9d0f09bef7485b245197a046cefeca58271db4dae1bd2affda7794ad126739e8e0e88c6bebe0fca2264e9fdf464a716239;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6a095eefe5bb1029335e737e985a6f4119014d8b5f35d08231f75729a5dde6c4ecabb7d8eee5a0cb1d684e8dee921e3cc1056363739712cf5e5e0ff3c72c54e28c13413aeae8815bf6377c950838267a9cdbdc800b79885ce9539fbdb2bd18bc075;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72689f17c0601cd70230d7079672816ae8e4923dcd701be162fef62ba914eabc595117de326e2e24de724beb9f8df95f0d883575ecb377977527b4a5fadd85edca5f443e07bb6f6a156d69af1708d14f5d074e123df3155721ca869b177182f1d8b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26be0efe7bf1701d05a0f3af78c8f8556b29cb2f98b70a8ca779dcff828f7729906870c936dc56c41ba25fe66089bc90d3979e3e1015f22d833178e8d470565789be9916901e0987f37af65eb56c77f19f102e73959cac7868b21c7215209b5fb086;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had79a4ffe2cf78868b3f08f4542892244799abeb10cba4e61ff69ac1e5d609f4200aa8945b59b4339749911a3257fb3e884df5d106c8ab473effca0718f0462261f4c73697915b959b42ba4cfc6af7ac0142fe63df872e9b8cbcf9aa44bd8903a234;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41df36eae347f9748a56f496dc9e67c09782122c66753aef313cc122c8365728becf14c3891c85d25c7497b75486cf716e9f81bf84f94ba1edd2fcbae1c0cd471274bb0d8a2575671b42d55b04a286fb746c49f4dcaf681715fd8554c16f53738712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed3090b4fb689320afe11b21dc6423836e04cf36387dca18904dc9e7e4b915aa6eece673e85041ca1110e3a29dcb87de1e86ddda38d752c5e0c43bd35709e0534bf6307d5183e272b3d722c913947eeb0a2cf50031d55c4d355f4611b451eb7967c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc087d33bddceab8804060dd769b87ccda256bafce12a3cd819862b5d6d9dac1446dac3dc766153e45d459d465581c378fae4c8fa3f7dc23d656b29dd9a415a4c68b736546b12cc146db489fc1df7b8cd66a1ca507c3b369003e4d45fad54b646f971;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf285899dbfe8c50851be4423728f5909d8f0b1f87a8cbd07e8c706c62e0df48c948a5b9620f5e29e7386e32e15a5b9f84a460a1d7f4b8f42aa0cee49380b2e8c60c1a1773c21427688b3e365e4d8b6b2cf6f6a8449abc69062f1a1a9ed4359b7bc21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58b5615086348e296abff7d344324d7c4fa7d0e909c0ef662096e0c601f0a9a183f094b2b32a36eed8a41a4eef40d4a9391490674dc8eff97f0a2bc4ffbf74bcf525c09936a2e9551232349af8c986a42656996dcffa798168e33dc79def5d133ff6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5930024b7ce42e967aeede611562f77547fe8005f44962b928cef025705a7394610d1c8e74d0e50339fafdf74385da8fae9df7a4a138dcf5a85ec0213831f4db8454068bebcb0d99d207e91da73b3d5183e92afa3e9cb7b2a4a77cebd9487ea4f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7726effc5c660f15daba6ec69bed7eeb1c3243e95e13bbf4d46d2ab488f3aad89c1fadfa1fdafd69d2441106fae5c211f095f6e6ad1cf81f1ca553ab1d045d94c878d0487c310ef43b44fc6e3f92d46645285d4b37f3742ce44a32a1e613a188471d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h896b080fbcbe285937af375c76828dfdf4a3504e6437542c8e7547393aa96d1ba343a4c5b287b336e6a44895165708e17d64d8b18744010dccf1aa0394f8463e3afcd16b9dfeb6fcfce0dc6cdeb5c0202a599540b8c46956486f2577db3fe6846b5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe2dfa25a96a7282423060a33274905d3cdb6b68d166925bd3ab4a42e8f06f7cc34ab9f44a842362f71747c6ec9813edec0142cb66c099dcb3bf4484b3456586a1965f822e30d5f6995ec6e49764e70f1f34a3f1e00cf88cb67656a8832b93635bae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h667fc595b72779f19f03be36fb32819c926b40e1fa9190785ee09267ef820cf534eb451000ec11241df9ee03bf2cc4225286463de8f2bd1fedb40a7ec1329f0760004358d3d408f4ee6b9187743da753f57bc11dfcb068ecf9ea62bccd45cef8ea1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h964f58f61e82d8568c6b02b8eff481a5a1a3a605663ade8df8ca9152821ca76e1222a41572ab59a31e33274ced9b023f012c31566381d0a0f72f5686f08acca19bf9712efd8645ee3be15adb1773eb1613c06f73804497d4e7c1a2ca83468c7fea8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2c0f9771e0be9d1d18a96cccf2be6a18d9f1254712efc77a1b77bd6033e6d020dac84c6c7c580a669a33599e37354e803d9feb6548be47f353ead1593d46ee3ab57439e659268ed071808ff1c8751bf39462aa95ad405c9153f580d52367aa32643;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4282e9e6380838094917e4d58ea7f1d93438580d42e622f94feb42d01c5762cf0a37209abce92f0c593dffd77a4eaa770e486d73cb5e0f839156d8190c73905ba2681fe58d2c2acc06f9d315e17c5791ff59bb4fe1bd577c670b6f7b16e9cdfa222;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf59ae8fa6c8d2882cdf7ed839a4d70426740a4a4a9b5ce05efe2a94015a4ab6fee992bee883f48b6aa02bfad2a7591076373f9728b5eb7504e5adbce0d24040915bf7dc2db85df18629e343f713230679bb76a8a560a90c6157dadfc19929769afc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaed6e927fee6e73d233c11bfb02956939c678fc8b712c68dae18f2942b964583a06de4e12a2a60bc553be9804f730dec72eef1f5baec3ef208f2cae5ab9f92ae6e10152886b13d6d4f054850d08833085c1e6038c9df1ff82ef92eb6a2ae05be973;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc59ab1e8875d40cf9c2452dcd1c9d53a186b94a4fe99937525ae1ee7969f923d4d74312687ae11945672e673d1fb5bc281f1ec0eda9ff802287cfe75ac521923c7cebe50ed98a5b03bac2cfa601cdcd030144a7fe5a133dc40ef9e40d1d46f697f07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77d7b23d43c19910a7fae21552fcf1e12afe1a53d13e32cbb646d867a5a0a953aa3a71d132bc65765dc76ee1f6d82639c8adc2fff7867acd03365374e8530745a401d86b413a01a4279e32cff582cc27e4af35aeb1c0d1501a188f6b1f2566271319;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40971b16331c4c7cc38abd3bac8b13b8cb09ac441fc2642df98097b1498e028cb8ea7f175c8f96491f4dd5aca8a4cccd93da9cf26b259fe5880b550bd5d2354cd2d0e71000ffebbd65dfdf0400f8bdc6bbbd697c6ba9620be5c585317c5f78b2614f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98c607f5c69522efe0f4a92bda43d195b04bacdf27eddee118af2999c13d72d83ee4fb6fc21537c974f62901aace13d74b4874a300b54724a2e65dbae3dd5052122f5a654f7d8f2a0efaf15b14425a7bfd37bf09926c75ed5632b7ee50389afa31a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h363097b1808f3712d2f2b50f6d72a46ac1a3ac5f297f28264b0a9ecd538fbdd6831561b9d71eb27228458c371300fab60d35cd273dc13e65b24e2f84a1d922ecf998642c196683918083dda92ec9b07dc54aa55be366ea200a40d910087f7c52360b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4523abe95d90f76fb501de29b3ba6224f2d4d6c32b2d57f1343cb50b4ad2b75d6b80e305821d0c48743d33ea7404856c8dbe5e4000245bbdf4b2e0831355956b2205265d4d895d7d5e73f2f31ce3325ac27a5389d08b990bfaa5e06d61f9ab780d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb41fe8a7cd3e46bacfe1d11915218c877c680e8cc3f1e495e1f42d1eccae9228c96ca93fbc4283e2cbb04b67e66c92e2eb6d103a2827cffd1bda37d85bff4dd0e9f4e2ad9c4e22ba688be8587cfe25fc5ecc731b99299054d7a2379f85eb8014dae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5763e65a3dc2c4b9f7b75804063e54135060937e4795b0b27077287535d7224f3776de12a607330b4834c3a67c7e3eee644ba1ee197dc411dbd01ae92e898e7f54e57722f546a9fcf5c73a8b6313d79c0e0b05657f31954829647f89dbcbed5fc22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76eefd212af82dccae2b03fdd136a9abd616830b33613531f92a5bdb2492d4bee4405c7d7316ddb1ea9f6408a21704c9dc3db183b847d78341cd76159c1612ca596cd290d0d852460e649c18197eac25786ac946b1443f20c14012571e0dc7bb6135;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ac6d2fa4c86da43d89efd4ac0d3529bae78b300dec314a209c2480009ee4b60c21bdaa545fc329c20b70d3fa88f825c249859e10ebe216abe0c15bdcec8affba1fd1cc627cd2cf37c53205dbef59e07ea1998b366de64bb2a8bb2a03e3367f905ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4abd0226986f73842a1a48563cdc069be7ffd3e3659c0ad2d3bb312d87944b2cd8cab2398b13332c83c10a6d8d29ac5a620444012af18a48ebb42100d0d8ce6f640972d65a9a727b0fb32c74006916bac61df6ff1439ae94f790b2b202f7c5645c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd27bba4d455b521474459bd4ee331f1a2445fefc4477a5d817489b3f276a9241ac27336537ee4606589b90a38387dcc4553731b1f1e030a06d60a3abfeba9063a8aa86883e58c7423d7cfb1defe16efbc21f667af5895ce010407eaf803ca87ee804;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d56a1626fbc2d9499167e554de57f1277379f6e1965b18dde2773a3048545b2b7f2d20cc6be4651bf0237702141d8cde6b906b921eb3686e7b9b26d217d889f2f39f1db69cfbf07e2dfa48e989a0fc8d523ef027c619f5e20441987c7eeda90a361;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dde91e37da3b1a0a0fade41101c7e7d4ff171678047e3369ef57c224dc115ff594608e940d6f1a97a9460d60117cf39163525aa7af9105ac2050f6db837a6248287ea1d991f1d512a6275de996ab5e0d2fc47d566b451b1c8deee9a9fdae51558a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6f1b52da660b5ad567f4011412b52d1721fa0f58e5a6e642abe73453d550815c9731341d74fbc047cfd8a89bf38b3b3e87b78f71587930a19cf0ba59676c6d4c4fc7ee4549c2908d7922c30cf2511c50dd3a4b330190902fa2333ecb9e6dbe181bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3af068ba69ce344bac12ed21032af627caffda37af9b8eaa53f8b1dedfafcc98702d0cd87a88085672c5ea35db056ab0af671b90b3bfd44af40de010be437bdf4fc4024a1bca54ddbd2394d699e8bc60e97678248fba0eb3868c00192fe888f39009;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8ec446e33b34341ced39e33a295842473556939a93bce4cdea78df4c0b581725d4e4849384f2fe65917021ebf53a64a259206389312e2e1f4544ecffcecfc556f16e080bbc08d056b1c86bb888e1b0887f0983e5f229087a0abbbf33bc2dfb78775;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bb758501e843e769cc99b5dda1f3e4d73c1e700584a2afecf539fa5152c26499a4e0c70d8e2fe53611e90de6b236b3569b5863bf5579127c402e8d9a74fb944919b2c5d28121d7c893d558b4b5b67473c9228351b7b707ef4020eae6d6940845896;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h408f0a813402730a0c80407509ab54fdc50010592a4ac209cce7c3766e8123afeb0fd5f5da6b26385bcfaecd5e747da765b5457196c615deb19c2745e75e1625e1a1de382574b3e1ec85c2d7ac597664be2c5930e844fe92ba7d9786942198d2f2f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b3262e3cb8f38542df5d6c6a0473231ee4e3034406476e8e0bb24241b87b2e59cf6cf7afb3f199a06cfdcc1aecea81b707b929e88f21e4ca8d41c437aafe1d7a3bae076783ddcd0b0b05cce6138aa8ec2fa037163b40e24b0f498505c17bda1111a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a529e3b9d01d16b1fcff3934dc338431ed5349bbf491724c7147cb35c7fb4f8612b28e08cbe235ab2355b49e7193f655ad65f4110bea0e8723a5a86aa62703cf2c9deea96abd03f2edc170767caabfb38fc4451dec5006bec3ddc3beaa42d85a33c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd888e9d94d9653ea84b6f4b7e7a4571f689ce7b53aa3ab1b1371e01f5b6b99450b2f87dd6e9dc63c4d9aab92ba20fc3b1c5986e00b52ab8efd5b2b01b9b75fc0b6f2f11c493a938e2842d6a60a8ab59764a6d569d2a97b6af38fcb6658bfad537ca4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6eb038bb7bc3654a0c28ba415a3e2520559dcddf0d5aa34736c5692a12caebcf80905b8fd6527e3cc6d5cecd353e073692a4b6d2d0356a03366d61ea7eab09836658cd0d85956d7baeadaef6e6606879e981394dab0f7bb5604c639faffef0c69917;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he655b3bd6f956cc58b2733cf6419ec218bacde0b6db390aae92fe0302d4dbe05f89c7875fc0ecd6a626944f55b35072c4064f0524bc93f3d389a997865f91631934fc66bc310dc66b6c7e8e850bd221aa30796b8121a47bab9d2e9ecc318dfa65461;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1817eb5f393dcf80a84a06290a2068923fbb573950a4aaf51ef207e47e92a8b11e6b84097aa85b1b7e64a587d3efe9a771ef866f15731f76cd632a03c137b3cf0d8c6e8aa7c25c6a8955ee2ab9dea248f747b57347b34effe0b2d5908bdc60024e19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31daea5309e832811af0d2d388ebf09ca362182030d3fe6802eedaab16c210de8bc964ed666d364ca7ab91f70e4f782028fbdf75c4c5fbc2ef6134ffbc8265c8207953e0ec4ed28dca5fcb49f8f88ec1eb39856781beea3548a694d5b67954f6e384;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb2b7b58d138227c6f60e96170052c0ba9e6b14c79fb5ffb25952f1bf14a6ed094b8174a91b22e0647811af15a39bd61bfa0e1598a81191645b0c36ac71dabbb291af12027fcb9eea0375deec4309373cee2161853c006fe797620c40238b1d1cd5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf3af25807555c57231e0e654b9ba4aa3a4f8b83f18019dd8225351d67b2eb6c3562b40f31aa5d106d3887c8eecfe4904daff83493ba5fdd92c493e67f0573889579c3fd30e0f08d3ea6561e8e1960982c0d94bd761e9dda80ca37bc558416825e9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ca4a5fae0d6da1a7ce032156e8292d98f5ac95d5bf57dcbe4627cfec51127274e4703c42a1e743630edfa84a1cf7a2330f61f23d5465ee622726effbca608a70e1e7e0514f35e4659c80017c8cf573306d9cf0ea9447d304dc1075df70f4eae9ad1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16e31d0ccfbe6ba7fabd2ab72cac9f4bcc2b370729ecadcf1613d38a250f0996c5507d2c4c0e60d738892a48e9f562651117ba134df059e09df12db88fe8951ce257954eeb2f56c475d25531939cd56633cb5ea95d91b236787a19eab00d1dd6b7f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha85a600711a2615bbed6bfa6c0c75b2425a287bca7cd36b700f4320419b9078cec9e7ef9af9e5ec5b55f273e140575a6d3893338e88c31f67d8a76453320a0c00e2be24b38f9ae5d5e55a70bf53efa74735e204b08a662375f6a9739b6eb37b63e52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7d42352e635c7a226f4b1e82afd897dde86b6c4d1cdfd620b9ba428d08395b66ac30865fee98b0b2cf3a7ace659242e5261f7b32549a0faff1afdce0eeaaca91b43846198d421075a4ea197f2c6ae2c6b4c9691f9f35c16f04871eede9e8aec6c95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2898c337c076101901d79497826f280515e5aebf3fe02852b8a8ec959c8131e9ad5f97c92504d7a3914f1cefc72c6b84db0ad3a51bcc9a681548dc276d6f2058522d1e8b1293108b3ed4dfa6ef88a3fcce2d0a66a1b29af6cd0e6e02b999ff3075db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h886cfc9c3f26c7213f3458a10b422c46b7a383fa53cd238826dcbf75c6876953413c40c9d6cdfb2b4f128bc37557453d63b0595ddbcfba2bd42b093e598a1e233aa4b8e7424f26315c722cb1b80f392ea332269eb7a5c11529b4cfc353b2fffe6ce1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49ba3fb1fedd19d604ac2e58d6ce3a5516a024ecf5838632b1b66fe8b28aa3fca3a4b66f5cc08af355989e7581bc3d8f183b74b0456d8524221a54c9793a322ff17e1f78fc5c7a5cf57a50d1cd76fe6fc0c2e252dac9b3eda6d3da01b63819cd260f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd27a8fb42ddd6fb87ebf87b83467f38b8df10d17dd57f1c663e78d866e90f6c5690fe396066c893af4231106adf5fe1594e2708fb40eb4220f9f524f7a1dbf8b6c6f6e87f00a55e65ae863be3e8e7ea60676ef630ba4ccfe88722c47799e924bab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf08b78ef75e029c918fb1bd2276e42ad76a48713d0b17554d1bdfdb52185bcca4df183ad6b4199681e0d9b5b6581a08fba54aa144f66bee30dcbdcd8bfe87852d24be153d86611ef49aa3c1da9dcf62a9106e72b503e2eb8cb926de9292c0b3baa37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h278e899d02cd4644cc9b536edc634de2ccacb6568ca030d7eec77f8a8aceda0a8a0693977c23bca80248982e9ee0dce23f4228b8cef5a25458453afb847f57e4a00b71248a6ac6829f6d9c7f9712b5778bf88e9ac9beb3371a1126b48cf9c3db3d62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10e9987e36338d8c01b12003a2096def2c7f6a7abf788d1645d893f51d5ca181a38002df5f331e1940667fa2c64671b3b14555a0b63741d57d0dce07d137b6b0183bbc30ab74225612010c65c620a85f73aea07a0c1cd56cb895e8888a4b7c94c8e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ccc1c7921777cae8f10c97a850d76f3632e4986a5bad7c710dd0a3e4573373e14416b7b769236ab3df1c86d8fe63acdf5df1306bac87010d7bd342541802f04e0747abdf5e7a31c65fcd405e9078e31a87ef2031c5d19cfb3c22d0e8700c218e9b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebf2f0135ec34d6fd14e99e87836ee929e6017dd620b170019dd43dce4d983f639ba30db42d57fbf204510f91bce5ee76f2443c667106d4a607a0fba7ee63bd8d41ffe4fa532c532d8c275fc55f739e1d4eb5fed67145d5f7d6c7b4cf9b4da3710d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0a8969f7b8de5123b13244645a8febb89af9643d4b94e43247664778212efbc7f6419967f6425b0d3d3cc645e75ca2f6cef3f8939a7e8d82f041663170030593b7e15543e97d05753ecec08bc9e362ec77c1871b82f89317a649c71edc6adae9efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2421f4c4c6163e8124856af333a759c6dde51cc0126aefd3e0b071b8caf705995122b695744ae5a21cc2a9f7e3ff4d504cfa8c95d9989d8b7d273d650d3dde5fca6b322b04f98d0aae1211ccc56f0f913e52b36955a9faaa2b471f74002e8d38c6e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63ccf4b7f177213245ddc9503f1692b123741ddef452a7393cf6381a38dfdcc5dce30e4aeacfd713e62d11b84d1eda8afb2c0bb6805fbd3aaab29cb85db7ca7099d5226d0e1c4ecd929e0f8293c65b1528e82ca7ac5cea9c10fa7e5d4dd05e88227f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92c3c07b7636f0e7030a3a4ea5f8da5635f43ab8ba5613fe9e64dda7e581e3aae67158d50e20c24d8814803d97d405bf429bc8ceded7e58d666aa91b767d7c655ec8f59a348ec4995dcaef5c7899f010974bd0463a3d441fbbc1c25aebfbcfdf4c3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdedef240638a8a2b077fd799f6158b16b6a80298b2245c5d7105d782c685edce6c216714a74b085e2256ce64a2d99726eee81925fc19e8f55482cb1e5f6b4d525efe163bfd7d2d5a19f4b688e819d725d1e3aea0b99bf5a6ecd1d449f2857844efd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94bc3196f2a077c42bd3c929c45e320f27d6d776c56efcfd446d5ca153f600353f4e33548a6be22eec7425fda8d5852b6af0028b8c9e04adace3d8e6b102e728f7bb9ab0718d7143bc24aab51d444eddbfb083db118de8d5614b9a4a20a2efc820e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49a4822054919f99df0ca6de11bbbfde532f7bc748a35e690573d3f48f859c1bbc4ecba7439034426c83f258ed935d54861c6a22e860ddba72d3c793bca3a55a8082d7ea8d50a6d050cb591385422504131ce9b1416bde7b1f66bbd7febc1e5d498a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h485da5abed4b0e533b16dd23e32572095e02835220de330a025c8cc5c20f02948fcfaa500bbfee9b052da0e2a6cb3c5ba84f8fcef6f4afc74b220764984f7f6ddd502d45da2489af001ca8702d4b621e004c4d0e544a1b97cdcff5ce5fad43f25445;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8140e8f72cf60b46ecd9f09c791507475270f3dd62ae7fbce2adfac3b5dc4bedb53513b7de1d1639e42093bd3053d254ca9b2e2198638bc576c11145bb32112a54d877f492896941acc6bc5c839f84029cb9bc3451bb611e2d5c120dcd296d38ae1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdff12f144c1e9a603e8d46b5a319dbe9e3a705000d35696f859a7fa571a197e6b28dd1627590cc951a8f324d424c6a4db8b4c8b2b3e5be335b69473f0b28d99c176aaffc0ddddc027fde64c6764ca6a12f43394fe0357c867459a094d27138103837;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b2e29c4b6ddc9a1c39430a892b7e15451ffb9dd0923b4fb9fc8d4fb2bccd1b49f5ebb3cd47cb9c912463840a9cf574d4e10af8ee775305f2b2cfe17eb0159b2554ee6cf398632c95c1a51f65312c927b6a396d124d20488e0d6fc6f90c3cbd6d8cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98ef5bbdac6b04d794e44a5e6f4647aa619269147cb9853e1ede983ba7e4283480cd21b7beaf8451d786c459e6f43e84778bf8a14e3cb18219438137ffc46306a56c0fbfd238242271eeea4f7ac13a2ef0cc5dcbf3e0433d57bd42d933ada1eb0e24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfcd5813188b512c3497fea6a4016ce0a0b880d6233e009bf77b5f767bc7ddd205ed1d7d2412699d1c040ae13f8d8b203ae62922f9bb02bfd187d772467e7299a0ed79e5f07d5f46d85944c2139e505a32b9e867cb8ec377ca853f40774808813b5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ef56b28509adde04dec26f1859cf4c73e5386b210378db4c6deef33ce5252342666ad6d0733f92908ced8a85d9ad2496a0dff2e68f163efff6f24f6764c9040886d3441393208256b30a62258036648b23b3a899bb035905e25c15c5bbdb4e02932;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeb3c4009197140e0316a69f534cf3b45ae4da377711254109f79bb158cd64c819efe897732d28d29b6ef7519894eb0cf44d7bf788299dbad6892d89a0735b0eee987bb983e859aaa38cc417ebf337c54e59ff12b34216ef47c8c7359144abb876d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab391f0f909123adfbae2d22562ff0f2b725dfb2fea1126ae8208992334ae7764c599c37eebd18ce135098b694a2eef2e25e27a7f6d0e9f712d8f02914fb0abd936489c7a3a131b4ed5ed64c8ceb37cfbf5bfea894b76480b4682d084157f8ce9005;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6fc4de13dad44432ad0d39dc1132e8dfadd2f3acfef1a1383f10b05b421a2fcf50506c64fbab82f9e939837c30ac067e9d76560e42ce7ece5db8b663cefa1c3d9aca6e73f16905c11fa88449a03ffc28385ceeb3487626141b0c02dfe43a0c906d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce8722cfdcb5d5110810a848e80374c816bdee46728f3d21e85254cebd1ab5c797b0f5216f7111fda573e18cebeef509437689d400df9acd09e64e27d8da080051ea7be6512cf46d4d03faac77c516cb380b2d0c831cb036e62b0e1af5af5d41fe62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a8033278ff95c6b7894d7516e1beac5cdb995246f99ebcfeb249dc8bac53a551012474f561b48f5bdb67f3bc303cbc359727d18156f062f28d3541f7fe03527d94cf48e20f7f95796bd8b80eeb23b00ecf44696a2cf91089d2a2e979f562c4225f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1cad92ae2737e6c03b50114d343726292e27bbed14d297964ce0e891a4ecd4ee597ca66eb8ebb17885c307c8b1761b5ce065a651616cbdd6fe96b6e5fca7e16b6f70708f3845c2406b9c49a97b263f1f890c4e19d2b688c2d04f39cb2c43c5f013;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61dc19940c059952b5ef14151abe42135046c5fcc4e82d66c38ec04422e451b6bb94a1cabb9bf75c3ccf7ce2b5bdf190d0efd0f0fd4051c70c6e660e01bb101ca15a21d06abcd0a0087afb2488a4cf59b85df7888bc83a25a0963eaddc3780337d80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd482dd4f39f2eb41cdf089b12d4893956565c1e19b9ed42237970c6627f2e2a4cc4c02ebe401d85fa7348ca0cfe9bdae520bd663226cb151e56c68e998a85d3c4d3cc6763eec766f554d115ba2f7edd9f668ce4575da7b5c0859da0f00758c13c963;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e3454d95796a959f4af1598909ae9f9fb42258af88e05b732fe0f8f2b3d6b89134b39b4d83a72aa3b199c108427d995a1ffdc67a2c0f60f74f23e86680822bbc08631548ef32b629bb27256ddeb10ff745d2babf5f9dfd0cef04577afec3f9cbbfa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha038aad5e821ce458253b7e6ab9d5990b28ccc43bfab6d9e5e597b53b5ee319cc82eaac151b5819fc849581f10ae7e3898f3b961d577a5f01046c630bcfe5a4edd13ac657cfd3e62998b321ed94212b7797960ad70870a1189a5e2a4b3f61c34a0d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d24b8e6574effabf400d377ef24294ce423a9e52fee8d63f82dacc9d05d543e4c8f58da247b539e4dde32cb74501f1868a017c88b1e0dc5350f1dcf8f7001b46ad5153645dafea8222c48ad1c388bc59415e73e34270e04988513c381bba7efcff8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e056da50b1b04d46715c39cc8cfd616c73d46a7109641590c3ab658a868d528ffce28c5d47de47c8c3a6ecceca1b2508b142819ae07e278b233703336440180e8224202e77090e707c2fe848fe85bead2f9bf9f31c6d348116bc79f72843991ed28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39ea421c2e184f814d5cb8c26cfb47d9fd7da66dfd9cc7ada0a8cd2bf7cd4f3c8201f0f9fd4f919ea3acf0df0d7cc01ea05800a5d6443bfc10bf90a064e2fad8fdd8416bc637788055a96bb8e77ecec8f4707ad8e77e9136baef6764da73cd1d35de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2efac091d4e4c261605c4b421a603e9e04319df9d823537a044ccf2af3a386199ecd1d8cab3147ce139941c26813361a16beca6e84b3d52877ebbd7f1dd4ff375d3ac9c1b6bea16faddce28ae29bcef0c220ed6b3b916ec9df2c4d1075750f7de147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ffdd975dc6cce5a94384e2d7a513f35e007b0a96144e9f490efc7d7469a3d59b3f19f2791d0aafd1960f6f719121fcf2447d3c1e4217bb7e850724b72e2cb31efdbc7feb386b4661966bf568e266e9efa036155573dc8a8786ddf8d78d9eb12f8d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee5e4c7dc639e701815c952909e0ded2597166121c9d69752ab908b6ee3d43b793bbfeef3e147c21662c501b2a150b16d32d3ea5c3ca62269ccb81e74ac1dba82b7e99ba7f26701e533d9fa6b2c3c3a6b7748a1f3b51b2df6aa0867db6bd215ba62c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55a5b710e2a36a9df61dd9cf921474baddbee1a5604bb0c4e3954c95d5f55cf46c5488ca1641dc4360eda7298ddee515b9508f9913a6d076baf241326c80476ea18209a472df6a9e22284983b739fb4b31ec69bb7424d656485c934829a2a187f1df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3ec26cb44390342cce28832a5b1b667ce459e9d8e7b3705f17e6178b50a8cb510a7dcc679eac1bf881d2ff6579d31d1130f16aacba3a4d30ba200b963038f64584f1bd90a7eaaa911a04a3348ba9a9c2b5c0b87df23352e5d7b40fce5fe3ff729fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d67a9d798c9e34baacdda5a6f09a9ecb836dcf00f9caef1d4bfb04dfc0ae13bd7e79b7c148f1b5f180bd9a233e1f6ccb4f65d317de95c4cd4757bf5e5c4e48e674ffbdbba9cbd65f690fe20bdaa949082bbc34d5499c8a848a948a18101bd9ceee8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d08fc8f9e0868d14ec2d78763f7d107ead72f8a64cdf51aa6a3dfc7545ada40c5caf26649aa5bd62c309ab279b0264274edcc8e41a391edd3b149e09cafaf8179c0dea199f85e22ad0c849a97d88fa2bb466278c0accee39fed0e2767ae40787d34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40d5998964675545fa055eb947188b682ed24befd1ece7aa4b93d9c721b3d80b10281f11c3d592010491a4161729ec53a56429397c11c3c66fc5bbe2f12797c9bea4df63fd527f402c1918a9d0b429a2960fe2a97e093143bcef54c2f58c3a77db7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6aedfd0836a5c83b4715412280dd370844704879286dba8efe04fe756fbf1b2cf0d9e37e59485f898eebe06ef3df97395427b518c82653319af584eee5d283d2564b205741b74869e9a7975018a66e399ef9b1c67b7c9a8a666f1a6d8528c140efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5736e914e4d3f4c3674f273080e22e462cdf6c6e52cf309ce7aff44ac981d129df2b42b1f5abb2802d6e446c18bb873240739fa6cd8c8e1effb361d32c435a33f6d6f9f6a098784bad82940c3a4fb730c8c3c6642f780889ede95536b130904ef1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedf8501fb1b22ee93dac51c6f20e3da067b1168984beb316a7483db5aee1a0e1cff44c8aedd15d3b73ee33aef5c91654ad469707470ec9801a442681ec151fab65963561c03270d2bdc7f98b8e8318256f20656e950a7148048065d0331f17b47cd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11677ea32e58fb82a563af50365f8fbf036b6aa48fc906a50e84144015982fc053f8a80d03f50e184cd488b1746efbdff28efcc31c217e7fdcf33f825af51002a2420c70006194c0ffe3c5e75e94fc407420e5ede3e66624c622dbf9d8f75abd1a54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7c9cfdb988156a14516638da647e27ae1204cf21702035df39fe384e515c509ab68eae666885653dc86fbb1f8d1f705e5a228df398951d1cb78448d34e26baae9a0b80d7b23229a9456f6632199c861dc458a240502d7347d97d62491ce764d01a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9229c5a7a5ff0a6fb5959e55c409ceb23ab9c587987e21a0a967d61adb25ccfd322380d9f5988b20aa19092abdecb42a44bb4047aff1dd81ed359cdcce8b156117ced7e0201ee0a87926bd9ad45589ba478c322de46d88926633f88f9a6963438306;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88f3063aa04e7226cae181aa025cad25e313e599afda2753353caca390a2ff3dd4b0c6e5eb1bd293f221623d36ed50b1ef91f8d82e04a70789975eb08f5a997376486cb93830c74494ab835409fc7b6483a2e37185bbcaeda6e01ce6da60c1dd64c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6953158fbea9860dea19e53e8fb562e482812af7621339d7602b27cf529fc361cc9f605dd0b416015f93de4ebbe8eb7e74c8a4cffe82c3f84c0b25fcc95d89c0bb864a670799492ed919190aa6324caf0ac8d00766d6c77a31f9bcf052e77eff819e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bcc817f9592e597842c491ebc80dc9e3cd12da226f467c8a5669a21a75d0aab8fc444344ed6764583a11cfb79c6b175d14551c690fba637de356eafb4b47f77d6454a8a9743259050fe72b6f8ae35ce0ddb7e6053ca1e5aec44e8a7e03dc77a038b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe8e3d7e058fbf1f2487f66aa2f58916731584ab6b55a4af5fe6969daa8c89c59d4a647fe21ce7bb0180c3b674dbe28b3371fd380df1548b475df6ad78e19322db8c5fb1a86b292e0f0e104648d26773c9c0d8326fc25cd6a410f2298d0ef60006cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ac9d568d7e7935b00e9a54421ab9f17c254473d994a2eae6507f9359e932b2e75cc5b115a6d84232c8cf74ada8a4b8f463e22510708a6be8c799dd846234eb32584b49a322de3a661781c00d75126654c754796d2761b5a80dbdae16cee2e22f8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h155f8370850a0cc4794ae1bfd01ca56fcaa43eb14940a987fdbad22a6816530da9b5ed65af569e7cc67e01bce0a62727d65a3e3fc1b3c8f1d12ed6b64d4b0eaa83d3c9e05cdf829e3244e3b713c71ccf9a11d6d5f096b1941f540300b159339c0ef9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h416639ddb83306cef31cf4964457b07230075422d2e36fe3c9b17b4d1b9bebbf18739bc3c3643ef8a92ddabfc252340d96ee91a1f4ce22bb5d24097d3e821e946668f770b74d94b671cb9f9d5cb76e889dcc5d3b2032551c9acaa5045636b6c528f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb757f130f8bc456e98f45fba2f9bb3dbf13653646cee5b5931dfc2782052b6f6b7329322404c1ef1a24ba520fad0747e7e510992c380c2b6c8d894dd94f732dde14da388d4f6821f13527fe17e54707b464f5798e05f20811930ab4e619f6faf4c61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37a10a0e943da49b8c5ee8a25e3138eac9c5c719ef3e00adf65c8881094dd9cb559adf91d83169cc1187cae35761352c2c45f1fb1b15ef084f2ca84be93bdf5b77f9736cdf0f677ed3ed10faf52d7986625bcbeeb763a2e540ebd96e6c5df6259a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c546a7f4b8d54de99b8f535a43a4f9a7171d72c4eb9c982457fbbe44f9faf1f061953f4f2fb7a3d4d1fc8026991334e6c57bd0e419b011cd89b2bd18aa913c1996fbebae6e025fa6b26930360f0cca8f9c4f57e738111fa6259856f1cce7c457dee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc750c043f9c158475e5d518cd194a787f1e0e86cb95055f4a5ed862445777a4bf752346ef6186f1ede00bb34cf5d6aa550c7b932b2d165f58b1512c34b5ec2d98221200e0dc859aebd0a17b61318c19e95b164f74a2a4356618f855889d860bfb70d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbec207f5ab4ac94c1c96e20af76443ff0f1b864f4a50eb39d60854d8ea586c512888b691179864270c9ef8a3853b06cb35c02c0fd9949afc60536fe2e6df4224cd4cc97822e3f306844b5eebbb1c19c9db94d349322538d90ecd61475efbd66458f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65d2784703719ba75110eb3effdb39eb03a66cc6856e00d35062c5fb2111c80fd37a5f06e96684282b10c6490af20d4b844d66b2b64c137c59b8190b34e610a047809dc8d02f08e782282c6474c1199f8f9153dfed0c88d96f9ab70fbe7edfea29a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99f942edc967325bf285bc20ea0702e74bb1342c938581e4193d15d68642d75e0135732d5c2e3658077d4770226784f31a2a0044da2f18bbddf27c8722283b50f2a1cf8906c7522d15f3372aece83c6abc7aad7d6bd88ed0c5bb22e3c387dd54b524;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc42df2c2996665c95a1799c6d9b3259078a26394da0ea2a4032e352771e96dfcbad81b1973a63de6c5e4e223a8640c2073e259ff2fed61d60d89d2df82040ac6c7789eb1b7c4f0fab642cf049053f11937bdc37a0c49e0bfd73bd471d708e4e74041;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b5b029b29e81f11654ba912a9d3178409d8f1ece9cee1a28ae9a9b4dd6ea357cd41550661842b3a22e4926d20429d7e455cb9aabd4c7f2807226ddc072938deb796845e9822aa2a36a5f352579f62093159c2bbc9b69e341371e4830a7fa162a55f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4336c29eebbf7fed66d5220384dc35e9a4b8540a611fc3213bfd37df17e86047c78b56ef665baa64e9588eb40aa7a64bf246ce358c4f9ce0471ceb11ecc6168cd1da6008d5939e633a7b7d3280efc213a0a680489eeda29f739e5d79cfdd84560aca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57bceefbf691145cf6d4bf6cc1d4c6915287c02781a3eba9d5e3bea97d5471a306530590db2a6b68584ccdbf43a508c36af268ad99571c32dd4c5dc6380e4d81abea77867e80f7ee7aa46dd69d90f70cbf2d0073d04e3536cd5674397cd84803c3e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f93ec63f5025b6a80d0419f0f760d613b82ff37331b7b485118e9a5fd722eb8651680d3ae4b3612230d60b9fabcd509c2d124ecdd9635ce4d2d9232f2fbe37d436aa1859b3a1cfbe1051e3181b00261fa381e767fd85005feca1e3d9805930a7292;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44781946a206721125bea1c8f37501da3361d91bf6dafc07f26cf5e8077c95caade690ddac9db2e50a496f0db47333a277e6a3e083121a2f61560d7b86fe171bcc6e4430da77b60384f2b2c23d6c753418c6c0e03fca3cb7d45c87d81ade2eeed0cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c776097febf2d302af9bb7a1dfc7e8e1f30c47a35da52398fbc82e96223aff9a2cdc9b29dc61b915ad9037f7df79012268b8c441d277149071ea85c2da787b4d7d3bcf2c3a319b08d1226c257521aab710055bbb5ce46b0ef6fc51403f61f8df52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3834a8e06dd47c67236ed42efb67cb11a31d8561fb8e1070da590588c335f0cd4f4f22e38a22b553361a5df9243876881f39a18c36fc1516edeb30c9e6a8eb54134cc114fd37bfae7820adbce046379add7263a4943acaea53876053cd40b4c9a05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf616deea710a1cdf5796e5f6f0adc014ab3552157a24bfb73273a94e811d8e163922d9e523a4ab2a8b7f1dbb40035a3cb9f895d038496fe8f901e2ca06eec1865fac4cef98a0453b5a91e9eb80273878b370f217fb507fa4317ae8f7616d08d9355;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h235bb18afd30b9e80a4cf1e1644e6fbb1aec9fa02c159c8079042a52a74a8b88329bce9f07cd758c941a354b71c36f2435a27872f7487a786966680ed2cd10f9e4b998e0839a78838a8c48571e6d9f6128956d08cdbc8c846c5a85cfb7fda3ddc760;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c9603803f546c7a7382c4567e75c0222a81c45f83c7bcf3729da4ec413bec52fc6cccb5eed5a3e0ec3883eeb5125922a926595e895786e6af8d22f0c59e15d6bcd7a40b4d6daa901bab759f9da7752375716879c42aa94421751aa1cc4be0d0eff2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1d15aecdfc835ab664e8015acf95d0ed279c688b24d6e90339488ee9f9398693295eaca12bdaf166f149c4361e43f1a5f2b2955c306a0c66335285bd4005c6b39e34b967b07deae1ba3048065d50117df5fda2e27a069b337ab83a62616d0eaefec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1681d26401b2e5b6b9abd6968271e6d8d3d68bba632e2e7c6b5d470df1bc34bf2570a8e7b3aadc7910be1e2f5744910ff33e45763c24c41462c5c158281d559c6f44e3493e509ea40a9c8ccfd7ccab8312ad19cf2912326c5a37b7a26547393f8aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48da566ca05cc6106721ca781b938c498cd3b85a1fa57e9c247af58af68675a5fe254e31e3dff6bdf5820d110b2a0588c5db9b2b42d96ec2f9c981c6bed5a8cc7248b088cc6ebaf3367ef702e23344ceae3ea9f69d5d0d957149acbd073911cec2cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63bb6698bc58f74afda639324e0074b180f3b5df8f9b507ff253ab06a8a202ae02a83d57d5dba32815b605869d2a0b21af7ba8242fa64332155c0af26858309aa93795aaa909dc5eda40e5d2d05978c029d22440eb22a81a2f11e172f8c95d16c9d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1355950181ca6f390bcbd24366da19225eb294cf0b12f4a3d4e7d0c87e0cde7683d6a9dd8893fbe33b4b513e2a631adc1b9beb895276dded10290c5f063605510b21e10c25b1cb049e66fb3df686349920d37da2773c46d0aa0f7e574d0183b9334;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a492cb1658f3d6d7c19c4d5f10e65792edca20ba68c562ba054f316c67b31de42a4f756b799ac2dcb865da44b6ad0a46d32afee13d34f5a871467a2c673fdd868a3ec330b7d058c5a53629f2adc0f320c096850c632e8e10df259eb408cb374a935;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3020a579e78012ac25aef7da79b6287ebcb3d15e4ad78073cdc800423deb22ddae567ec196821f94c332be690560f0c08654a3ee6560c773d97e683c79b860d7e38f961a101afee792552f3452f7b9859e87b8ed04bfeec9c7e4b9f8c2f2827697a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bcc9dab3d9ccbb7f1cf475b628de9932fe873e26a89a89fbd74c839574609334b58e35f3d5d90e6ac2b7b5a3dab014a93b99799cabbe7278b479b777068f10f5ef4cdfd7419f5c75734751307c50dba36caaf1c8124be7ce9d1aeb9a83fcae821c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d5adb32c4e78463a8f4845708bdc316cdcac194d658e8eccc3e8234b311c5c20b5148380865da4a4feb790541ffd124acb7e995cc573b91e66a1c6ab27a62d5373a1c3f44ba2bf0eec7cf8356f2781850cc3bc3afb7cd959b82f33bd1b5dcd155eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9d1db9d0b69253af718cb7df414d76cc995c6a308909cf2bc79e3f57724de72f89c7c7226d803e22c1f1f3f3ff3382efc82d5d65b2f509d3375459ef51210a80d1c5077857e0bf3ace9d5f225a8d722386cca40e185510fa2d62c4170952900a8ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e35733bb893dbf17b21432dd2f8f8d430f289f44399411fd4a02c6721b275e5d9eec956eea6fef03145a2f98457f9988831b34444c50d83df056d5ec91f7346ae35e92f7ceb9acf53a5929919ee2d80639637639c5c8db3f75c9713d197c3017146;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h794115ff46a4203e594243ed1c29ed63a5a5c1844a6fdd8109c5367ab6b2f48eebe6980f2bf1f7f76a8eafa763803bf158ff58b06d19623ef3a337f6251790ea282f0808861fa604e4bde30d0e2b1b73ef754bbcadcc5a943f52c5df5d7760f05cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd462f9fb605df6918f070b11032050daa2a520ad5728b6e94474c249b6a2db202912097cc78e13c40571d7b63a29bbf9d3b4c80c8353618c24c58fe1257d98069e4542fe023717b5e3749a2c3810274125f66d75c93897b39f4b769fb85b976add39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f66ec67f116455aceb9f81b150b3135d393db215e2a99b93252523516d19e9b938ee877863e22e6ce89f8bc2893e7aee74d8eee08a1f6e123019c64218c1b0086795c51988d148bc0d438e2e30ed3d75f5ff14efe12533b0855e8b6b1b1e206301d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ae1ca070e92992bf9387bcd77d274c289bdd69e01977c53fd7a32c1a9ffbbfa79009d6b63f850ddb28e1c0083535c52ba002b55c36a3c055f8d304117875c0448aa6b6ae2ab8d6e9b0f98e391a6fc64499bd56a0f8f560be5b2a301a6bb5f1855f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8073358a25c4f96465059a09a7e06f652c2cc05999224b711898f104b514cec495587d3c9190ca2ec39113313501fd80bc3b0a2b2317056d4bb4786b53216185cb9b32e142bebf7a07ceaf6a620c4f1bd3fffe3ef5710e55f761e10f6b400315ade4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc66b91e289689f5c28d076657d12d99fec5f7024d4cebfa9e3f4935b84badac7e63caa6a5f1ca70ce83d8de9a56328228d924c19b753e8572b1684e036c95ec6cb66b88e4f313925439d2152a554ede9de85912b77fe38559ea398bd591aa4d0ccbb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d71a60b8634745a4f8698f53ba7139e00c44f939bbd76eb8502b1ebb9d3ced375b655200358862a0262188cb454d78e82d3c51e9d6a7696da8253aa32da136daca89983e94d675ea27fa4bde8aa90148d1dca241e869e413fc8cf5861c137f1912b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacb03c4717d68a145c01c1b4b4a62a7041e336a86588c21559f4261e4a5dd1f1f8e5cb045436d5cbaca5f80a15f8a69039a1fe7948f74df688aa94815fbf9ab3b3763c7acbd3cf16f9dc645a0cb9d2f495a6f0b5ea1f59ebf2dea3ebf555a1ea1d13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d618cd1a7fbfcdff48ea7872ade036b1368c41a6064346ef6304f1ece16e94017740a30d88fc25416c10a423abb315b0400baba00f0497dd06a2033909cf938a86d3d4891b06161ca77fd41b938015d4cd42934d1089cab045656b1ccc7bd4842d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h648ff9a40675e6ea9c6cd3061a11deafb2f7a0bc759b761fadf5e171aa0316c5c9f6486d6716f8b0b46ee2e5ca2c733e1d550a050d26bf70d2c5f126242b6d14d63bbf77e86519e5abad834b029732d290976662750be7a5e632a0bf81d0f3901017;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3b80802003b50c70204914985b2461962fdea8c5ce43da7483cc9d03b454225aee5d3904854bb9fd19b81473724e35e58966dfde1055ba43fd0869c2c8c50db049942d9f98ab21612bde2db5e91d8e5e22d8a736a2beda00e172dcb93c1dd21f39d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b7a8d9da2edac0de1c86b45ab970cd28cada9dadb7882a4119e3653492ff5b5d9310772819a72b411e3f5d8918afc1027500ba34860dfed8cff57d9dad4ae44beb3601ced208e45c5a4f03c1a89af6cdb2d0dee0523688f36d6a1572c3a3da3486b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab97ac0c0d70198bffc73bdd1442a584e9553a640caa38d05a430074d78395be5c6cee015e34d9e33048ff26cf88d36611dd8352705f8264de66ff845e57a112ffb5b3643eadaa284182bd32ed340815bd190da9e378f7796a2c9fb2a15cf3fb27d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f3aff02e598bc5100e17073c9aceb0daf2d6daaf19377de782ef39ad18097d148f0922626441f4c3fa6831a99405f1b369644eedb23eeb09e8aadf330108de682c033b79965c88cd8c9a140e6086a24ca2e722ccf7d0643f2d39b1fe5f3cf8854dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3c69e573907d82a5b0f18b6c1c98e6140560eafa8d3e8a0e0f846bca03aa6e20d468e3b882b7c9d84bb59d4a8388387c6bd7bfaecacc7cc52157328e6dc2d6d2d8d2f6ce0abb805dc4b336bf707b32678f1f76a186732ff9aed802b0b87041cfc40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fcb99101e1d32b933f6a2932df82f3935ddc0c0d8ee52234ccc0635f2137e74d34b4e2f4c7aacabbd201d1f4745b682ac84709c7e5106db636c5c81b223307f6c876440b1a54a72d722744ed9da3dc7f5b00ef2969b0074ee578d72a1bcec8b3ce6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb079868b8ca4203c782f9e8dc42585c6a34c6b8e3b94b25bfc9f4dac33c707883a6ad3438453b97d0a44667f085418b1751e8019086877167ae3bcb2e8284db61d19a2ff8cc898d8ad6bec7d494e1a32f993885430fa829d1dd25b775904f87f7e41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b709133a2a59c732f0e9f99535435f2933096e0bd292f301691f08158a61664d568451bdb44dda12eb366823ddc9cd1328fbb9b94c667d992a644c1f1e98ebacb107370e7b6f7a56185ba431a0bc72ede449fb6323af779d1cb2bfad86499083f34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f30f4620fb6711c8b200d73e36f93c07256751174fe141e515ce418251c3625205ec72cb69a3fbd8c396f1021bf954bea4d7a16de0a271e635b4f840efbfd255c4375ca1ac4d07548ca03d2e472653b703ee77eab8dec3478776b49db66a38f997c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c3decab3de1d6a812069c7fb0ec9d901b77b4fde257589eb6ac8e94e8ae92b82863c81697d59c9e9cd02aa52166013dd87857ea11c7eeb00d45e870ebb84883cd02d6f486e25b0aaea59916be603ecf4bbafbb460241973167f6a0e21a87fea3843;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96b1bf14ac5d1b2cd3ee9ddfcdfb15ef9362e94335343201c3f0f77a7df22ccf460502b921ff732d33c27fb3eb568185da046f3175873591107c0aab93bec827124e311bd65114646e1bfb47790a6390d92aafe8d12e61a16aa38a61ae6666beeb80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ad5ec6033e5801fd12418ba4c4774041c0ada1c36a968c18c5761bd952f3f02a95519ce5bc82811c5e2d467df25e26d13c28cf5511c06002a165736bdafb0d0a679ec3b0319eea78e2bbfc1c6361f363058dbb79ebb9c5f4717b97edbf73e293b55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h738cafe4c7d49475bf587ef4a5d9bb5daeb032c09bd1b65722d40b954b7b4c0608e41aef56a02dd2346d72259c5ec03e84882e1c6414011b1307d78f03f84cd737d0978812d6a21abbd70e4c9b409774eba4f7fee15e3d116d060f3f1787f5e12edb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77b3fe0015261d1bb6da97591a631e26fb0908c82cae466a0979af5c019a097c83376679fc89fcb83972f3a1593403bb2a308acabc4c83b519dbb35f6846a5ee3ce5bc59a6f674c031924327ee5f6410fcacfb15ee959565c01ba5e2ef84b61ee10a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ca4bd62bc982642ef78995cdf23ddb3fb91fafb4dfd44619ca043dcd00a33026aa3b851d3f34eaea8244ff0f72838a0eb097da53d6dbf74edce0e7d4dfa7d3d6c99cb5b27f728f27652346323d09bea75f14407b9d6aab93354f516aae273721109;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5c3000c899a85ccf9b003bcaca413c6582c2f0000584e4ad339531af5085dd56b7626c619f7009edcfc1d476556e32ee76eab68bffbfbd970134ffa4ae57796b37491b3191c0bdefcb7ca63e543f95b13a363e89e7e0a6257d4e59430dcdad53c4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35b3538b560360c36f7c6386c29b49d08d94e3d8f7cf1e2d60506c473e508d28c9df9df6b7975b2ba7c7b5c0f4049eb6256980ffe3e320d2fd58e14aa25ac268457243bc8a2b9c5c2d980f0d84d4da86e024bf75c00e14af8ed942b5e92d9678980d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e6cddd2a720446e653e68843afbe25fcca8ffe2161129da947fd167c25a8327839ff2a12f648ee64d24c4db60ac90dd15f69d902370d85987ce678a20ff4198346fde4a33ca9a4fde4ba0fbeaae0d12789dc4d7fc45e1f2d788feed9be3058b9a2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bc6765e79ecf4197975723c43a0073d485db2e8cdeb48306aa7743f719fd9efaa1c46fb948589c465f04c55a4e4ef6bb39b4fdaa5061d6f4bc85dbf3235d05c4fae1cdd2a1bd5068e31e734357c9da3439a2bd526f37c95375efe0898d9f80dc90c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79c8211a337d42582f9015e8eb4a5e911a282b598d089505622c64f3b956c83802d82184c2101e52b49e29e96f9b4be6d3a380193882714cbfb3b9b88e4bd7168d88374b7b539bbeb3ee09c7aadbc192b2be5b578b2a79afd92de09ef801f324d234;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f93f602367a50a5ab1c41530d7104e3f2b3f44ee3671ecade41e7f4258576ab2b8b194850a6c21637ac6eeab3cffa39aad5e88a1047f7a4fb6a05d65e424e42c448abcf3d8ab803278e77dd424c8b2c02ad9917216672a4615a37684cb8dafecf74;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c2c094052ff5d944ad3dbb9ab3f9d9e81f1590369e54637e8989b518ba6d934a3a4a98b3a217063ee6e28b5ee857ef9a9b35b41afa5348c14edc2a11b19af010c288501465c10b81fdb4964124799a5225c6ec9575b4e7b554b8de6a62af6115b7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h999bf3d06c419ed08c12d5f26c893ff92777ee36e93cffcdbed68bb36b8fc616a7554d44a9af356d254ff03eeda33e73d7e59d5c8c00e54b873e08fd2bc40b30007e08c787bde611280d56dc1d036ca76231a67e080f22bfcea401c1b3f64a220abf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5995f5bc4169f2256c4720b4316ff4b701dc0548204ff99f68add9851ec355e58beb08d4e4cbd9c068d6a37f394fe1e30a59a0379fcdaef27113aefbd51b9832464b6c3efd7ee9f76fc7fad33b9a6808ce19fdb35831d3323c845c6adae27b2084fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7552deabbefa592dbdbcdc3508d9832963899c6df8efbca3a5db36ef20c8941c3dbb544e3234e833e6f6dbc45145888148bcf2e793bd8c50fb9f03b9dc07597acfa8de2952c177ab8491e820c2225f9f9c45bce128137e161fdd37b50d70790f0ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b04496da8f548788454fd00b5129ce1057ce2421b4430f84a0576a0b587365ad3f7d40941f06aa01d2893cff53d8d61c21c1a6d76746f69d1ade1041c7fe2d11f08fa5cbcce03a04273893fb1c1b30244edbfb33815f2816683c885d7461fefcaae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4f11582106514c8160f4cb4df6eab7bc4a337826cae72c8a94b720cd3b825796d547d5e839981b876162cf5b49fbce0615321f8b9662066fc321973d5bce2456eadc1b76d01baa87411c938f738cd4fbed13a1a473b9bbc2046cb1670141cea7f04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7d034447cbef55bd154ebb628c9b0aa082a67a4f4ec1ce455d2258fdae2fc5008f9adc25ee01730c6cf7d4e15ef002a8d40969962fb16fb415631dae400b3ea412a771c584cfdacd502e39173b27b46cbc6c402bf9fd7d4d4b8da52e426da220e47;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h797b1ee3f560b9a792e3ab020e4171bffff312d4cc893aaa6aee8396c61ab61e962ef5df329805cc944809124cf6662455b08e3a4baa85e24b4672d419e25ab0a7997b3d1df2fc32e26fef254d1e3dfdb2a3bd1be6ce5db0bbb02217480f8a558120;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3df24c23f9c51c8ab77ac2288daa39fabe46724d1e9a60f9b289f94f46c240bf0bc6b0e6cac08ebc6439bd17b2b6d8d516ca0296a33c760d44f8c1bd5697920d8d04d7989b91aff0f04ba27ff230f6a03d2312f4a94be0ac0d9738b385400e647c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc425180d5225844b125adac95096c418c211daa40361ae24bc41c80a4f31d958d14b8296be8989d377ec2d89cbae18927dc684a56656ec574e7c840f05f45182d6d33f580abbe305a8e1d2b02a9150a591aafb57b3764297c8a549b20bd4ca3ea467;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f1b73da94f2fdfc888c9e66ece1715822ebc77dcacc10b4c4cb1369f4161d79355c7c6371865b54493606350951c6f040f474684459963d899503daf78cf6b789b05e66c987a2e8e3d101c7805704ec6e9edadc49ce0e11d31d976a1d6e79c4efb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aff3df3df9a1a0cefa1a5b573c4729de84619059cf5356cbf7626910f6c5c1b20bffb3bfd3cc63bb6d34aec742e126d7071bf59b7db6a2e16938f8a8dc93d2a2e50d384307d69af6daa52c8f4b7da7b89fac61d37fd5f30d32a2c995ad2cdfebb40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5f5bb6a4ac848730c6458c483a13e6df9399a41a64a0cfcc4b702f3bfa91a0cc931503b21952c7a57c1037adc6ee435fcd47db6c3904400bd7a25bf20b0599d31bbefd9f2511768b6e5478faed0d050b74e8376b2caefb239c142dca6ed8c7afad3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha63c09c4072b70345899fbee1e612f2ca19b81e468d0d1c3e8c4ae07d36ac82249278602e4763d85b5b8720e3cb7b34c166571d47a5dc9260f746ae769874fdb5c32466d798359f0874420d583e5eeda33125a1a72fda7c49088a1dc367e21c86353;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93da078630c5f3dad7cbd738991f40cc26039cb73baf539e0f78f2378ef38a59070307aec447b2d07e35d56824cfbecfbce01cc050c9389a237a44917da831a91ec72cbaae091b855271c3e86f51cfc0458140fe7a67715445ef4236ddac27c3eda4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ad5efa80fc1afec61381aad76e96faeabc7150d68ce569aa0a204cfdeed339c350ae94c95c9618730f3ae0e12f0a81955c37e681d1271075acbc7655e5f92eb5614425b18dcbae0f72fba8a99e5b52697ae3c348d1329a596b160500a897fe4a1f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff05d75edfbab75859807c5704fdcccb65f8ef3a627fce9a23d785ac91251082e31c8d33f8b04718f7098beb7b8bb5b84c973df5a58fd6e343ea3596117e25a90cb961a3214ee49559681b09fd72909a035b060260bfa7575d234e85db864c82f474;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fa02480a3819cff79b08ff837edf990c82bad2ac0ba43c8a983cac79a5623818e03aa7af9561b3e8c271cb5bf39ef5aead6d7fb74132e1a7f8fdb752fe105786247249bb498e0659f3cdd45aa2fca58a2ae8ebe0b2f80c5ec13790171af95b27608;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa1518dcf9bf0015c540deced541c6a3f2cb181ec7629adb53dd22545e5f49f1054e6011b25a0c875cee27294c47939efa392dd6353d8db8a5df8f90234b15794430bca9a04dea81dbabfbfe91f6055666e4ef437154114ac1962462fb8930e02da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc84f6a533b39bc65c1da2ada3faac266c47a99a19f0e35e9963ca16024c1570824efef6076ef782107ad09b0bf26064a665289a2cd121c2bc85059742036b1f154b968cc406e5a020707b2fc1dde1f608132ab8a366ce539f57cf3b4a5b2117f926;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3db033e481e71c31c3e881a06f1b5cf3504e93ca8b59aec1559bcdd9da4da63580863f78d677f4aa06facc8961e551c6a8815ada11e9ecaebb2c4bcc9c532e8447d6faf573bca721f1be260aa0bfe18cbd43bfe3d81778d57e362b229e2058a7b6b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb0c7620739babc853caaef7c18deec6a82cac4173f5620a3498be2c806adf704882c4cd8c3f46eb6d5c50423687d3b18392b04d1594911ac96635a8b0381bc08c1a73a544c6a1a111f4ad4d1c63d63ead0e6a67b7491552503c2c12af095273965;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e513a73d44829b6279f2da0748ff2ea982b0d89a181e5edc66b7a5e06feacb94241821797a08ac4a5693cc38d89024604bcd1fb4657e458fab56f0000caee1da02462be47a0be397e2c1581df9fff56132944eb4c7f4187b241d89e8e26f43b097;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e1ce4b681d8fe2baa12f3edabd87f3d8161f4d17a0671bfd504ac45d23ccd8249890c9855e23e57fd754df466aa326fc713a1971888cfae0ae45ea420c75a0709fdc721ba422d06594ed3d360420b17501447d68198d3df44eeef64f093828ace0f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb166c4ba3085324aa16f2cdacb6ee6486c091f47bef338642f11b0381be2417ca32c9505fd965e5b1cbd2e5811110877e1822cd4ffac2bc7a525204fe12b30bf72eeacd6a1e49eb4f8dcc0de13d7af1726f207453d6fc0d4c616707c6bd60117946;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc958f0cc8fab117c015f0a326abd0b60dbf414c7ef3fb08b11fcb460e47de402fd1ef440f20fa802f82ae73fe85cadddb68891023337e77d42c45da4c757c7eacdcfc82be1fcacb3a981c6b4b9ed33e1bee825a64d2176e0131890b6bede13fb0434;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf618ca1286b61b5ab1555f010a06b4bb27c6891cbe60fdb7b5a194a1628c3c57ba1d1c4983d298926e488c338625a31fbacddb70d5b664b05a7066afb352df094b5934ce132a011c0b166157e5921d911357b19e9dea637b39c349293fff342ada62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h249e119a621ea4dfef43530a8b8550c1c7c50abbae48d4bd8ff16febb500fa312deac5c294f3e488207ccb126e46ea875835c7ee44b478d8ae4ac1a65a6ff53923cb85342e6fedaf73cb1a7edb0b6e307d6d8b38c8a04a382247422c1bcb0de4cf61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56e6d526eb960545a2201a9b10061c6203e42c48655ece7f8b275439ed0b1ee0681ef2028de861f9d1357c5ef165fe69fadc2caaa4877a9cbcb28cea0a456f53df3cb9b0ed9cc4e2e3ff03e57e8e25a62271b8e28267a76ec00e34e5261bd58523d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36104b76273e2c2ea84169a42bf154d29383b7051c4e0f8fd1de710f785cb7af28984c8c573610dbfc7d3d21c675f55f2622a767041d989ceaa0cc9970869e1c30bb7c2ec7976ff226c1458a4a245a5fd998afc02952d4cd4aea9d359be826e9246c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc1a6239ae21c62ca0a913e7bcf7fe024431870d0e1cdd69a57b52725bde6601aab0d5d2cffa84fdcbf901a2a1252c89f11661dd929d7ca3ff2f52c165598b1729bea943fb64a865d61d5b9bd988d02a6e63e024185f94d6d58d47c3742ede3e193d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8372d22aa4974ba8b9697714ea509a5d3309740b7c4170a225763c70b7a3ceada488a696b2f798c0595e74b6cf947376ce625cb59cf4359e0cc07893cc13db703e46bd737828b6acc0222a07d48ae64d4abcabf45f5c045734d3d5f3d1095a1039ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b29059f1a2a32e1348e3ffb4b48ec9a6433a93b74944a576567c4caec22a12e020444433e2431c746a4af320be91750c2819677a1f1d53030e1c9b54b7c51440b14544f8132c354a3713066854709bf866ff61a46e896e55148524e0cce15202f1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7a6a94ce8fb384ee9e6eacb023ae8a053afa95163b9f42a208b26ad11c1ffcbcb634bfdf4a9b822390e5737b2c9bba3feb05310d7510c4685c77b10d38fec197bb23eff89fb6792d43a9ebdb2620f2777d9811a74260f20c183f1014bf1b7798d07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90c75f5ef4805e1419c3aec6f27bc12a2f55f751a54c31509cb5b0c0a4fab796408cb2f6731f553c8691d64baf0aac73268dcb816850a3238b7be1cf3e2a575d500274bb1010e71e4eed6f213ac4ed57d3799349d2ffe99ae2998c553b8ade0e9d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55fe4428f5f9b1828db384cea24c129c9158de000cf6a49e5a20aeaf07821f93a1a434051f64008dcf27734459fe7d9916d3ab2b7608c75fc9a188420e7b9f07f695f5f04c1c2114e59e246132912e9c7d0ff1bdb4fd3d8bfd939cab9ef311a1d7a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2088e8c6b25c672b15f301929104f260beff0efaf29647501ae04df66b2b8de0c23f335b35ed66d290fe4b8ba6f18c7d88597a7261033fdcde1f019155c4f76c1d72c77e00d2bc29cfec18d2260bd62204f8477a82f0997f242fbd22b8da01a02b26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h505891ebb531e66572684f66a750e990ed1df9ba73a8cd532caa4fdf436433017a7bdae81a50f33bb61418731f8f79175613520e07f40c85a8fdf5e87323cadeef68e0f694ff0310029ebd392eaadb4679e9511d0068801629b1e59a20c196735a84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d066ae870ff8b6e24f6d6f167ef06770385b4927d698eb7b561ea54f3e78a7a22485f8159764efd92c922dfe24ed125906e839bd225d1eafccb6d335408cc644c6a88fec659449b86d2fa5bb992f018e45518bd8a18b4479a7d8164fe11a493766e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60c5bb202d58392f3e1abdce57c0f6f1000f7b713d0a9751586e2fc2e42f09ff279d0d41055ba8866cc590699d3cfd2883eebb656034994ba359cbb97be6fd44551bdea9b7d3bd60625ef99a597c51118ff79b592a44de23f9ff2531ed21e64203c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa5f2d2c357f2733091174e44a97a4e5243a31c22b42dec3c660333e9fdbdf895abe88d69783888f00f2e315a16d17a9fdac5ffd73550801326cbfbedd56b625ef859082b92f3f3895e09cf413466db97d2525022fd7a5fefdb036d92b84503bb0b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9063b6fb13ea8172be9d62464d8f1ccdad8d50440dcfd1cb87366a965fca4e9834d848f36f341361474091de03df07fae2c2b241dfefcb0d638ec56bace5a12ab7da3d4ffc4b31a9b6da116240d8626ca3b5fe6bf8d628708032aee5be532bf150df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68a2014c74b99231a0d8bcff3b353f63cc5d1dbd330264f7479f22282c800995a3214a95362a1572d08ea8e26ccdc280cabdd8e61656617c7a756b2c68c28da31ead7c54ab1dc3fd71dc806b2826e44c24e822a47b262880d8e9ba71f06a30397626;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6f98db08c3966b4d1a31425da39d16ed87a66da79b2c83d5d27133a99287e499e0fd5b2a6c2ea6ca2d820c39c47df1702e4e8269f1a58c16a9031ac826de0d93ea6e54e8681b93f1e57e6ced771da98d80342ede5f9a535d11c5dc2f56fc8312b38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d05a17e2d7073393c215fde880b92b602dfbec4a55bfa16af6f9ddcf16d743b27d797c3986367758413dadf58180c8d964ee30c425326867e4872fb99e86176cc4c7f65fa5d105d822002cf45c0bbdeceae9aba2565b884aa4daa6d92faf9f03e70;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef6aca473fbfb88924947d2ed85a07c670f2d959494b4ae9452c534eb21fa51bfcd6bac58fd029ddba9aa2c4f3067bab605765d43b640c6b6a613db68f23a0fec35762e6b2325e13f8d46d17b8bd11d287c12889190c942744e25672829a01a23ec0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee92e8fa2f726aeacd9c85046c8d749db5d3bdaf9465d2a14fc24a3c7cb9ad10dbc1d2a5561c8cdd4a06c71ec73c85939d59a9516dadfafab206f26a16a2bb8fc68ac40fd7cb50023bc4b9b4d087a18a1d4efbfe9122c79a7f8f60ba556249d33ab2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c28d1c824d5579152f4ee44eaa59bbaeb0ad17aa7eca015cf6886c948789130d41a3c9981f70a3db6b2fafe5ebacf6a9cc354f37de822dce2d2e908dabfcc923a2bd373d3ee13e99deb1eb37b5645fbb190caa7fcceb13f8723739d5847bdbebc38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8729ff84b08a79c2fb6e1d18bb12db122f75f52309f2122607f7e2e68466d1afe8f58ba3c24acb77ad580551693ad97fdb472031c27c199487a57b813076650dc9961f1bac5d2e3e34360b064b114b20831d23af0b44a376d77558d1eec49f1db615;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cbc3fb7c6ecba001f841b993630ba0fffd9e94d757e1add7446a01530702888fe4b2213e0493ea528b89874ee6171f2af318ad5c4ea089d99c56ebe2587cb9ad9b731ec807696e9b4f4ce6aec600a6e44373d36c777e5a2fdd8ca8322a41d701fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf28c735973aec7707333ec94bc8b49350a66d3484fd1037eac22c8dd55d16c2e763414cc61d43acbcd5b76e2aa9870a6d6d4f5de5060fdbabeade325039474706f6cb4afdf4a54232c70369f2db259cd71989a1355a990dbe147084169c388da6f68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86619e891b3ff99329dcc18323d4456163503bcb01eb7713a4b1d84be2df0302da84f66822b3cdbf0f74c5b17e010439644cdb0454843b6eb43610fc1349af833cbd4b1c7c00e2466b5c847ff022c92d713c723ed9edfa77a39d47631a822933bac2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92143f5e86390d51ef67102f0678cbaa139b97ae22a69222103420de7da770267c8f3cd0ce2bc44fd6a42dfeddcddf880b9d6e6589b15e77b19bebd9d9b15c4009bc07f3258e16b31c5521c27ba96aff53371de30f1cd3e3386228358f2981d5672d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h683e4ce6baa2ea7db5139e34a9fadff93dcfc61fd9130235b2323df68446870d83944bfc2d7f03dcded4485af7789c66f5cd87b0e62d5a22cf06e2942ffbd63e25d6d09a714b593bde5e6c2cffc6bb8d12a4b3f62eef8bbffea365885e812deea735;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8ab29af1ccb4678c56ad49d2736f5dceabb61cbd1b0218dcf5327f26d9c8b7a2fa54a9e847e5f9144b2a7423327a11e16c2a11a0cb3046bededf1113e951ca01031a8de70bdb06e9a93fde952e51a171e61f04338e7173ef2173f1834ef5d5e865e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba390789de0e89efeb8067ff819b3528e95963fb5307b293c6c8f07c6786aa9569b4563e1c36300809ad053218968799f05c7f7c664f68983ecbc9898b702586799f7baad78f23462249c06762ce7d0b575b824440746eb9c719e6ae5f3d095cb557;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a64865798b68d20cc5da72f6a2f653a0cff127ab2f143b512ec1cbbeb26a0a147b90427c8373e8836f1149cfa72fd433d4c31f36c8429d75be981bc21184fab0096f2f22bb3b2ceea0474c43e43144a1c5507ec48e403452a847a298a8e2522bf51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89771a8f69bfd58799303efabfcfe3ace42c1d442efdb769599fd0b519305234406445ca7681d83f354eb6b9291b771aea58ef7aefd9339455f22b6fadcdd5ee108f848442ebe2ce468d23cd3292e4bee359b009c5c521b133c1871a9811e00d79ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h284a4b237b32339230f93396ff5ebc8b8a38e8ec9afa022009ec8ef907644f052b3fe62fadbe3578113236f7dfbeb1d78667848e2612a9548a0a18042fab56319d17c6fe3ffbadb8cfb2bc1593d78d66f7dee2449b2eb92f35bb8cd379497935c5dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70c170c95da351eec78feb92ac6416c62487529396bfcdbf0df9b7dd1b1c9ecea07fe9a8e65ddf4b8a1fe0128c563287cd3d9818c81fc16b3a25131793d706c6356932e7f71e7674c5becd8cfb39ca8726ec7705e85616754da6b4dd81f4565a42f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8499687def714769364317bfae94c0e367590cede306bca8258956cd016ba4721f8d7fe64a74e06e6cb14942c48075b63a331eaa31c59a1b3fd5f6f61207f2b4ceb5f5ec883e78cdc2d79975ed6431861cb103d6fce04c38d937b30e8668542d2c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h998913263bc29e278f3876b87a45068b47723c5e1399c10308e4562e44fd0409a3b9bd9a05bc13bf5a1a1ccb61a81a9de57d37b4740d21a2cfbd4698a74778f22434e861830b2075f9cced63217554b4836fa588156b854969ce89dd48804dc624d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f44649590fcaf9b44196ce4ef9865a542a032defc8bf8d3d4986c64b8b8dd4df065be2e4da6161ed94dc005bfc7cd6c6ad035507d0700d078166b2057c0ee51641bdee66ccdf760bb488d36f4864e1f2f967072c1af9b6d5089da8ea7a30a33cdf4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h815363f7c9a3e31fd98ed2fabdd3c954cacc569ffed3cf816a2ae385a8f6cb71385afd359be8f1ed2f49b2d977f117d0ae753b49b0bef0c4b83d1f5c610dfb90c3c45175b713ab072a602616e15ff08176755c7e0a63cfa0b457f5ed9a30052312ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he123f8a9f0074027e626bb6c8212f022b11cd4d8123f0eecbff4d17d70e8aeee05bd3b45886f2a9ccbe7920397230b77c620e8024ff7df2582f8ddb8e487ee00dc3c7640ac3fec0ebbc29f975a8ead1035b8ce5fe5150306b0b64fef5c23554d1563;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h269a232e1d35926684437d989fdb26a954b7d8de2d571b6dde8878c47321f1818591ac7fbc877b8aae383b12af6ca7fa7ab0e2d0f4f02a3dee18c3dc5df8a23f8eddb757a8f72e115f8c597cde966cf5054f81d496679ac7b717d48479953074dd24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5134ce5b29063632716d9b7515776c32fcdbc7a7258069ebede66c09555bbf46eca70eb0dd4dd6c4f01ca98c6478214004f8aaea4ec510b92a33849eef0f8025720f2650354f48f30f4177098e7f3a572cd2c21afdab89669e0e0e10911ddad0623;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6335951e95d0da1e01e2d09e71c1e02e35029a036684054b2c1de1662eb6b5a9e6445237d5189f0b74cdeb8fe9fdf906608a1d8479893b68307eac39cf5c5dd2990eec034a3597a3f27501a51e601771aa788af99b4c57f33ca128d154e314a1873;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9becb78e1a8378c8cbf319612e36b92982f650edffaa53eee2959759bceea5e3bc245c6ff0db95371e7810f34311fd52c08a499803773f242477840357f1c918f48074d1b440813147aa1cc292c14b41a8fee83fe5c219ef3388befb41a0d2b0c59e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea15d6e7b5d0a25253b2815469b2192473c046c8b0ccc1557d64afdf21c4d8d373de8494be29b4185d85025977e1cff6f7e0699f1804ea692ac977438a950f67e799a26c96435ccdaabbb0d96897e6dd983e8a243d99eae0ab527913e916809e8186;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h266fc97d99024df7f4292c3f475a623c27b3d4e08be245cdd2f79f886e930c0074e00a455ff0e614c34e1282ba48065d114f653375934560050281d79313dcdd7cb10f8f886ef5020dd5772b8aebf749d38d03cfaf764da03c6302aaf039e587e911;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bfbab9c30d6153fb28285b058753ba998d6392fc33527cb533fcfd82e1b6661f549ffc13b96f780723ae4153700bb28f043d3d8da1e8f2da9ff5abf3f6880a238b4228eddd1b714b839d092134d9f8a1c16f024a50d5ec9113e83eed8a3f913265a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4daeac04d721177f5c5a534b1b4c0215335a6b25958ff3f9521245b05f820d88c24f2bc602b1e3e1613937b9b918960f0ef763ddde28759b6250e3dc525b823040ccd263410b014ee4ec5d819623f912fe4c826aeb8e3142eafa4454745997eabe7f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a9d6a319827d87cfd23cbe971bfad5e84d280321e575a24d01a60608e8ff0c21c52487aae1482d8acc76be354fb6849da8bb9421fd892406c5355385eada736361e61561e85a7842e1f7f7ec9405ec66cc5ca30527e94786a9e026542657f74d779;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda63af0a3ec6ac077b55f5ff80ba2e706c76eaba3839d46c94bd58f50e821e2d2e04fb1e3f8b4302cee7b3e47f7e3a6364f31ea6841458c03617d1f7dc1ebee5f99b611d7e30ad1b4edacfa623208231f6306e237c80789c1ef37eb49fe91803eed7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20ad96d6531f7e18f8eeed254fc2c24352966114977c33a17d169244b9fcec771cb366171150e7988e6a77368f85fa32478c231f4d6c01185f69ad584e52f5f69a0a0a88d4d4f79ef83a6f0efe05ad1ba3cb04aa06e55279eeeed507a6e752e0304;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h265042fd8f3c88d0558e26c2037a56d2265f4fe1298ad4f42067ef07a4b5bd0f163c59a4740d35e8ca249aa3199ff151ed8ef39b9ac1077aa2465ad0d547515fd399928e6b93966e30d2664cbdf8a89d0801b9da290563c4f4c1a7b8a1b23f736dd6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf99927500c9372e3b1655f69d1b993271570b7df5bc01048e3f624dd52ef707a46fad961292ac7f987b07cf46eeb1cdf3fd92a9cf4eb14d2736423e73e70d3f3bbd5ba93540c5a2683980b1511a6ac2e4aab8787f324b22d4a6be28afc71f8919c64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2385ede05da80ced2299fadd16ef57b9295f28f66279a1608158a82b2f376d38289d9e2798d1503ee575fced1764371505557987b8abfeedc0cede8ae75e82bfd214f9bff54d49dcbd1b3994981ec8c0584d91fabb7689c8da9cd1e64da76c089bdc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d2ca6a6f75a6e80ba170b9037632ea303a5fa2ee8e432f1ad0689098cb85268152ac37ec195491c604e732b616670d69abf8817de5ae30268cf02dcc39e7cc3f27e4fa8a7b17c74f9170cc8584d6a4b634838f0091ec552478370335d2d9571a9af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54870b71a46ce1034ceb613348a3308afcbef9f58e4099b8e638c662551c0833fd9a028683dd5ddfd240c1353198c39e7742d68f5bf3601ad9e36636aefbf9dced874b942b1f1f797620024d9c4c90ad176d37f2e228895abea5e3470c60bb781bec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefa2d982a6ffb866f75f62cb95582d1f887874ca2f06d9d40eecc96f84b586dbd5c9733dfb361d96cfc57c470b0133ca17875ee07c7d24ea05bd72f61246d2546ddd5e7e5b4e77aeb67aa977ae63966ec340f2702b0bdea05b2e9bbbce25fc0c64d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb90b9c1a009aca301e3dfc2310a3434c3f91d79210952ec54183436597ddb4f7d9c36295a5c9393b68eaa8d405ab75148fc49596f31a11e026ad88957fe703bfffee9cb86e59a7a597fb304c898d13188ef81ae77b38250462e17ca860de022a08f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b6bfb6a549188ae4678b13b4c49451c93873314750a2ef3be0acdb654802c6ed391416ebff21b0fab72fe7daa314decff3b0632870a4855c825f08502ecd04ab726ba02378b529acb43669d292a1b81ab6813f79caa8d1c41d4db6d8caba76ef64a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82137dc2cb888b2d38949868a3c73bca0c4e00ae31a298f38700c632e7b688cb97ea2c4710b677285f9cc7b02000280bec02d07ccdf88577027ef345cc43f1549ffe85d3ed85c8144aeda9056634ef409a1a2db2357fee33c7ab1ff951df8cb3318b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4a118da9aab8835545655bfc8ba0420082650ea9a64a58113adad9f5f4bacc58c4b012524a53ac049679057c23b7bcf16f7235a0858eddb074249d7ddea186344bccbafe5940b79d1e26b004e3568e38fc7a6328eee4fd9d7bca4ca2ec2109d42b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb280166ac98b0a29f51791d21e3ebf3c8b154eab6742e4b8d2b95434500738a92ce6d52867768b668865b775159bbf0bbd231f2067e88940a223bb1ffb166b6985881e2db573a7659e75034e300dab69b85e57d360582eb3cd6c135f2e46ba4f8274;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa1ad18f876e0ca0dff3d2d82170f818f53683da855412e88a2632a597eb91793e6617f7f068b476688a88a3bb6b1fdf01196b48c5c309dc899ba779037d4dd59d9e6a1db7e385780e443cc5a8a6096f211b85c4501027dd732440f32d757ba805e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf66d86ff5313187481d1f28869964912d14953ea9b7bac70b4cf600bd90fafbeb377795a780a6a50be87dea799f7ed1c0e84179e2950c330a382932923326e189e06d2c09ea4f4e5fb079445e79db060b123058fa6a4a50a3c5c4357831000ee0896;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h565ba0fde89ecf3154eee843429a7095f0ad068aba4207c38203415cef73c0e10b47f4075ae167b39c450e8d329591a77ad3e81a023d09abde7f9791d562f1fc95089c03be1141f423294ee39788df48068d5803a9fcdd729b0f2749142d7694af79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2f57e3bd830a64cc543e4720ffdf7f564902a525c8200aef2a238a730ac5eb2417acaa719d22cfba017845e86155994117be6f3bd8838e80dd9175fff8aa9d2052ff15af014e6cb6de55b085089fbfecc6e37d8f963d643fa0031e2855b935ade23;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55a1ad7867197f49bad42e84bfef650b3962920b578b19e4373a3365752a9c42cef50a2a925d88219f744cf3a15798c076aba92b03fccf7e1cf56202c8fb4f18a3da3b9b3160d94ad2b0a99bc1ace4d373f512435ba37fa9c3c0fc95e08cc5746911;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31d969e7cc1d757b376070f8354fa375aa159ba2bce67c7422c3e033d9ee9a7c3ed10c7d46bc2614509eec46eaca01215f0bc417e12b56a3f3ed07246032ec3a21be710bd71a2efa31a29fb03b8fe9d789a717e3130bfdba2ae78fd94c9ea8e99a53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3fdda4bd0f69d9ef99c4b2656717aba2fc83c34419e2dbeb81752c8860cb31adcc4311d2e333879caef41f434f8c0a1636608262725f18aff87994dc92319600cbe1a15848e9ea2030f8ab7fd2ca3ab41c6ed28fd1a9f8b5d1de9df0e198b9c02f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e9d775275ac51fc29ba296ad4e73e874e1ccfcafe464fd1c32fa9246a0f7e5f7ef06230fd147cc81197dcc82b81d21125fa46aaac889dcd9a308f111435abdc015dae8d4d1f13371a8207c31b52c176beb31635f6e7316f0e1c817d7e10e7409ff3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce75693e81fb8cb6a4f6eb0704472b2c06ab544d07dc52af8458d65d6413ade58e09ae9d7b3b9a48b1f6f2a1baa2473772b7f332b7f615fd10d025d0525048dcf156590ee63426eb3fdfe5ca5469c2672872825ce5e8e008d2aaa36404fb7c6149c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fcc339eb8174da05e997a85b083f705f6f5325fcf4e20bace41cf2ac3a36a99bb81f108f6d99000f3e06a1d090d83cac6b4b85c87126da4297a1c26f476b8da50d4becb6f09f9f682d4ea0680a5a3f7c13db10ac7465b03f6c61b1122811b62d7f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfacdbb3c1f9b10766005bed70c0f6aee36317147726b7849766751a149721a288c27674f9f62b7161306169c7af5cdf9d8cba3ab70b25c91a1934cfb8e19a6f00f3af7533fc786aaf35aee13d27befbfbb3f8f724fb9d5cf7551c007d2310c48c29a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9405aabaa18a58f6aed4eaa445e9223e379857403f371c405eb107a06b25edbc1b0cff06f1a31b8de4853bcbef0b02a4a7448a73c5d90fca5a64f51313b27589c2b87f14ef4f2fc7ccafe9e6a5fd1afabf1b2cd4645575c95f422cac89b3b2caed63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h589d5c2b72d68adb77d1e1992e9c1fb14c9baf9fc0b5f001b35dc305fb6eff4c6e8d97abb329c6025ade2e854069710bfe36c2b27e8b4a522cfa1b4c4740368a8b3975c555fb908b839ab3cd1561f9a9fa709bf8c1de573be82f6239bd51a20861c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fb6cc12824622d447e4d58b26b52753ba075678cf2bdbb227d0dcd964ccee66abdac9a488f6d3f3d9ab9a0e12b31ee3d287b87ccacde058d92cba1c5612ac7f11fb68318bf6a24e0ecf276d7c631fa5ba90d40cd30a0e8850725a34ba126a190881;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he97ad6f7b596aa48d6a6add4318206690d005d3bf3ed7067e5729dd26ba755367ac639b9a7d5d4810b2cd78708657291b6454ef04910f1b83e664751ab3ddbb3f29126ae00445502318cd47bdfaf7f98fdd590d8ce0a7925b32d76675aafd470d3c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2b70f34d3ae2c97a7bad9d24e67f99b9d577c84d47f0139113df7c87076ea1fb22c8eb87cd8e841235ca3df04cef2dfbd9a2c36232e991ea305e21de27e8b29d13c3e0bfe6e443ab6d7f00bbeb103b90f0919a5b69166e943d08f6bc78a58061458;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1810946268d0a01690544bd0a71efb02a6f806594df93e0de71d32c045abac02bd45c427b2eed5d5955651e011740a78a81da80ef311c0deda8509616d7a6eb7bf1e1e272fd57213ee3c24b7fd8af880be9093328f3fc84b856d007951bd37139f19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he794b8e1b5aa025bd974029db16499b81014b1f136a1f09dc3d887b0f8534a518821d6706f3522936523444e7efc0315894df05ba08fba935411d154c950e53e01123c67b88b5026c6249e8e877aaad6af8eceeb55bf35eebd03dc227655efa2d2be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcca67cfea2785a720fd11adf9a5bbc8a7512d2ce50073c47dd6f8011d5172214ff9b64044984e96db3db1adf7e14214b9f28e74b26c53a5f16c1ecb77df632929bdc08329a5b806b220aea0a94487726a021cb69d43bb2691a753c4d7c1575e3a8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86efd638ee1a2ea3c6bbce38e8568de97ce5c272a75a8aaa0c121b4259ab62fa230ebfbe76b477eccf9bd57be3c8c90f1b3a901558a700b23c76c83c6076455e0d297aeb5fb306c40a38e73de77f6c95add22b31373387a9efeab57349a4bdb7ebd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf801d934c4856f05d034bf25fb4cd34d87c9c0ee45b0c24bd4144cf4751e1a52221eb4b8672c6f2ea9ada1761d2a3d33aa22ae75bb0abddcbefbfc86aad7f20d04432cd7ce776ecbba4ec55bca1683bea4444c2d0e2f3c7f0eb7da3161950c526394;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd869419f417ee48f42936ab66fd922d331fc4990cb8cf4d415d53c044382a180fef04e3baf571802569106c05ae2a50b28997331cbff645978964300efaec1c73488866639c90f000db117d9d74d1118e56f6e4b6b4e40ba6ac83f681ec9def80836;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h201f2b91bec7d35e267c8c4cce37864ef87c18576e79bb1046314abfd22da26af7bbedf2eec6c5f0d47dbbefbcce13278ca20d6fceb1a64de8a5792f6a1da279b7bf5a834bbc32fd41081ed6ba2efa7d19a146ca313088d10a018c70a2621b538c4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb77b370d33289e787720781d402e273dd5b1cf26530e6cf6acfa69e70005e946a11165cd4fa52abb7812c50a87b8ef1a0ed2952d2837078424746a1db5abb9be69d5d3ff869d301e14c9a52e314d5f99cb24e273d17b3648c6aa7ad53ea707a2585d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15a466117687d17e748719dd3937520cd85efd85e6d75cf5add0b72bdccb6f2d8ebdc9128cec0bc9deaaf961d14cbeb965b89bf744c6ec9d091d48479f6be1ddf01e5e30f6590aa92cba184d835bdb37a4d37183e7a06217972667f76cbe96398e73;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98f66331d2b8e3f86112da8cefe659782a4f9e67d76e5cb67e03eb9f53c938b7c70e3662f912e86b36e63fd41edd13a3c3c59ab0c4ed108ccbb479891b05e9c83479ad0434d6e579f871618c7def4b9d4fab6533daf8f22d322083a6124ed677d2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78abb2fd35f91c81f57e5061f0a9e2755afd2177e98ac86d2bbcc54b6b5a4662ecb1b16c2d36db4ba21b2ebe901105a20eab361fdf5ea7ef274ba1d783d39a3e7e600a61d8951a6705e5a0d5096985d67cd455ab42a602d0ee2f828e5096c5862ccd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf11cb75116b9ae395809f87794057193d78901713c0cab11c3291281cf65a8685da8cb7450e1c869aebe1f8ae52efea57f62e6d013d7049684b23537cc95d956405b2eda1c3b0a54ec9d827356c71635258362055bf207375d2e6920b4ff5ead0ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb34d308109ba4dc8caaf196ed19b84216b47e39f7631fa6789086f2a577d022d30ca099410618e5e8bebbe614afa6ccbff0b03f6fbe22c42824de584092f0a1cddc9ac863cf605799b46b7e21dbc45ffb305467a302b73e4089a1d9b1cc367816da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb97d76de3e22d4985994398bcc064abf37c9a6ddf8b75b12f8f37be51f5e9c23509bdce467ef3ce740756003474c86a1b0d665fe58f933e99dccc125258b824e72788fdde91d844c5be5ec3aa50f11237b931bad8bc541d56eb53c5f9ad48315f08;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d27216180bf4cdfa9953b596765f8a13cef14a886d20dc78ebe551213eedd10454bf079cf102e220bdc442471de4eb7350395a87908bb887aa9b4ac354b3c35058198e61a60aec08e4f2b29d03984ff8e622e9732816403dbcd56b94c207ca1f564;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b4927d6bb467c826fe42eae051d531633e6e5d912251b847aa72a82fe916cb552f84f1ba83eb2ed9bb343e6e92139a1519b908667cd9b9eec3944c2c98b4b329bd25797685676624aef638815494a56e73dc0a232595e606b2bd562dd495f80d675;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d3599d836fb3cf3e8c39122997a6ef94413f0766619ea85ac9c940e3c94de2e8ccc8d967c1659f70f2aa42536aad2e4eca1932c19881d8c557313d8af53d6fc7257083d3ae3c7b830ebf1f87da1b459d6f6ce9407686fd33f892859dc2a57ce1c6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29e44165dd694229f30806b3921ec9b583caa2a24c7092e91341db3c4b82efe41dab614ae8348eab0521f5faa8b37609df2bcc38dc7760c967a333750662af6c6579eb9b6a70b57958bc0eba7f9ab94b08755888540a2b77b6cee208b475d59a7dcc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ce865b9fbe0c1f5559a85b83a5b651a0870f1aee68fcb489b98e8904fd103aa02307ba5894fa45900737f46512f53ac98bb2dda4c8bf072d03131b5d519130f337050fd34a2826235dba0b892c5b776d4bb3e8fa7711bc3d5bd196c1ca0b261e9e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2deb0a2a9ce667141f510139eab9c92db81deb19d07fa8fdac53a8d354bb4a285c2dcce8394ef615e03e594a39b1b030ad1e35b1241b2ed33729a55aa918541cee7d00834ec8dba2d19240f22fe4990f37048cadfbc07846cf11c268568e1479d537;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29ac68a7759c042752600365a6a4e1f52a625b245c06bce0640bef6d46a5f1f4d58b4efd874fb8f1b5e130988ebd8a70f5fd55aef8920e726166372e4cb5d77e98beb6e4137e129e862e63e1cf5829066a7883c6c8b88660f22a4ccba127d57996c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a3c564fb74e2e1d6692b3f486a26af2d891d6bc4c9bafc02bbf51cd8ea6172dee3b53a7d0b4d62dd729991e99f74708ab64b926d38121299bffb4cd7ed6d46d37060baf85a8aa0f173fa916e2f9b75e9a0d9e40cb53e8b7b2b9d8cccf835cd96098;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h702048a6cc358a07f68316690610f426020b99a71e9e21cba2487d6c789894694ea73a42e7c4745bf1cfc59521a94bbae00721d789b8030d4976f8527454cefd3e7006902926d501aa385ebbd85db965d41d229b636e6b6f0647a7f4a7720b7cfcac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2d2b52c3aee99b6e533583b52bc1705b1be56b4d526483b41967cf29d28cac0da28c5ff0036669c6751e38195e3f3e800ed373a38ef49ca17cf155370077d9af872f608ff1cbd00fe157106944e78f21b40aec42f8396509ca6d9e0251f3f4aa811;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h439616833233a4d5651b7ca7bcdbdfb2a8023fd0a7b4909a86bb8cf97371ed14ed12e31dd12311bf8a60b2a5f7277b7505342f2c78729cb69b41efcd5d3e636cb50b2666acd067eda37e1d3c5b078891ca9fb0417844f0f4d38aad60a9245f263879;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8ddd5dd5db6e33fddf15b223e589b45b0001bd5e186acad1c0277178db84f3651fee94bf614f3d5655ed7a3df2fe81b91f23dafd73ebb4780995e36ff009347bd3cc0258da9c2d29d7a0cc187d55fa1f4a1328abbb4422f2fe52103ee7f0efb6245;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h648543e0aa8ec1e60e208d2d971589ffc4ae6c1c16cee053b7abc490da85de7eaca3e74d68184e60f0775800e440a29fdba8cb5133393db5fb23ed486940552d3a0b0172115540473893543c8bee32d25a196a61105d7e37635fd976d5ca9685d8f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heab3584d8b9fcfbc0521a508b29368a536fd420b94e53d5aea66da98f0d818d1389b57f0b86bb24f836c7495b6bc986a28fbc69e12d09346318693c8c28d4cb537c3904e8741743d913782231e49fc4de17a5a6708ede546a41b8ebaae3d94d3bce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b8375e7d01ea287a24ec43dc9745c2a33a61cb1b49d8bc65e0fb40c6e27e16a16c8e509190c541828c82e6d06d207df5578d8e38e19e9bd0e32334a7dc4f6306c05d79a1870a77ee295fe6affa62d228fe6e8e692dd3a9cdcceff8074e20d8b0f82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37e01d4e38e7d7e068bfec8282a665e18fe9a80138a1c0ab8129345b6e6519205355c595a9646c3cffbcf4013eb56be593168654de291558f929e9671d5f21fc3172cf2fb95da59634d629d59d24dc895941040e8593c1ba3f074dd910bcc0f74734;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3ac1983fe35af98327fd494e91bae52b2441ccce7a4e3930723a5204e14bbf18f741ca1cfc9711898c86a9c39569f4455cbdf65be6b1bad52fe3c4bdad5ae2380b948bc308d3f7ea66518f5f4dfc98fddec647726f6e7bbbdca89279557abe2b9e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2434e422b00857742f906cbc7039b287698fb9bb4662d795a08388d40c4d69d5a6b6f2b03c196d924b7f2dcca5e6e39ae77f94d6be1497195dd7f0e81fb580602a39b9ab025832ac18c6fd9ba1d9819d664ac9451f7fab12a5482389ed000d48dc5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ac7cf7405cb9da13da2495f4bbda513051835ddf06dd8bcc7c75e9e138abc8ae265123ece58dcbd0fd9dc5b709672110f39c05c40e053ad6886a02b8cb9ae5e3d9dff13ad417780f587548ad1ed6297a4c744faee2711b2bb91a1c387f7bac9577a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18f091300e604e8f2c867ec283d28fca5bb1258ba43841c5922c3b77cf7d91b985b0b88cc05535fd85c2b68163f959caba813e4a3b09df2875b32444db72f1a3fadf1b28bbc90cb07c3b75f7bb3a655b8a3bbe78e74c3f1bca331c4cebe8002fed8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29dfe1d16e48e27657e3504e86d1021cdc42219d5ab6cde5976b78f68437bb3c733f0c4f04c2cacac28c37ae89c04ae0e061b35805eda2c8260078141fabb1801c01b5de91248a1f621682af24d2e3822cb2e01d045b9e3b5a612fb3f57c572339e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ab213c52bc75bc2d650b9814c589c22824b556c7b0419e3bed610f363feea4f51f6c0d7117ab23d75dddadd513d39b8458df31fe640485cfdccca05b938f7540cd35c99f88579a1afd05dce6db0af0a899a74668d161a3157c24e4d00a9c37931bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3bc053111956c6e73febcf41bde0af8304b850cb178a286763a670984928d09142c2c41492bad38da479c4363b57f25e491b65418ef1607d0e489809835ea7c39c61f663c4c359fd1e0f803abae0c6eb763215ad9daca6ea841b2605779e27ffa2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5dc7c7b1f038c8bee2464ad510588cd887d2b01112b1cb2f0d04303be334c8cc46cce1d0b23a073777d5e18fca1ad4094847ad4468aaf2f29406a87476c48b3457a9b60fe061b7f6164ca5b5a7c3264a16207e03056d0a427731674fe5a79180856;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h277a5a3e8ad1ae60126b3bfbc85cda45e374bcf17c8010ef6b492e761de9bba92e71923e644eaf8e9d444f66875d22983fddf4713271f561e53f1d58cc6b0d39d0417422eee2ab81fad84412a0ae672d077f669433052796bf093d4280b2a8388fd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4acfcc2de8e91d67d9c2895d79c93a40f6bd8e26b5476460c519b5adedbaea3bf7271e796581b304e3a516d862a985c082aa741a1e4f2cf9acd9b8a20a2f389742017d7b2d4a5b45d5479e627d075a1d72fc78ca0b2523491a591ddd0073efcb290a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d99398e428236dacd2d5c82ad660417461cf7a968aa974caa66e8b3070b0b0c968c360a0db7062d06198d42f85aa984d28a9febd197cfbbb5c27785faf0e6bc237874dba3a95105b9dd479df498117acb8f1273da3946fd92a55cdd3f411b700d98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f9e43d4c0c955cfa6a615df530c51a435fcdd906b287b4faab2f900d13ea33831a579f5103c90b218c710210bc10f7b130a917d8cacde0012842f52ca4b75278d2415957c2d9344bb855dfa1535fafa10c3a71d3a1a88398897435eb28acb062dab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf43e880349d6602e92b8d8b6de578ff228c23c9c9ba53afe68406f1f8ec2e94d76d29ca0a51a0544828e01a0e2885d63815f26d9d8994ccaa5b7998cb25d70ae42bdcea74a43adb01c017046a96ebf8b37bd3858c7c35a189dbaa30a29257fc26712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3f8baf4fec82a0b9f12b159a982c9e7ed916122b8fd11497453318ca9856af71ff750b00a299189759e7ea0f04f0787df97f2226bddb908bcef76ad5b628f40b3e8d3b34b8a3fae15168cd3b38584a4a41781c56f56da80ee0b0884a92794f8545;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d19b336f091cdaae56147cfaff603e32007cbe5ebe5d9b29d835d4e31d906a123400dbe2cb0b6ee8bea8e3f365ae8c96039b90e2cd44179a161cc69278c4e47637478b91d65cad3dc64ffee2badfd065960759344f44c9e27f1c06bc8f40ec24a54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11a3d7d05adfe0a53115283d8c58402eec3ab8dc7c55374ee390a893f3c36a0706f428b0c6842448007dc1cf79e787d729917c5c0dcdba1e1692565655174634adf4336952440086a2169a9c5f22716ad756f94bb1aedd2f6d0ddf934fd0257954b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h716a6552c8732b895d579301e8514f594f112d9ed7c6404261da618aef2768bec897714732bdcce008187cd5a3d69870a4ba1a7d485b58c54b9ce9510cb0880be1eff68758e0422c0f676f12e04de3f371cc415f2609aa4d52165c363a95b1f60edf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9d394067fe87aade3b208d7b9f1d53b43854be1df294cac98dbbfcbdc46e37e73f05db9965d170b4db0b582b3fc466a03044e14deebdeebd6a7e3a5f40de24acdc125b660605c05f3bcc09f838e20a78603720e6698c73253da282026ebb7a103bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a01989dcafe595f3517a89d48ed75760706a82fd4bc59a32fe87c1a302d03f66bfa476c800001e2d02a295af33fc1a756eebad317bec4ba0bfdc55e56d147cc7945f14622739020b2f068f895e3bb5458e79a0de1ec5c3511c484592e87b923a3d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44d496edb32d03c4fb6c2bd57382c0dec0aa4b0ba5a2cc2215cbb09a0e6d093d8b87866af07b18190ea758e2d5906c5bdc7e6e2ec3eb4390ea8355a324d07226a3072134adbc934fd97fc8712994b6d8ba43c54522f428a7d7c56179eed40d776b4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h569349649321b158ed5f72980120b8da1f793edaba1329e4ce04d09e2bb192232a560cc6582d15eee0118c5d4e57c8ebbc80e45484d8f5c639ff3e43055e388d57ba4d616d7423375be02244c3e0803c25b9d3c8e6ffa5fea69405ae8c931631e97c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h120be367e5c4149fb4f638d22e8efa8c81eb0bc29a93c2ecfd7e43b27204a64b2a4d423e35565915ea1503d8d44e71de69e447bfa449050b3dd1655c08e4e576ad40f6bac80f34c226ad6e5ce1c12861b52cbe59b9f88f30bbc8e3da5bae3015cbf9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h221224dd6209f0b042e3ddd79e217d4a814ccde384723d0d79dc62dfcb0ad4d00b9060131cc5e41f728ab0d4fae82eec0390e65ec3aeb4ed0e0891bbda46cb0a35f08f466d17f75cebd3c1084e0245d11411f5e3e47bafac16809afe8d808df5c15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac6a3d387c7d8621cf3922a7c53a8e19aee3efbbca2f6f18c10d59ae6969159666a3ab52079bf6a3d7a49b1bae929f173cd847815b7c4dea1ba329abadfe4f9b477f8ce0ba276e1e0a62909df71c0b74fd97ad6f82f1d062b059e9cc30a52f4c00df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c67173018b74e14bed7de9e3d8496291c79322cf6f1579a81afacc3a825c9809abdd5f68fbb88aa52bd0be29664b43c92ac333b559da6d9f91625762e9a622c2e7d0c812ab60dc9a3922f0a25fb60d78115ee2339f618b8b094a0dbddf55d34525a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf1459376d0f7f6fc0003fc7770e26787bdf0096cd4e16787e2b2cf4d76cf8d6a847b692238eb08d98efea4a0923bf794184e69f0e7bc80ec3adf72af486049b11633e1e8f30c51fc3150ff545c52af08901ac60f11ae759cd86f0ac6b9a9f9eac2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f9253171a6e9898dd49d1b3e829beea3ea43c748a1c91197c6547fa577d1220ee92572d23eb63b89120d8617ae9059306dd86b34a38aeccb492dc16c1d99bfa8a9d40e19143ba658e970aef3ea1569a2fb940e1a7b6ec5c5ee630f46a99807467a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd262879b526214109b43f1b642ebf978719eaa42f26be06af19045d0d1db8842d77e58c74ba49867fce82e830cdd59557324f7481d4504212d496dbe92f72f401c7f8a8cc2a2445e53a0151eab6cc2129b546db0efa096194628e345c98a406d5db9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10bdb418f6517b45a59f3e61f6a165cb8fdf8fd50219d30f0603e6e57d1a93dec5a88c728b212a5852bd526a08dbbfda3b977a59d5a89f8f292f3a174002fd9f65b22c75e4848e694f1cb3f3df4fa9ba69fe1d2393be9e25862876c23b9e5852fb9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13d818aa08a37ac15921ccd5a2d6a8c04a8ebeaca20f700ff53ea8d2d7b641d5155ec31971b2cdcafc7f7695b7331ed1a080a6758d4b78454bc232a8fd4f378e503b297d0a035a90f05cb8035b3973007375a08112513f2ee58bd8646db79a0cb47d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89953fc74eaed1976560f2bba362b53f9ab43c7e14e9c0eedcdf7d1e1ecb95ccea4c428a28ee463c626096f4f26f5beded8e662fed77d886cac805443add8eb7efe183f89438da28f5813e651b68ecb90a0b82a73cdb61f1422e8460d3bee5d7b238;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf326744d7e5961ce14a19c57c5384184bdc3a94e7998fd4ebf71b5896b9e946bf3162823f8aa8bc46d62ff9b0740f4ccf0cfe0e4ee471b5a1bc0fe28a333b497d1b81d6f1550dd5b32c628a3eea3ebc707c8708d643bd5ce19257d0f2928338b6fe4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc750a11f76b76b5685d1a92039f662ab1cadd7eda92a826c48c1e604dcc7b3e4bd1c055f003e1282b82a07e294d4728b7953a486bf6f0f587b37565f86429bc84392f503388d4a7d0fc76c9f19f9314856932c4bb9731f148d98b9737c8d4c7b9d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf909fccfa52525f411edec6c06a4a573aa105b414d01b9b1639a4301daf785f2a25ab3792776134b2de81295b07684ff451f0c1c3c6336aca0ac1db4080e122a01367a83225dd10f7eab8f7b980f3de04a093c97bd85068eebc253c278af7da5b0c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee0aca5d688437c2ad95d946438c4fc2e987d749e9eb5f5f9c51916094f74e5dfc8aaaeb27d480ca0ffc52be853acfe49635541800c42d3f9033a4f67ccd6275b056cc42119bc2fea20a44eae05a96724314e9b17e38aa4953346ac7fbcbc307ffe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90db703f4d743d42167597917ef8f085a38fd52b5c2baa1d3371480b15e16db9408a73c7e68097823f7219bdb77d765ac614baede2281e42a814ab938dad93d6b168a15e323d2fe215266dcc33f88e0c9d00eb5787e9feb5ca9417861d4a35ec3a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77494c87c53c96e2f2aebd8da2e4999bccf5c1220341c4ddf99214265632d1f8774181563fcc36b6b8d773a4157c7fdc1347ecb96d793566a0355bafff03c9303814b46895508fb5db2df78937dbc5ff369c2677370d2dec8408b2b7e54f55beb1c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b96094bcc56360707026fba4a4ff3a7ed22a7c6e8407ef26a5b7afdffb6ec31e80b3f3be78b3944ef14d61bcf095109f2c3eb35121760c7d62c50d760fe85fe562531e3ea7cf3b44f95b9045c783f12cdb50bfc551a3926e06f722ef163427d01d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf81f8f29897040f73ed1ed700dd25e98bcd2a64526b1b7ae313a9fa29b3035e945a2b06d887c96393c186380bdefb6b1a17a6350db6da46fa9d71810a3866e40657bd66215d9c027e5f098d743731d4545d4bd19d3965c9c75f5fa2d4c51e4bddcf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4a050648824b435f3c7c70cae96ac7a50d817e188b8b41417f7fc3b80ccf3147db047c23473b89799d50aec534df7d8a95061ec4e1572a8775247d6f369c8b5ef5712201dd24722d9418af9032b31137ccd38400ddce5447ebb4f29fcd6abb31147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31b0576111ff01118907eda9f82326a41c2848ae8a247cfa2b9d6fdfa18f4e62438d21323c801987f97eb94c1cd4e1f511faba2fd4cd969db8f087931f50f052f5c681a934e47a66c246173cd456a3d83203f8d1f154b9bfc1e47290c439cf021fb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ed2f12f1e4a1149ae62a6ab6a4a93683e703c7617c7f94e97e6044fe4488feccb5bdad93e00de09566838d35efd8b45ea10ab5210e248bfa783de2ed055331e2615befc336740a456f57c2c2568201610da6c03be49ca94c625f30f25e00b4b9a7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98e774a7a1c86ed6c0d2588d8cbc55a2e6f303b03bb8d11cf1c5774e09a333f8d8354d5cfd7a6258e051f5ab12fbaa90e2033a1f0faf3412ef1e61514cc59acdf711715689d5760326f0cbb79a30450a35956cb1a77355fe80636d0e8477e3de14a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3aec3d560976978cda560912a18365e7222821db0ab26a2477ef105d1cd07bd74330a803ac2a1b30a56714efd560971044c4797c81504b9602d8b0b22c9537d178a07a5c302fc71be2b946babc001e05b51329517f694f480a28b5f1873deff12163;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaebde04139637137c72715aa2c91ffa0c904ef753a1b3cee5fc15cd76218ba7405933342cdb7e8175f7f06a368106d61822370cff9182870ed274195ebabb57a562233c5cad5bbf74f747f94ff0aee158ad72f197f69aa5f679a42da37ee07768af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4db2787123d0a8d8e3aaf8d6ce6ba2d475179cadedbaa6a8e449948a66e4f92f6f60230ef1e33ccd629e3a55477e4aeade9e71b403579d60a445d36fe2cead6ece9bca8996265ba81a73f59f08d2a46e5b56276c64883613e78ab04b52596aa013a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11efe0d188553338ab8d84a6fc7f60628d5266236d6824f365d291b43391d3477a6c26f5b6e8907eb1b2f629f9c0cd91d09c3c10725b38512cb693ba11837b5032a34fb3c4dddfb6a95e026e9b8f9a38d62ed1176b645e64b3fcd3a3dcc714379034;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c83f23047b6eaa9c78b56f7d9bca62e1d0102e033a19f8633062a080d2ee073252fb34691f63c53a2ffdac5bff7ae91c93d627de45c942535f75fc82a8c99cdbe3bf359f3dd1a8dd66e02bfbe22d97c094715868cc04ce0eb41ed48c46511d1fe70;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ae72071500a2b5299c237f14274d928b8bbdc4d4bf22ed7d03699899ae29b1e2a0e00df2a83bec53afbc447db7a7ed40a2ba54a849577ebd5f354e325202382c1ed9aca3336bc8c59cafd13572a02d7a75a1fa6af3bd630694d7cda5bfc6083f6a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56b64a5c78de401ab4ed4ca17f939baf1c6044f525d846edcf70b697708bf81ec4ae286deb053a5ef7d98d2b4d5c27252e7d5b6758555642776ec1c8cbe2c315fc2ed9806bd579c472e553d83b8eb42ca57cd03c18f79783fe97200a4ef2f39ddee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c10c52ef53c7f234db73d667ba95006d1140d465c1788440c7fbedd6c61ab930b2a32c2c18051ed30dcec0dcefea24ac78fd2c70a8bd4c793c3840eec76eb770338230ab1883b8c633db079cca32feb6a7c58e4b042568c17d60df68539c02793bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca01128c5296304bf8dda3f562d4d31cb0393d5bde4fa4eeb67a7b523af00c2fef0381a72806f831969b8c9ce429f673dd9dbb109d7788c8c7681dfeb78aafa10c1079cc963fe72e3b41801e08f3b46f1be86ad2f6c3a86f76023e18dd142691d201;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98ddc1673b15c97b965d080b6d9a0bc8184bd81f9741581327c0da9781f2cb9cf0a5d8fb1f24c0ef8a4930582ace179ca04ded070d98cf0e4214e345e5c13d790c3ae3182be9f8f11982409592373428453a34195dabd6e3dc94ba826c44deac9dc6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h196908858e7242ffb7475fe65baf6e49d160bfccaa360808de2835edf97ab003cebace8039f0b0cc7e494b943f21d217036e9e05ca7252d8798675bb227e2758ad11387a21c4f1849e81b79bb786f38354ebfaea4238152206cbdd0bf66ffec40c2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ab9e35592917fef38d3db038cab5a4acd8b5c1ffe2dc62e6abf11086cea85cfe9e3e35f0abe2438c409bc51876be302fad0f828cf77a2e3328647b584d0d310aeff9f9d81f4f90c0a2a2ec7883d29d2ece70e7e767897b2d6780a99b8f73489aa64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94064bd6ed111c92ee31f783dc24b76f5fa8275c9c892e34c7a0acc9ff357e0d2b20e5d586e4a3bfe255c2edc2e4bd6c05ec0688525c30a04298bcbd9632f9695cf8233245db4b29ee0f09516f30c157f0b7b6102c292b7b1159b15b6d1e171890c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcea0121dfd1b3c76e2f78cdb0dd4f440983f08d4b8649a1d2bbe76a3df776adcec116868c629772a0b76bfc973764d772be47ebcb7db69f86240badff4568083c552795b394cea2c814fecaaaa04050d96131a1fd4339588c029cffe3e51b83e39d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h275c2beacf1f7b02a59fbc4f6e25d968f1b6dea46e9c3ad2039a95dd5b54fee2df74f820bb672f800454b0d5654f9b2f81c383210f7dc4226ad9c9576a15aaa1b4c7904610bc6248ae101bf304c0d5614aa44912582ae32f17bfe2454c7a6e9cf057;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15c17a121be6418a5a31e1cb132f11111f5e1ff9bffc1f8ee5534a33ebee8bb1d8b09a593bab628b4c3088b30cc17f7619b2726eff83449f0519d6d928ce35da4c5655a4a45d9eda49890dfc9f01eed68062f02e77b803c78126e463e661f2042298;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb06555099e2cf7e81041b07fd99f704d66de15b693471de076eef7c5dd43fd9471708af50f9c9dcd8e70f4a90afb6ead82eda320a2f973cbb32f9f3481b925b9ee09de9106e6b17487e90e2024cc3ef2a7ccca97658b701561a6277050a99f9c1317;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc09687618f957ce0c40dd63ae53cf55417db086883cb935ef6e75c4950042421794a1e29d0b40d49aaaa4d1f1a98b1929a9e8d1d1e1b6a406a0259bdf0ebf94289b46eb5707346733b159d790d18d8b87ea68526883bcf4112fb17b47266daede0c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd8e5f563f7004d1b5dcacfdb45887bbf46782c78a7ec8bdc5372849a21360a3c523c70db6d0d930cd58d3519960c1f7f366f729e1f3ce54a0078aaadb3ad0abb27f91f131dc768f2cf13327d9c340d10664959e87373f7348e6a29822f286fe7e94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1caca9c974424006f80181434b50545a257432cefd1ee80137f72217f9675ea475faab0d02a25d13b358eb9ea2e9f977d0180ca9af4f2c7ba16a3090a6bb56dac9df15cbbd33bce70963fd69d2afb66fc61d9ddc1595b10d99eafa83954f12e109d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h395e0fe5991e53e4217c9115bc63a311305174e1051890fa658eab57a3019506546218014d83ee7788a02803250f4a8abe186219a1ea1090297aef1710a8e0762c5ffee26d5dfc2f3c65274d874d02778f9a61f132118bd338694682a03dde570fbe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h186697b3046fe907d34d9e7ade2d4404bcc0fc68c595d375c96538851506580a8e996fde4125ae267687dc6caf9f93f56995fb2f94a92508bb7cd4117b4af88dc15051d3096ea97df8622b1d03a515aef98521bac8897f645ae1b0da000d5c774ebc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h122edbbcbde912267b737a0586f04e32debea9a3ec33925d1c7091096211819cc1afe9986f019a844616fe753c147be55df7419cf362ab04ea50b9360129b366e0108de49cd29310f72648a263a295b93005c8f33660ca9baaec6669ebc1a9b85d6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haca627618115759e68e34c8651ad27ad8abc9f6614a77c56501c811b8c447dea8ad206884d519013cce3739b46dac35a5eb246249091acb82355bcb691437106dade5bbc9b2322d8ad3d22ddea8721108bb8445e8deb6c09d2a34f7fe2f2ba0a1e30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b650f14825eb973f9184fcbe9f5d0ea0e943b46d244856f87a9c0cb360e4aad02d452b7624deb926f6710bd9f46d7abb6d20f43126e4832c0b01fb1b9ede7ad4f35017877eae34264ccd7966992155f1effaf4684d8a6dfd4001016d531398a2e5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63615339ab17a8873c3c84ec5dd33714f17580ea8b22bdc1c8202474187867b47793ae8958535abb6c73274c6433966274be90c73a0f744a34da1986e7808656c23fcd35ad1cc833cdb090558ea211509c2819c5551afc815700e841da098f8a7446;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68e1f37b9fabf3b66f36aeac0527cbd75feeaab40edff3f93a9e0c5f0c09601c2e7835b085296b95b7e4cfe8840b6d9f3436d3137b15616b72bc99a9e22855484caf5410d8ee1ee627723cbb6d4644d39c1c5dab073d7cd4dd71322dc1ff33d0c45b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aa9b29f12bc21d9347b6652fca5a04a8160aef1dd95a633026fd132b19b893539eb49e5767e26460d062d8f8beba0e0be84c672513130fc17dae19f1c715b879d3a912f7e827a582da3f6d5541170a3780df3753cbbd2c6cc6d56902c7243b7d23b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h487baec93ba269854abaa98656e54eaa8782a37ae1be4d2e4d0b42bbc158e4f112ff6a2e764cbf8ef2017ad10323fcb084be12bc44bc6c75ccfc2c3b5b893663853a38ab98c64651ae585afdb3706937cd8ea942fe90758433d5ffcd838175a19181;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d1ca0fdd651d0c4c04de77eb09daf2746e389474c421dfc0a0b8d08ff41f7c8ad7c5a5b58b948f4fed931e7382abd09979a67bcf563d1ffb858a75eb59b3a4556d31490474f4b028383c1547aff0089eb0e22b1287b74c8c3a646805c8eebb79130;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcba17accfa46a7be4f7155bf5af0022a73efadbea1e5204099ee5be1c36c316cb56464399bc3111b845098a31b36979018c001a2cdf546f6a14b6965475bca68cf28b66b3ef1c49614905d867a530e7ac6a4d435a4dd52a9d636711bb9d7fe014089;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd382d64617ea529a37065430fe0e29d716abc55e5edc68348274c49919d2ef1d2a74807f685af60f9eb32f931d5f0511a6cacc55f2a1d2a28625544b0b31283fa75342f6dd68d6037f59630d0a8b6fd9b50b5a9a51328e719ca57600c3adcf4d7ea6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ab3fd15fff5985bb9f8d08a8db84d6c7a23d7ffe04beb2b438bd5843ebe8774b72c4c0a50946848c33670b4a9f423636674d6c1e8fe07a06ba10996fe01df5eb32b87e6ab08aa716d0031133849662c04e6a9ae15ae39047ed06c3d023d2249a4c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25d97d99c668f1742448335815d66f4455788e8931d94c4aa71b3b6e44e6bbb8ebd7c71b381b5c979747f2a383875e2b049811d0603e41faedc4b610ee4c58819caf0308f5f322a10b6e7ca0d46bc1dd3afbfd016347f88d3dd7bc73fbf8e65b6377;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a233d83dca697b390e6001bd36d5c5a7a8a13a03b34eeefc63a255f331c7012c7ed087e542ed3b81f85dfd4dc9f099ea055386b89568f83b3a0dc90bcf71fc28ba829cd92e760dc874013a407fc6c80a5eda928ad1e9762973cb504f4b3fae5b029;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2747fca3494e1b00c9f5cbea66ded9cd1f1393223a0f7d15e3054db8baa9994fa464eb67f4ae9529bec3fdb8921ee858ace5f7d9ecdfb39754bfc0c2cdfe9ca67060625944ccf1c5b43c37db6f9c96077c6ab2579f92c211c8f07f34c26d4553eab7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb73aac3d5d67b925749662be3edf7567f18ad384d73345d6af4e7027907d8a70ecf36f4be4c35d54d9c792499c6d5f0e11f59002abf3d8312856cac3073a1f5f7bd88f2abc5998e992be14778ab8e3a52f99bed62310aacadb2f0098333e3b0de776;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91cb0afcc83430947edd954ed000c23e29bb4ee3abcf3de4a1531b0611e91a55238bfeaafab48f0474bdb860460a032246ea6100eba7baa288cdedd80020f1af3cedd4a5d6ac73118baa1c40af4d7c3e4f752b2d89149375b18bf15cc715943cf232;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0a4bdd805ff115a2fc8a4d5a4bdc15de041ceb6ffb1c0a30f623104da03941da71f4d1c6cd7338bcd75e2a8592407f7a6da5b87368948e857ea9bc6b310e60dcf9932658e8328f38a156798fba7c25c78044a0ca02443af672ed4dfdfe073730f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he14813673fef81ee5907141f985ef09554c68ca488bcef73adc74acc2eac81f9ba36b12607f63ff039b0c426b7cc2ef07a43ac075382d3c01df56439065c8935648775ff38faafc912030bfd7bad330ad3ba7eb730bfe5d8f0f5c792513c868f1cb5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he374be1fa25e29a54e1aedbbcf024aa121018eb577d014d8a0b7d345098681f638390c8666bf496fe7285e5fc4ca7bd603530bce925a8104e2849b8c6ac05ab0e382077dbe4c86c22f20aff6e059094d0a9b52e204ab13f0fa3ca802c9becfe4b385;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he07bf41a170a5eba35d998075b3bcbda545a60d06f079fe0d066fd3c1e022b4af75131d06434d8f03cef7d61731acf004716b18e421fe1fceea5575d643ef019fca12ee4e5fe760492ef929bc3b2ae59e73a19fdd8c5852478a155421ebc79eb8de8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cfdc3f65958927a67dac43bd4174e6fc8c6b4802c3748028f20f8bdc61dea7498b3ee182641157cb40701e75083ea0f3c80178a46cff93f5b98f64700ac4d3f4e225c580ab61e5157f953ae97f5c950b08e1aed2e3648a12537c17c770dd971f1fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d7a02ec2f25eb8b66c9195958a34b728e2e4276216505e85de6390dd550ab291270c52fa81ab987888bb69b673e9d2bdb1a3aedb417c3cb3c7074434d75120a452984728a570f523224bb69be4a9a52ce67901ad179111d240383502bce65bce2bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25c3b7ad4e1e18f89a26cf0bfec72a376e6cc5d2d7db81b0d2fa278ed638d990ef8747187601dccf7947488163e847bb5ca2974ffc455a28cc40ccbf4c6c0b777936a4a32ff1feb21a6d7d45508570333545fca2f7a5834325336d36822f75e511c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda42afda810b88a357b1b753abbc40192a84a331f49ba272dc72a87376a640d45605715533eae8128fe2182c3ea3876b9547a414b1ca487b33daa2d880e9591977b1c89d39ed3c258696655b05ee3ef0a25a3a1cf77b3364fbf179ea847219824f4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heca35a94bb77fe5fea9b4bac5f870cb9c59105d6046fc05e40ef56f4f7f90d703acf75654b62c9ffada8b3b92d45161be2d157d2577bab3d94fec266302d51101fb0c519489928777dab5d975e4ef5ed0575c18dbdd213e1f3726a4fd0ab46d91688;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5bd1eeb14877e75e203a1f42baec3b3c2bfdcf837dc669153317f772d4de99387e3c0527578003c6fe523950fb34b9058c3ed71fbdc2143071455b4b1953309c81b8376973181fd6f13683192efe27efa41124f29803ad5c258d32f9ce21dbe053;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b50a63983003610dd6c9fd67064f9add85f4870846a4c34059e318400b5fdbadc4180500a49cf17f72cb352300a2592bb6aba623d178e31d1613f55fe5ac7d92a812fe069128be4c50ac589bf8bf93775cac9312384d3f7e0d3b46ff063ca4c297e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c686e85c671e204f01c59ef069b532b62afdf9dcebb30c42c2f94d7bc60a3fcab7a27ff030344248e809764959b84f2f887999d5b540f952d7eb97a7e2bb2988a88239775179c1d68f774c87a92b96e87ae751e170664a0811c8618e4160da935d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3ab42f41641085c585682f3eeb74b25420d15747cbb7c4ee19d8db09f42547364e08abaae3d9d7d1aeb64f4496442b1d0c4991a2fe1b6c4a5434f56293fd93f86b683e01aa806271627973448e08152ec521e1db610a69386834b70c742138eefa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6be99dc454f28daf381cd28c0a20e7a980ae820e3de0ed5dde81f9af30d144f25a8ffef42ee1898407e2d9549a7aeabc3a743d973080264c782e83deaae0a378de4cdc4849ee12d2c6dc8380821d3d43cd6079a6a8eec70ee3da0e4e53bcfb064cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb140c56dfaab8fd6e28f470eecaae789f7b4c2b09b08132875ec4e03896337c7d56fe4e6ec5901d6fae0567cd904178aca2b1d68ce6c65d472067d82769f37c5f07142b3b7c5721fefaa1c14da14228605948bde8060f8ab9a8d72b69f6b5ec36f84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f8b611700e37e7d6ee6eb3711e34a5ae557d6d7626541607d844ddd0f4dfb70656fad368242adc5fe2654219b9e6c34dd53a051cc6370d99d39c0f8038dcbe860e25c24ca47391d36346b7ae0d9afe8737e371a3f5c8431d07c84f691144c31fe62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c9877a5c34f9e0bbf9bfae78da6e10336305f9c0d1acd5425e989ade452b7490aa41d5bcffeb95a9074e214a00105bbf0d7326ea8ae7900687c39901dee252419feebd664d59406cab62e459cc6ef8a84871fc5aec64aeda650c731a6dbc10cebcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17437eb4e73767bcfb52237614a69c840a46ca3d4269f0ff740d95b5494bcc237b7fe7b9c14e046793f9cd6d9683d90402fb9561d3f4c208e64271f702d1a4a038d72a5933eca664c07885435aa0700ca1f2e5164b8e48c3f3284c61d5ce9d1fd191;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8159939cadfb3f7cd787c9f56a54c3500d8940afa835b795c20b24cefc739b253a98afc66789c99ea9c5b8391cabe858c96f1ef5251a27fee7c0cc0a89d8ea14c84fd3d85464e05ded69bd395a6f7445d7ef1fd6d67dc7917caf936f16abd81539;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12bc6175cd10ebee205f9cf54ef645c48b47aa3fdd43f36ee3c270278644fcd2369be64e374e3d3277d9f2872409934ecb222c6d5e28185311e47a8d79fa8ea9076485db35af9d3a32233f817dac16bab24f1b8ef3ca83a8c3abf0f611ad83a2441a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1d0081d3e72a652449ca57d176dd267cd1ffa67c21264d2b044198244b50ed4d5bd06c227dc2d3137cafd7f265702fcdf361956fa6dbb652c335082588c6855cceeaaf471561ca7110a90ff7e971844f1d1f3f6474cd5602e6ffe9faa9ff78b5975;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e8b8589011e4578b1664466c31dd552a202b1b69c45b2ca9457913d44d6d111c4b87997fcea7cb7b6c210a13d5fb51cdbee82ed1dc76d5f0868b0d6b2c3f08274a9afeb1a919edfdcaebc9a8596324d07470761729fd7130d469654e7bc396aa88a;
        #1
        $finish();
    end
endmodule
