module testbench();
    reg [29:0] src0;
    reg [29:0] src1;
    reg [29:0] src2;
    reg [29:0] src3;
    reg [29:0] src4;
    reg [29:0] src5;
    reg [29:0] src6;
    reg [29:0] src7;
    reg [29:0] src8;
    reg [29:0] src9;
    reg [29:0] src10;
    reg [29:0] src11;
    reg [29:0] src12;
    reg [29:0] src13;
    reg [29:0] src14;
    reg [29:0] src15;
    reg [29:0] src16;
    reg [29:0] src17;
    reg [29:0] src18;
    reg [29:0] src19;
    reg [29:0] src20;
    reg [29:0] src21;
    reg [29:0] src22;
    reg [29:0] src23;
    reg [29:0] src24;
    reg [29:0] src25;
    reg [29:0] src26;
    reg [29:0] src27;
    reg [29:0] src28;
    reg [29:0] src29;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [34:0] srcsum;
    wire [34:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h882ddd8a1d3fba99e53e979eb5ddd80fcfd6aa10dd9044e4a84e435499068392a0fc52a61927672c7e96752c95c5f71c4ada72642b38f602dc10d5c34b9c88d1e5fac42591062a3972a3956c791ce34a45eafe4fd1b71ae4060aaf374064eb4936396eb1568ae9cddde0fc076e101c6cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cd867f299b2fcaf058392c03930df2be3b3505409fb4dadea8da3923a183a9286ba437b19235a59454545ea6b7a6958161595daecb93471ddcfb05ae510b4037b105b44cec2d1f9e6148c4c51ce8799dbbb2b8b210cb3f2ea93f0fc2ed4cfc5ad6316f8a8fb9f01b2c4f6ba3839d2625;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88f079bfd343d06a537794754f65cecedae03608f2fe73933d31a45b8cce4116f802631048ac59df63c8672f81ef0ca7da8334dbf96caa87585d5d5024c8051f8af29a22a74fbae69f5715734b16528ce6961c530bc94db00198251f691eb0e93d20ab7ee59eebf4d80bfb41c65b62383;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0656b84b2ae6c740e4e121d55886bfd2d7176c1d2b9c8b5fdb7b8716c0cdafb3773fce3398b32dd19634c26289d0e4f7c1ac55b01bd5a2b7b01dc66efdf6430f0c8bce3f00838143df883feebb093df0061fd00ed519afb20d7957d9097b74482810b9c8dd598590d71663b3b6f6085e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3c37803beed517318e55b653c3f1010e41d09ba279a0c5517fce7de5e0bcdcbc1290d5da25ca35074e68dc355b1f40ffcbd754b560a4d89c278c8d4eab819d9dab3efc8af6dacf86b240bf5968619a64b8bb9c0b4bf9aa527843de0a7c79b99a46df722b83e7e5b87beb433321da301;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4b92e5d7b16c7369821661f24b67140e523c01bfd41a809125db73939c0f88bbaba9f571043a01e5fae1e3dde86e7e9aba65380a7d47761475b94bf79c169b295e907c5e1fb46804cebed8a149c83b3177d52bbfa99ea1cb02ecb5d008e28ac98b57d85549138b7906a73851645d1c43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h178d68d4d7cd661f2027139f8ab851cb823fc2349bd8e3f4a4e2e7ba4471509d2c0298dd1a51593877a587960aae1b198ef6274ec7c6e7392e84354eee63d3d8918ffd248a70d85551a5de725b7ff428d66e7f8a24adc9e7be7bc52d7027fb904fea4c3dd6f48e1bacaf6687651eaf0d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h787418dbaff741e30217670a089fa09c5be2f4fee25adffe0531524b4d5b294103f25a98b5d880a60a0ebb10d407f3e2a97e8c6b9c3028c45f68388fe8979082b7047611500b6596cb758325515aae19a7257561bb3550debef1f6d018018790b31ffc208435f5dfd3976e44b2bec7b6a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32c40bd1bf68b9ab0b03845a7a086db001c0d4f4fb6059468ecbb858f5e73aeaab78247246e877b7e028942bb57839d2a13fcad0c7d876997c82e9b4bc62f1e075760a2057b13b738c7cdf70eb26fcc6854b6763dc2d4955937deb7a0562173007bee39038e4bb8be27cc50391dedcddf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed01e3dd2b9d80483daeba0df56299ecaa56e3a9e8ca19f939d1587db8788512c4a916ba6dd148c7ee7c025db920a7c20bbcff6a8ac8e3b0e52a1b52f0822939faf56d6d038868c6c1d99df1a00491fef24041ff3248374f88876e3a49cb61cecabdbe66ce8aeeb291d6deb607a6aacf8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42498f5bd7aff27db08bf916b6f571cb509543072fe67b600b44053f4478fb67f09828a592ae98ff229699c8d681de96ebbd37095dd473c57516cd5ffd60a2431d32526df447457fb267ac6075f4b1937d8331de3a160780d548bb805de1de37c5961c669d2d975f07640e940ae05026c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e351b9be23d6bb6d766768a46a2bb779053b4fdf2e8028103aee61e1737f610c677b191bb4e1ed33bcc57abdd8d43a9011449881d17ecb2e943fd1f85e9dcb324c7115ee7e7db91b456379f3ec2d53f26e3a5162773e32f2588b2392aa3e240112fd0fa193d676f8143203ea35a55deb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d9a3fe42ce010563439e03791cced615ce69cfc51c59979f6a97a76a7b5bd8bbc8e1228fccfec79b335191196c72fbcfbbe9c517dc7f0842b27160afda9c365ea9b2295541289a1b9bee7a0ab6ec2834d6438b5f565ed2c47cb6976d0e50b291a3a9316e01131a85fc77cfb5df9e6025;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a7ca71b10c258acb1c91d56112d91db6d12e3046df23d9fa254be4891158c8ef4f8d449dfd96658cee5730e15fbfd4699bfa6da1f87ead2dc1c6470ac0906e57146e187c66f3cc54c520628b4568f33f3e43f1e84dd8030a52d23065eb5a8221c46b987e6dc1b044a72023791c392f86;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf63c8bd99941366e8b8bc9425e96d02d935824a8818b4b0562587baffa343cf6b86f09a77eb50975458765aa35c76f0116ae3f9d5d98c75b4ad2e44df463be8d3b85286596fa991d609dabb2db78f4259bfc51dab8f46da908f45e7bae97ee2dee7e13737267fb314309f6a156555b4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfdf0794eb14cb51139e5292a504fb01a6ca2d196920feafbb8d2bc840e2b2950b11f8dd8e3bf7d73b7de225d46958ed85a3f18b61848405d93b993af7ebff99d124862c9e762fa0b31fd7256c9b61a97922400c91cae0d4695cc033b2575daf999251e28b03e439a6f1b6778ec5b3fb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5dacf10f800f5d63a3598f855e6e04dd0301f847f2b6d59c0d85e517ad8ee2df39c37b9813a6ebf0274d6820eaae279622917bca39cb49e5bc4e793660b015ff8c4eaff4acfda1da9333e49b73367edf8b854dbf157660b3726fd2a25b7232e5df63cd5e1190af6f6f60c7f402e90e97e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h434b3576857cb5d6c8d6e7b1c16b1606d6260efd8af071888bdb69fe2e7311745d7d309159ddbeb6de36c5cbf76d41ea564dab5d2eca4832471d5adb7ccd73c3ba266dde09c1fb4ec0aec161f61508ec2e4fceb57e8cd1eee062c2c33baf7994a2ace6de7f1231b688be79588e7446dae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceddb695f5a83d1fca87d6770455742b69d27a64d015ae4e3adec918a9718d5f070458ff226a74ca7094173faf5093ec387cd912f57ba5eb10bce26b563f8f69a7adccc17caa699590db9543631ace24d23131bf9239e7851c4664549692af61b199e9594aa352ab436f4db7f672ebae9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc9d3cdd3d8c560a44e5f9fe0d89b7b02fbe21f06f2b9f184f2bb5fa457ade018dd2ac251b3d0707145323ca7f87deefb7f6a4da8b755221ebce78f3e26338129a736078d4676c776aa38c24cdbc2f23e0998b5cb1cd7f1fe95d440bd3804c3104427e02f5893b814bc404e6960ca7cfd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ffb3a17ab698998fa7a3e97e4b61c52ad784bbc811785f60bf43e5a12198878b488e45da72fbb201135497c113346be6b699d9d47f1adcc2bf1ba3ac36bfc16ec334cd1555e3d3a4207b92bc907f49ce07ad6f5ad9b676b16621fd6017eb9e88a112397e2b3ec7a4c7b9af5304c762f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b029c2642c20f0a4d02db44d161e77e9a18decfbbbe653da857101f2ef12675cff7d0a2edf904860a0c94e4d6e80aa537c0f7d4909a029c7b0210ec7531019b27b619d4aee9fa913c6d77507ff70771eb36c474b0eee213d13d0848d8980289c9166d0d070a3c9f942757493f5f4457c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a2c68607eff189f0f39ae50a0d6016ff20216cb129d6aa01c37e78cf79b07bb7f6b3ee962d391b195d7aa0c4924a775926e5074cc52256a785e247f58fa50e901c8fcf5165fccb476512b16772356d3a70e55be5e18049c5c73e100692f4b03c3bd50096fa48ff2114f17478dcc6cf90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa97889118915beedfdd5c6c3c478044d69bb72944f1791b3efc1d4660fd0dccf093630921643855869d4c57c151a0b8d28632c3b1be4609af8f5e6b00325578ccfac9264351daa152ec6cd40f108faa5c35ee38c0036e1a5d069dca9b02fc977853074e0c25467f66094c7278364499e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bd0ac7ce6e2d980da19770485a22d5d01d8925ab218211c15ecf360641c8f6809c6a5493b13f07ddf8e8bf45862a0486927a42f431f2a6a2d5c1e48d6b35c777dd881af1319d12897ccd8c07bb1ebb3b7ca87d82bd84d9336ee353e176f47f1c27d7a81f9754c8856346011930475d2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9d1729e805ed8af787e30051f508080c0b367f324f6e0f2768a7995c3d0da129deddf66e7dcb123a159e4f2b68b27d1a7e9b45f32c07126b997cdbf0cee6eb5e6092607715c9ae63783b64f18a1b1bb9297afc5278d877b120d755f14745637e8a6af829f9ca7383b72d771af495b10e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29c8ccb559082c1e3644715efb7029cbe591e5a1ad288e638d41127d2a6bd6565d9fdd15fe68c712e25eabe30cc13db1810865b1f5bdef66a96d6f1ae1e90e4d97e672eca77bbf75c41f3a65eb6aee3a7f674e4e743b3094f299549bcb9d43ba22a0f7de7608a7bde33b425ae4db7284a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5234bb18b03e2e1c0bc93ca3afe19bf790d20c039d8deae70fc43b247301b711bc586099ad9a10eec57a00cbf9d80a70bd9f57a4b0d909160634c6d8d24e2311252103fd484dcbf25ae8ea0bea3dc6a6610e331f83a7efc3033a978555b9a94ee7dc5e102a3be8b213c4f5f6b8e2f448;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcaf295e53c8b8e055780feeec67a1d99af85d341fed3f66057e28869021cf17364fca6458e11a47715084b9ceb7d7a0d10229e21cc7de06c00dd0f07526e28120a8b903837fced07f982da28896d45cd971a1a8eac500f90b277cc5de9bbeac7a1358009224fc065bffbd23e3ae4f661f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h607f77d654fd0536177283e65fcc3d2798d687fa06e338a57c44d409cf787c1d5ff111e21ce232ebb63906a9f2aa7a5226201358545e930f106ca12f08d79db5c67420b38bf983f6d2ab747c4c35ecceb6cf05d24e43c0ce3b8320a54f5b366e9311be65993d52486d4fdeb62f7cf7213;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba254902128d73e10abe2d78e106af2f29b3fdf7de7f6ccd394c6cd16b33da68c48747fe690f683f7799058ad4aba7570cfbac7a3045e4ff86577df7d851910898feef2bbe034c9064336bd6edf1e7061a9a0a207ad50067515fcece6de96dafec5818f9460e26da5a5e3f39b3c69ab54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3687eeaa4238f516d19b059a6612e45d6e316b712d4064a7730333ca75942d4f66e000907e6abe1e7aca7d55fcc8f5bc20828414e24326bdaf9d9d98b003f4ddb9ac0f81420e116b1d529e15b062635f409f8e24ca3c5dc8c60cadd0b1d690106d67e58287fcf6b82ec10c5b091d9896;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he24ef0aa5a594a1b53293418209a50c5d0fcb5f33b9a959aa66f32c7a8ece60cb5c3bd47236398ac7f6af9b662fe32627aa4a2bcb95bf3eb3d8d54890f7a73f942199880d9567d2395f90b68990fc6922993336a7c9903bc1e46290b9908805bcf48a2cec34c086ff4b4276f7b8297831;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6df9e36b459eabc4e1d2b368536bb6b0a28caaeb072d5fa5485c76c432733a22452956755096d36c994d936241e89f6444434c043699aa24c7d10d7b87720bff31623bac6ea2095958f0c1b8fe51b0eda83ebedfe6b21006780f42920a91787507d97ef49296d63d4783a6a2d19468373;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cf36a537255ee4e7da65d39ae0910499d5f57e49f5050c49be3a93283fbff5ca8c76c37883c25b4a3f4ac99a86a5859367c9becd45db185a0ba4cfc8e9b99020bd2641d1ec78c7f7cda18f58c1efd60c8fd225c1c654d662a6eb20a1b8d02b13e96f1941c9447af720a62fc5c4eb5c09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa189923191c9f3a50130bfcc888f9c16374e014c6ad57855a14374235873fc51ba7866c9940f1c87f8471d928135f033d91fd98ee177c76191dae9c15e2f0a1d55c80323197cffcf5f93122cf9844e375586c2996c97a3d6c147dba62ed3c7f29f71b6de0263699821dc5b4df1364dbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4834fef28cd78c48a37eca7a8a8ef01028b6b00b6b04efd5e784e842cc1d485735ad73050ca1f9ffb4e62c05ce31acf39c7fa13b093293a203f2e39910a5681d3f2e2606e15cef7693fef99163c291b1cb0a9f8dfcaa50906730c138885037ee6955b0fe0080762aeb7518a85e513402b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e08f26a7b608b7dc6dcb789a95c31da186b0b9626ad63c5b5412d7e2ee06c53d4ea9f3e56df23478b01bef151ea204c03ac720777c92d6f9f2878f786454e4be836bc6df4c6a841992c7a08e625b15c5ec98eef8bcf26fc96c2226febdde06921a8ee0d89598891c8f48b8f24023af7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bbc57c2d7dd40ae7339d0caaba4205d9a3f2abd79821d65a127a64dc3a7eb7f2b3babc0675c6845193b10fb85100c954fcc53f68f1829b195c0762d6ff2737dd98c0b682573a62f8e7ad258d65de64118fa459a41a94b1c2878d6816f819896fc13138c36cffac13ea78ff016f00480;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f7b9b52cad13f7413334572803c5a28d409e3e819815ca50875d0e713a8e884c1a27554f7a4e9e698b4657a38a385d83677d45a038d3313c5978aac7c670250a7f7a12d4c687067cf35be0c70176b963ef6bd7464374dbc51c31d957b71724fbcc57312208f78f3298eb487a65a1932b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b9e94185de65031af605caeeb5c6dfb264142ccd1226b12d16a0ef088a3d69ef3b7f3e1be9d03b8e18ff698a068e2538838169afa7119354047afa7e80e7fd360292506ea7c9278c4adb1133fafe760ceff50d077225d79c4f9fc1dc879e777a34c62f3cf418308041df27163689e7d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf7172e4c7fc311df5fb422357bbead5e804d1dd539a1d407c5247cec0ce98fb1b94965cd8e9bed87057abf06d55154ec7e6bdd1f232179e0a8b29365bff5f58a40ce4c0131b37362f26f58190db1b8691f78ad0e484169ee225bc01cf163c55a5afb198e2c008e33f32bdb928e9caaac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddc0923ee0cfc81bf070af2ebaf59404ac40be5762ea2bbcef6d91d6a28ad0c7995ead5af1e236242164df563731cfd08f67e1ab1f68f696b59d3e39877aad143efc6c13c6041b61d74ef8212b9273738e06f3fdf71142eafd6617ec54e16b40c4ec2e210599820d60a6a9c52bf007bf6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde57b08dfa6f688d50adad1ca8289075c2cae2fc230d1d633f760a740a46ca37c86dc51eae8f884371eefef130bb896890138d5a48f2c8ea46c1e2429bc919d8248ea8cb97dc27c4e90a56d2af491fe20ca6fbc44279bbc77f69f67355b368d36faf6ce0ee90a4ac2bf86e7b1a4936b94;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3d8a90ac743a5ed3d407eee798ac92e2da22441f82b86b249e7209f78443073d57e0ac67c38c59ff42c6e8370a0f49df262a8543fb578a889e90b7e16a7d91654a5a4665178476f45d5bf295de2572c9c684f2071312bf6d74a5bba21b73b9e7304d220d8223d454073b09f4632ebe1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fc4d97cd11e39a5cd90ff3e5602f7ef39324c8c084b81920198dafcec0d05432724c1ba57a7190901fdb2c8f6ae9a218d4a37e3b7c9d8be0bf34af265f01e7d16cf1d833eb85bf09bce701649dcf3a3f0e1b04d3b4b559945345dbc9029a67f758d3bf37ee1d9463c9fbc3821439a4dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59712102ad2b90ee01edc1e10d4fc977b7f3db2e4a5fdf8cece2cd957884302731ee6abbd2bc8871eb393ba8471d36555427bee7c04e6aedf7626e35d1105da5d2141bed835b06070dc3611f9f0ffba5bb08413a9226f1df42a398e95bb27acc6465cb56b1b76120c330606d99b397912;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dcefbad54870f956092a47d81e3f1017472884008c11499570558f46fafa5c9f7f647d69b88a48e78115faf9394dc24b160a07649f161cc85eacdc6b095d03168396dfe0feb2d58607d45ec0725620345ed32c62e91ae375efc749e07a499333862d1f4de133b2dbbd7c6f71431538ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97c4fea5bc8b77b1df1faea3e6750d8b353b72b5d3e3e02e87cd358e6db69e58021a9570126ce9829963516ff0a3956ff011c59edf567a7577abb5fa3bf2faaf08115150117ee871cb7d2311be237c5812c93d1c2b2a6621cd309e374364d376012bd4f611865514c94640814f04a80a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a4e47645cbf562d01253f7dcaf03d1c903ff0a1b7362bc1ce8e5fcfa67141658ba0b2fbc976403f3e25469e609d676d7316626a25547d7f5f28ba9a6d6f7a085a51b1bf623410e54759c73c05dc49ee2aa6716edd426c6eaf7fbf65de023b34cdc752313f705a051bdfd0482213ddf9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22d534a65f6d35867548a713829e42eaf88aa3962f0ca30e9978ec84cfcea7786857c9bcd299515ee440e340c8353c532fa1e85e2b8525cd7e49cf1c79202b0f1216da85c71e5a658bf8d2c4010dc4ecdee8b7892fbee0493399b4e4b6f6f143989e1866d0918887973173736a1b47a9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bb5870c830acee6a112dba8e27181b7e54a307325d8bdd8aa0554e0b3623595ef73f7f249a0d4b6413c3cab019c926cd306e65dd449c4605f32f18f10e441976a2d4cc5df1b07c806d608e34c105126f5882a6ec4dd630f0dc8bde08501ddb8e78167e56a248b1691c444421d3c83ce3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d42e5bb1c658674173bb3eb7bd9f2ad4485061cc935e485a6b7c02b7dcec9654533d395b0a2990494d7512bc39a772aee1d6d8a92379874dbc978a657bdc2ac4f746ad353240221fcf898de05faaf6d944d636670c77a7a0de08eb286105ea63674231d7a19a16efbd817f98cbd66564;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h947823bd94162b6e4c3f488890d98adb010782806321242ce11a31e7f7b6c89b687133696ef57151351f177d9a90e0c8d58788ae766cf79cf69844d0ba87811c6b0c8be5ea318db2d972e20ea2a2483763e68532018fbc4d480517f910b0e5f656e326725a5dbef9eaccd29b1c5f874e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc89dd6e0a15f35c9f44045d172c7be7a4223390c293ebe38bb7bdc50c9f83b3563456782b9663ea5d896f1f1b7f735e8e0c9af61c74f096a7e0fa5817cc8ab1766648834fb25732b338eaa80d9eae754292aef586d8e3f7e4040322978b6dafd635044f99528123232d3691967bb7b588;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h953012848a66e6c06de02acdab377f6b6cba143d26fba051bb2997daa975397d9c9f32e7bc65c9edb75b549d03bc5a3954f83f43b6efbe5ab181d32194c81c97b7740e559dbea40c6bfe41e6ea0eff9777afdc1153279c1e6323e3bc4f37cb30661501240307ef97d461a91ccf625888c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95347b41a177c173cb5d32411a4adff6e2ca4e78f697f528916f690ba736765084a176d9bf2d97d4a42a74aa42f8f1b6f1499422fddc25d45238a8fbabe285c8bda06bd31e047dd12b1cd918053b945c57e1c09d70f38edbf2e42d6a146e7d7e003151de712e42928fdfd08deafab80fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75c8653e6434df808367c9aa74528812588bb6512719d5cec8e572c2c2f81d6befac72837f058d79288462927d957246e78260ce91817d3046dce085944cd1e1fcf838af3b39a89422ab6499db5e884959e91b4c0d4b0a63c5059b2e2ba820f316fc7e6e82aefc0c2433784656855c30e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc54156c871f7ddc13795c6d0f51db1b2eb5f635cc800cb6db9ffdc12fb5af1ba7e3bb7f949659de0c2a1ee96f68afa2532050368b2e2ffc9e417dce0e70c68763bac17ec3646add14a51a17973005406cbe87eb87019f6049d8e299483e452d8da9e994a5dbf46011c8219f20a8aa08be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd579b71d32fc3eae030b3e1af90a375f85cc72ea5ceb4faccbdabe3f12b2687f5cd2027f2078134d1a908ea7d55343fb535ac25eb4f54a35a436dd64f475d9e298df3c07fda9ffc4b8749b5bd9b070b405b7730752af0c535478763b8a010bd82b8fda159970b81ae913637d03dd941c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaceae88239a8ec946e2168943fbd87f51f708a8b614160aa80864245f26897ee6ebb26678762a06f87090477fa0f6c255cf24d5f676b80a768a460d1407bf9dca1ad23f34de2c23e819bf375d2dd6046fbf60cb4add2c5a053a93b13f7d975169daa8cdbf02277f812bbc8b73cea1ff6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h354ab567c421f40978c3dd441b563459d3aaf84289deb865bc99aee11860ae645f616c46ad59a64e617e7bcb5b4f79dc3f67e73af6bf3e4e352a7f9cecd710d37288777caaa7d24ac2d2bf28b1aba77b311511eeed4311fff9decd78bb25292164984ca0ef3d463c9962a18086477ee7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he34dc79014c115b92b46c3fe1314259bb7b8345e20dcf712e4d9dc8ed85a57f52139a5421dd7eb7b248e2562f727129d0f74b374dd073cb2b41df051955bde366a6df16d8312f47add805bdecfbae00fefcdc45be45c127bfbb95cd45d2393259c792febd105ce13a9722c0b1a99dd270;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedbe902c4ca0ca09ef3018cdda215db1e7d73cf10344a5777c7d0be71188580cfa4358effd59818dd7445adc4b12c6629d6515e63c26dce22f356d52cec884d2e266d8ef62355073be4bef14fcf3a27d509c0c6a5cdf4b195953b6c5f9927a1788aa4191c8dc81db57024625abc6997e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a016a2af03ae2efdadb473ae48fca98e226fc9bed5d9dada0e771c4c08fd15a1349ec54c57e07e7b95d787398e3d6ce897ac22c8048a92cc9847d344c7bf4043745397aad612e44c676ad865706ea2f4685dfdf9b625ca4b9c16935d98990fde0f884475fc1f604124226d2310ff9f2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb18cc76f136be6633f741413df77a5de1b1c72cddebabe60f36e5a021830bf4e272235f87322fd60a0f103f58e9f95d51a3a96126c1a49fbd0feef8b17f2c6fd85146db0e1b00f482e5a8ad1e788d309662b1a55ceca7b794949c1c4f263a8119080c8e6b3b776113c8df8057af470e6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cac1dda1f6bb30f37bb56fb2490058792d0389cc658ef0b5f3ed1d2771b89082f81b78e18ed0c6b91506c15b6efc1417c37e96e51ac3fe51b115e67ef9423bfd66286161bbba229c2b254a1911f7a18abbfa23dbc3e4c83c7065595500a0bf25599e7411a337eaf861e46f13f7e50b32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc29f38efc56cd7ee802c7891015f910dcfb8705d8633fc6ed5b4c31a28662d1d000d8ecb61212510623b662b9ccaea828d7dcd2f9852e0d2ee0286d11637635d2afb458dccebc4f7ef17bd1e348ef7d4d2cf2256cf1186a17929dc0d858e64bedc9f1143324c5c6f2e113e93165add0e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc526ad1111cf070a4dc39d2d067bb502ac25814366829a498459c81c7bc3f3ebb7a75e5b37b6e568b2c0e5cf8536a64ce333f3f4ed312a3dcd5a8473a93751c1b54943befdc246f6feb5b7be1009c9661dc5dcb1987acce2f34a112b13b4f9a243fdc8f311ac73d044807e80e097067dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdab20bed9900fad2f4083d8db8409a77806040e6a5ec210f9f4a1f3615b7fd1649d8b208ce60204fab7ddeff2efa2bfcf384d6ce418e39bfe52e0196e186bb4ee1dd136c01846955f7378bf811538fa4637a7e1d7bbc45ec912cb19bd7ff3326653dcc62978dbf724cc811de688afee0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h996854b4a05c7b2d5d17ee84eb4ea64efd26098fb97a208dc20b8a4c60f54c2f6cf352126349a9a4f431bf9a2e4364672b3b760dd0d2a4251f366acb2516e0c00e6d67fb2235b16090ea028e52940c0739dc788f938dab1b5cb4b418fa52c96a61a0aef7174eacca2cc8ade92682245cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h908a8839037a767746def00b8bbe7a71262a7fcc54852792dae07e450bbdde14ee032b7a3d3e93e708df7324e440bbe8df19dd92f53c1a35e3f439f0f1851163d37e56ac582ef912b1e04ed61e5cdbee96098e61089ab77548f6c48761584926a19c782a5fb71cdad59a81ae88cca81aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8376dd97b34baea3116a21850f8d32e60841321284d484903c8baef0f29cdfaf99f1ddea19d83321e63e2fd939dcdf743b4300f46c391e761c611b57ab411f6f22102859ebd9196f5e64ae3badb49d5ac12d7cfdbdec7f319ec0b3406102e2d73ada895faa6a08e034dec24acfc5a3058;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84f34181989ad4c481dfebb11cfa0942a81221d1b6157cf3cd6ff86241d8d890019efc87651a79974937d0715d3d96af10b3caf4e821e85703bf6164a748f73ef71ee78ac0df2f07c4cad137f0b48ac31c65e872449e40a508a3fb0dff3c24320b8a682aabbca3a3b55515e8682e6319d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h555f2b914942cec7cb2a79add8c84aa87a218dad8d9c578abf56d0b12a826ffe2e3f488e50e6c81b802ab40e715d98fe52eb031d783cd4314f7ea4d696da3098f1ff5b5fdcf80935e71561a5cd0c16b6aa2ce90cb4a6d0ee8914473182988548286dff4379db8e9db2dc150404eca498e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e386fb73b41d46a845f213f63f61a3d33b49b033827742b269ce07bdf8800678f3c4196866497bf530f1185233648d3934fd584b0061481d1f00209e26d9beb7e28dedfc9b7e4e821fbbb1ebdef67d7ec6e1d896d0b433341eb59780251fbb59e5e0560adc35f84813daf0c6f173b295;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha98e93f7c527ce2980b013a8e387e23f4b93fae08b9cf9d71c60b7831330ecaf1a00b72a7e705a76c058f574d2e4a1f570fca1f14bc243db1a7822d291ba4b0bf2337f46c00cfa80be7891551a030985457c2bc962616d6379bbe1fd67adfd7fa8e2296320d0661a82fb3b2b9d1ed0fad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h513d3714b98661aedfcb5063f0d1d6aea4252976d163e46a6ba1bc11659ab9fbc9d8ef66677bcb109aae273909a90afb4bbd88467695ab93956d8d676cd8f7692b02de4434c106555905f69e3a275d2ed4b2cd08bc9a8543a57c5910995d1ba2e8d71d071aadbab29cf93810583d701d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9454d3078429e8e78683527253b05864f7eb96fe5111c7f1fe1b9310119e645d05b3de42e2cbab591ebe0f7cf603622c916bd250987160b358d5d5b2406e428d421f045c57a53f500ebe7e79857284f2d011299e117ef658411ddcee1d64a9d5a75effd509a58a6db78eb2c6a69e33a03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4842b600ec2e2af6c142cd1c973d9bd7adbff71a21a26e61c00a7dc82225f2ff00e0f4133199291691d58645118230206740fd4941d1e411ccf2b8d50d319732336ddb18be254193265f534ce20ab55dc891485330c8f6434c6163e524e355f1453c762885d38267975bcb35c4e609a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57edf1096ca2b09982ebc8a80da0bc85d3d63afd84e1846ec9a7d57aaedab79545d6b4e5e5b461359086a1c7cfae1ed0ec413cdc8d1b739f445b8d32a4bb474d53e03f09a07faa03ede882c73825f24e070d2b465482b9b721432cef84f63d67595869335df14bc162fa96b310a13d262;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb12ef1e5680eb3116a5d697dd07dd88428a3d8fd4479b5a79f8cfb0c33104dda6cb7d88b4f294da9f17dc32d40fbc04837eb9c4aadb2ec85fcd6f551392660e12d85462924e5c86238f3a25557d196e8e425d0024d1bf97745bf075aae7fbff7b4159d2a941d0e482efb27fd7f4a765fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h713a7c5967b16bb73dc177b580fdfb4ebd17d7c7b5f38c560ff31fa78164cb4976ccbb408cca048b9a5268ace403d6cbc3f9f7c1b1b55a6d284b04f4896b132b06ae98ad1e12e54e09d43a96c50a1bb47c49c32725a83758c74d359508316e47470338fad2f6f8db4c202975986c384b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h789879f6b2fa874e1c97052d194858ea32db6c413b0fe97928121de30e8d9864754e64749da7a2594540fe8e996ca18a34494840f4db9108dd276057fe8ec8a2b17f0a0836e53d141b97b3c3b4c822a8e7f4ff6d79b0d881c678fdb7c41c9db66aad6a8c6964b735e278c32ec2334a4d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddbf13e97713c6813dfdf621eaab7d7f782f0a4eae8ab1b794ad8fe54eb421ba1c04c9006a4225aee8df6165f60fff756ffb8df4b7844a08954253cbb22da4466a7bc31d51189bd0a32c92a8705b6ad94f9a9ee644df96ac7462f62cfc4db637910f4fa15acce259b6006f1febd7fb11b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91af954ad61fbee3c5a2731d7f7ce5c1f0e7c8a4229ec46e33d98e0f5e386fbc134f5446500fa54330692b7c19fec3d9e44449f7b37f861acb1a21686e4eff6abcd3426f5280b73a78fc7360737657b130fc467d8e036e65a932f7f6a7777c43fbc829a76ccca8a38b7a048b215541a90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb032f1bd598cd945da1b9ca9a7565b589871f616b91c1bdb9e7fbd9daa4a61a7f0935624f692c131ad2f2fa971a142b3bc031bbf37650736a66e1024666fe490d523c280d7580660eea04ce8c098a3f68e4c6a10626809306cab682bf59043bfc9c9d44bb76c5a2da65399f363d6fbccd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9a53770f85ad7c026385f77329651053b3be5075c21cd77d9ade6e6e234a4fd82659b6bd1d4d5bd1165fe74f1f92bcd3f634fb688b1a3f78b3ee346ca530098572957b77bdc8e2b6346c40cd3b8f1babb374d085ed94a34aa0208d44505a772814942fd4af5160473e166f3195060564;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c8e4bf717bc608046599f768a729e51511e04dc9125ed137548a29de98ad6372bacc999c0b413449fa609aeee39a7600e41ba4d6deff57c1f0ba4065b09f093ef892858ace1a6019f60920115802987be1451b3216343374bc523c183ae85cd4a5ecdf00e1a47ce98c5bbe237336d128;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h309f970023fb64e3e9c82803571f475ca0787d545c9f581569b55a1b7eae73acf9038bb9eb8fa3ccec675edd373afa33e94cf27234ac6a3b876062b4322839f554c605f1b2bc86a73875d29cbf870f99e5d2f8ba3f5a08c467a840a03bc7ca0654e7328992c3b74c511fcdce9c644a239;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9c2dd7f96f2e744886be53f4097b086a1b2e0eae2159d32c056444e2f83a1a025f6b2200ac2edd6b26ac9d4c2fdf4b196bb80fb257da56d50b902fdacecbeb412ae99d4e694d6b38b39fa46f6ed05194c05e6f8579b59ab9a426e5fa04f1727b3215ff7b8f1a58c8265dd7f5feda92dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedc6f005ea6acb587e06736c56fdd5d16fba9bc4693ea72cbedfba3e2e7c7b596b76f29aae0dc8f29ebd3289d5b010b0cb3a58c5cfac51576a15440f9aa3915b239663f10d3b6e59ebd5976cc49fe9e649fd2e548de0a38ea2cd188e295bd5c4dca2f9a1c30ca768abbfed65e88518ec7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4ea164c74f8496530522b6100bd81fa98ae483e23b4aa8c744c17e2bbd1c26d320a4609c96f1eb273120c395175b46e883f8f421063e05e60ef31829d759f408344d800fad6e03622cfe902a2537154cba1909059d00caf065bb809a2aa0db3b1f57413b746aa4ed8895a692f067751a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h749d3bbf63f783df39c7d988d9dae2dad8256ef4107d2ddff4e72f3ec0a525d173b9b092ac3988a5a456c23e0901359917c6218c2afe807a8b1a132c100a14850facc95b93121ac452b27325a566e81341b26a47ac00652339e1b76348b0e1a63dd468f4e2d91e4dd1e7fec078a7c4ff6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7ade8d385adfe4f898d8d72b126459d9a378a9df4129e76813aecd19c2594708f7c23cf9bc0baa57d1c0b36d45dce9a4161e16cbb330165a785d212a2c7f02354f276899454ce90a2fc58cc99d133679cc3b4aed0b0583dfa022627c2bf9d7c2a12a5580ccacef07f448f5886577c2ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbec08ec997415a7bb95cb1052b9f1483f2fa267dee052dc3f11988ff735c437a82a8a52232b26e8a027060d4ff9fabd7115e51482873f6870cc9c9cca0047c07ddf0e9454da2af2d00b34c63879be8c2fb8537ead9b9153d5711b99fdc82e54bab5f173abd3525548d7385ec473ff9ddb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98e41b78c73714fd4977d9a2b4d730cf771de42b8477bed5442668f7fe9d6d7c6da6a1b1c730afca181ee8945da4e458dd1985bdf0425371e8622641f947357bb9601e6c2aa1c94deb5c8ecd55889defcba4bd2162fc19ec8d026cced0aeb48f9f1e6ebe875dd32e194cf7f1f9629e0a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h981da72af8d5840943d8b45a2294b83e517a224238adb5dca91ca59b265e5136c51cebcf9b44534ef3fa370e683ffc1342ee1ec89d056b8eaf6cd69fa0bffe3ef46b77f54ec61bce6f48cd34e383bfc96bb37a11f4915080b6514dbd236545b356cb71408def90ed1e0ee6b10ad6df3f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39d79fe2aff9133f7945d4b6c12d1ad99ecce51eeccff9f5977e74e368cf511216acee13f8718a80e72c0bf665efd4b277cc1537ac71d83bd2899da7d70c725e74c0384f48460c24718327a102159b5467025b97279f3a84fe3306151a266a54224d28b4f5f790c79402db64d475c3077;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc43caab529457fcfe67e1032d6cb8571891b707463186d14274b5e104ccafd09bd6cec6d08671d32146dd50ce1e960d8df8524f5d581b04b50ef65618b6b9b7169fb5ca47b85d99657909affbe413f62ed47bc228fbea02e4d184c856d7e645ee9ab93da9894c1453ef9f309db56561;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfbfce9ec2c6d358b7edac3f7537591c147a05f2271a063a12106f583a0db40d58d110503b793c44c4b0b3c88d403e18e38b9f38ada49902df7bb406924405f2dada33dd2aa7e6192ee7ba42237dfcbd8eb44cafacdb1b4c6e2ea68012ac76ef59fb46df596de1aa25495c2030aa04d2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bfe7271748f618541125bbf30260be2b5b7dcea26c91384d19e2ee09899d46ffbb1e910b7775e4c51fa37e4b654f784e50a92683ede65a71795381c249c0a905d5e51d547b654110dfcb0eaf918a1038a70ca1029e2fe3142f69e170ee505cf347e942360b865f8c31d7911c02ec504e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ed0f3a12e4b15e28ae159e04e067104b6d26a7e5984ec48887b8758d01043249a80e1c84a6e54dca90d860be67ff78e8c96a0bc4c548cf9521e71cf55abcbba03c5c4511757c96564266f396359134adcf5fb13aea63c34d4db3304b9253c0ea5458e0bbc79a55e96ef6754bb7b7ab7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4e1c4f56f8700a4fdbc80e49e54d2eeb42617436b2a79af02cb1e7203b8e3edf8129c1807a4849acbf209270635ca24ccead95c417d63d1609fae0407b12a5998b0a70182e157a7d4182aa42188ffcefb4785304c04bcf7b7db734dd85000323807a0f348a4dcbc852b1d35e7da8f65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd241a64897523ee48b907c58695bff7cf4bc1b07328144260960d33a3ef0e9428dbec4db4c72af1eee6fc8266915dd6ec8e974f0951651771c729b825a458514efb4a4de18d0e0c3f968f9cf55ac90f94b47e680699d6e4530dbba820a5dd99cdfac8db558f2f4e78aa82e7eb3cbdc185;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc226c1966a37af49fd58d11ba0e1edf2f341a2a830af637c5dc176e9c13ac34ed013fb65bb4c0ccb3dde2bbcb66d5d7da707e057468c0ee748ce5f92fb916fa4b585985a54e7ccdf648c76c202fc1e80ad41bf9e6d76e7d6a1a84e4624dcea2b0753cb069a6db2dca0ef796d3d11d0852;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90b69b82a9e1f21fcfdbb288531939e394ca39c362491e8a4a88a8b04cc4df7ebe078b46ce948b751b4a9d8f9b4800b204399938d5f914e2575a10d573bae669bc720d86048bba7a13b10a40deb56458c6379fdd5ff5b9a602374a38a41ede97ea2d3dce662392b5e7998205a37eb7e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0f69374c9a7089c89951645ef8b736c125c1dd198409285607f4d590fb43c2bf11b848b76724a6350c8e0f6a60087c5fd7b346b1ece2e92e6df2a6b35572e621bd0aeaa1726121a4b6a1d31becb5d422ef3c59f651bb6376bd34c5ae286bc32db85479ac634bb54e2cd528df501c008f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68d925f5e9fe4fefd5047b67f515f9a622ab7e3992577d1eef63c942541a5082d1b1c00d1b2de35570bcce93d3699897bf008b3d57fc0b2511492a1d9ea34e93336f98776198d7965321ff6121eaef1ad2643c09b5b600c5c9c932538cdba8d406a4ac90864d2899bc1b4eaf7888fe340;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b920805c42086178592f934062b9adb0a93abb68de6a80c858b8617f380efe0e52e59248eef1613856b69dfd0c0a9ba30d3fe91cfa9fd2e0b8d68223fc8b45c33eca8a70a7d3d982685ddf400be29c41b97a69cdf444b051cac97c27c0ee2cc276b22f2e523b0740bf912a6cd0205ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb359f6313aba88b2b25145f0e1a32e890523131f282935233e8f762505b8d530224368fa4bfde8cb03baa0ebf8e7cddc39a6b5d63b9c8c8170fbae94c115ee0d0500efedff8503aea5ec0e8d63f20bcd08e494ac140b894879c1af4b18e51aeab6bed70293f9b94014c371707efc4ae3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5552bb45791b58cb0463263a056e08fe0b2bf8de2f695372fd3bee0effeb3ba25155db497900c6ef97cbc93ca6ba5b91af7115070d4264da42bbeb7f4437c19752aa24aa359bc34f6b98c79b47e03102620315c5e7134dd59f687dc7a339c3873e1a875292e0fc13a634d2caa3b334af1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1362415b5d51d8703b574ebff0298d34c0279d3e02ca70600a4bf9e555f9d21d01151ddf64748793f45f3bb17aa8eb7025e32625370f4f2acde88e5a456a9ad51fdb41f2d4a8b3e05c80b3ac3c3b3d1c4d974929d19b1772c77ef415b66ba87f31f4bfbc559d5cb696ac8e01de771e95c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e92dab3806998b5942cf34c3ba25229cbba814f394b1763571073398f3a62b85bfb606d4db6747fd42121d95850f4770d536d4ce1b2b5184fde44865c213c714a61ba15246ee735266836fa0e70d6a9ee27e20416ddfe9138e3084fa25ccb1eecf3f3bf51b72329d7f1e978d6bd078cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf161f00f1b2fbbb70147d58c431e1c5a8a2600e38de73475d1998e06053470b7b4b49b66fcd8acd2624c75390710603f6e83171293f676936dd48446af84bc4867e45a694640f1347b4cd78756b9147867a94225c2512ae017bc69034bb66978c9ada3710d98a0960bd2844ca8cf6d86;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe7a1235dcbfe23f2f4ae0bd0d57f92d6887e56d9517f489a9a77559804bd6f9a1b7c97cdcb480c2c76537e518f746bd7c0fe75a1e571628342bef28002bf3ac8ae783b53a42f37858f2fd4144998b9b3eca76175006a62b7f9f8d644f3e1c3cf6a5f6774f0060e6d2a672cec4448e94c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62f8da08e640d8599826706223fc7e8013d867464b315c437d9770eee84215904e40eb6a132347cac7dff43d9e4a2fbd07f4bbb154505932de4555a4e0915cc0ae6035f09b3a9851fdbb49e71fa275bad18aca3feb6a629bd9370c49b6c41aeb354512e21eff3ce858eec0fa6b7dc9e53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf28e9850137e37516b80fa6e13898965f8acb17bfa58648648226761160e2fd2e5498d37036b7ea2d96e93827634c16a752685c6b61564c3bc29b336c2635b055978b427cb69d2425b291d81712e5bccfe321f1e7ce2ed5aa756324293f0c7f8007c77a0000c3b49e5f0e7d556133123;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c80717ead19ab03d63d83ae4a9eec02bd09076b2e42e1c227339055a91d96505179c3f914de62a3cf232b9f941d3220687625914ced022536428e71b6b945376df035fb55ba168f29da74b4d35c42ec334d86be18d8b963fa52ef81ff8445d1c1cc42b1a9f789b999f4bb6e41d8fc142;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a67134ddef5dae2634ec762c7aaaecbb8fcae2f0be9c9dfeeaae50ef6b5588343c5ed0208c27096c907858c49e254523c550386c3d1aa8d28425b14b4d44509f4fce8d8d8e38fddfee5ad539c03354226b7ed04d89c791f2dd5584d3fa5adab2e9e41dbbeac6b669b3a4a2e265ba3c05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb161c7476377bc9b08e88cbbfd14ab17c00b4008c0e8dfa805bf5de707625655f90a5d5d50f0bfb6779c83ade120fc062c0469101cbc4ccde4bdbf1bc35416e2f15d81238066cf51a501ed4796cc06f253711e38ba77e736c3a65b84a826374b1814ea4401d5db6561ba6aadacd94da9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2189a8473408334854499be6e127bbab23bbc396bfa854643689895299cd27e7666e618a68ea69b77d81951fd36cf8438c8669f92603c914a59df89691c80e042d4d6b2073d88cf8767bbb5bb6052530992f99b4899b1409310db6eeae83a4e9ca80033f48281adfadb0fdf7d5416b68d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b68bea9670f465f7a5109a047fffef9abe59a6843f0dcb279cf5ed2c390c9c774c70f109c5e4a32943c5fef60640cc680e0fdeaa250c88bb9e860e0820cbe8c9c6e3c51a046cca3519a2643da72387c606acc684d2e159836b20c0bb2cb87f5597e357a84acf9cbfb83bc887f0732c63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h196f378884616fba98e2f25a402ad974cd776ac265c62708ea4a92380ebda19bc1770fcb8c37274908b0c6f6102a23f3720c9cb8d967d37e6796af01e98d741c9ecd2f80b3147ace2e78214adba775608d1ec69ed95f09d720bd597d44ab9a6329f03ee201266108f278a8fe25c560367;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7b67a087270601dce5a840d5f966c2ad2b1cea6daa8bd9b02319239efb4b604f273d5ff3f3ae17ea7102f87840a046390eef3726ceddb6977ffd0296a6b72a0439f96c74f705fa55d02334db0c785c6380f8df7bc8a1ec69cece1752aec98e092c254f4440a93a9b09cedbdea4de7b0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d73544ba8704b96fa0d5c1ab922fcdd95f59fd27487ddb7a9ad980b8b4402dad8288f6953d56759af058cbb71220678b19120a05311d35fb53af768fc47775367345cc573ec69eb77c9ab8250aa2954d9f79e164edb74623ccbd452a3ba866742fa86602abdb4ec263e8cf70a8ca473b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cc2a3ed76ba5dd3d1225e451f6f8e9f2bbb5545bef8eb01144dcd9348b58b8e5b5069d56a255461f644b3c24f7b998811220dc261e431a5014ef06c77a9bad0a9d6866f3059ce73d70a75150cf09cdaa6d4112e6a2652896218cab14e4c6c47c57cd73d8986da151c4e3841e5a37137e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haade0af386d0596d97ce5bc78c9527b79fa7f0f9c8bc976d9dc53113d16447d32c79ae806ed7fbc8990d625d8aa005d9f1d501cd478e12762ef6ddfaf3bc59e35bd0708cd13204ce84c18bc0bc2120392b5cf4c7f33841c68ca031f7a32444f64c64f88999f771cfe6f3bbddf338ac8d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40c39e997ed4b70da5d9f76bd19fb3c867fcec28912cbf332559c7979ce492526213aceedd8cc06b48030e7b0550d440fb608775e5e691fbac19543ca962a2f7d3221661231090fc189737319790b298b3618a266c0b189457fa8c799ff0d29215de2634e1e696069dc9e7acf8dda53f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46b0cd310872daf89ad4c3e916332e43187dd218e88a78dd9167442e879373d77226d6a928357168fbd6ef10df5edac36d222f2f4636dbf3f95a5f47ff66c479ffe151ad01583d7609b0abf4a952ce6849aad61e6b0023370c0efc4cabb040f3f582d8e207c286bf346c6591494ec60c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb0a2219ca182918e5468dca9d51408bcf48624c7f5b92da0bbbc456966a034fedd5e8e3fa591badedc2fd21dd1023475ae0c3499e21eee10168d76d0ef6a8ab191c61ba660542b35307dcff2ee232d0212b3b8279f4b9d1a05f3a9bb9466fc8a5334bc06b5ffe7d10a41f8541e54643b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b4d802483742df636690dd3646c30ff7ce22842f244d618083c02e575629b2f87bcdae5ed78bcddabc27918bb98800d3a3ad0e31487d27694d86361292c38e075899368100abf60f17b1beff7a0ffef234b7cc807be91248473f8769cf2e87061876853d98820af11a4440b04dc2d1a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cc3c11cb4dc7f2eeef511b408c8139bc126cba65833d7c9bd191cd14e0e18345c567988347bbda172390d6eec7cd31e2bf7795b84e69951ebaee7c64135cbe395d36a8fecd49a46000be7995c6d7e8b34f40fd8586f4e1ee2af651568fcaeacda3a5cb7dab7056c77495f865a5f71c4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78aaa8420ca8eb720d36300d47cdd47f9600141b987c1357b87de1ca4916660664c6eb761a8e63b35905f990ae267b236df2fb79a59cc194cbe5de39ef34075c1c434a20cf0934c6afbbfbdddaeefa9ece5f90a28a858ed862a71410c843ce8e021f98eadf563f2b990f19a58dce1ae85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51feb4c5c8f8bd52c1a7e2a1cf7e2d482433054a4dd77c9a8db3d4194b06bd1bff19599dd9d07a99f747ff6bdd612ea099770069d7a9b63e3145d58f02c73ec7c8e2f0132bbf964cf383a26deffb2922554d18227acc2f735183b64e6307fb5acc3cd714c4073b58aa3b3beb060caa2b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91298a84ed80e0fe0b05ab5f06fe9987f7d7d1374ab44924319cdeff2120385fc0b2521553dc8e6a491e35f8e14771e746fc07d9b796fa3d8912c89608b292f6330cccd445e68e01f546190402f4880017436a24fe9686bb159f6bb7ae32864cc1a0cd2272e94dcd319f72353a03bca2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha05ad2266d2e8d048772e8c12e8779f9aa49b1ffa6ee46a7829b45896f05c0c29cd3ca9bbfad052ce8f1482b103f3d9ea1e689efbe288f76b68a1c9a70c15f11035c03f836c9bb8233325e8d06de7e373d016bb228ca9d2f6aae6ecca1820bdd95fb1814de9751a9a9fe1ee598789fcb4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87587059003e85ec4bbfce98d37f0a85bee4399a883ccecc9534ce68dd25bcfcef32d792b28bcbf009703fb4237747e68bcf57d69e9f7c427bc28c51603aea4f042390b9848953473db5cb75c408e9bd152476d02003d901978fd7fdc3cda52b827a206dfe1ded56962bdaf9181502ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a47da493f1629fd17355e307d94e5613ceb50cf0b03cafee5183e613f7aab0eaa783e48e23a503bbadb78cf6fe2c81fd935916e2ab5de7554317c110e20350aa3cc6f04b0edce68c0a844f43f9d85f9eeb3b4b482760174366827e60651987c210936269bc0641be93306c6488a33dec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78205872b24fa57fc1bad7af5e60a2a142a64b6b2189d40f58f8255fede29de17f2c9b3b7d5418f5a39e12f3bcc99a0311505da5027a70fe64b99d6b4659eebfdc4386cde62ac3424b03cd9caea83954d02c98d7b756b7ba33273fad79b3c0df9fb91c8b7fd487861172426b15ecd6f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd50d118a106b2e7ef21abd5f64e2ed39a41aaaea76d9c98b6557dc4f4fbec82cd6760129d143ff31f592452f1df52e66c1520509a46ade6bc999284fc253d64cf16adfccd8967a7bf31b3b01ed6c2cd7146e231ebb58fe3e74c9603647c363f078b188f2e178295d587e356b7aaa236dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bf67c6cc4e7f70f07ce1261b704a4aaa4b43d69296116ca8abafdc246cabebc7aa86a05cc0f775d9c3f78da7bebf2ef4cd39930e08d81b022655a1ae001d0a6098f46a2c7f09fc701d2a9d28502f880b864083fffe7a1fe86af84c1cd1e44dd8ceb4e7f4af935e19801b39519b057d2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h280c2aadd3016234764dccc3ba0ed2fac6e4dccabc2b36616e2e3c31615e2e48e2d9d27b4ceddde4562e032898b3c0db1eb71bf4fdae9b505e89fc24446c8d97181de0f0af65afdf948e8e191093c2758012c9c69a14acc12bc5128c6024fb1af77d4a9bfac01e255d6f940f7e610faa1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fe3e99785f5bc95f17698ce09f9b6c3f5590b236c3a6a18bdf8a93ae558d8f160884a20e9d280d98eec498afa7f7d95f9a34fc0c5e6fcb1dc4ab310e0a9f742797f3359a185e7d3624aee26f927daad948ab507f928453aa1a16217d52d4f4641a7b7f680951e4c169f1891bc3200962;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc522005999f29877e3f8b2ff6465f5ee6f76c4b12bd6d18cbbee311c1219daa34ea06b22d9dc0445010d8155d1bfb22adda8eee766d2d72b7fb2b7ca886ed346f7f6eb4885c9a665e0af081b376039f4413328736ed0a9a43e2ba8cc28b53fead77cd88693254df613b244d506c1b0c7b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3981bf834a264a1fe39e4edc5c7b3916fc754810c35d3092ae0fe16c1a07706c2d9197ebcdfab0f11f18f07695edb916a0db77dc8a6e3199964ffad7d4a4cd89db1741014863592173e2f5c1fe811d942a95a727744b4159117317005c5f5270541717ad23e3f94b095cdd8787a28dcb8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6145ddf8a9a0e01a6b24b17d21b7475d529b96e42edd74d386551b00b450385f57b0c169bdc7899dc03d0f5ca5788fda1effb8204226641d3670049e4f91c5ed7709415d85bd0aa3d240926c8621019c6b70323e071fc8d264e771e0654fdc0a9c366963ba5b94e5d0ec0f84bdc6c020;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d9340e526e4354a1db8d3506da7d1c8913cc113e9d37a73fa9f5ee0658b1801a9fbf313091aa43f9928621fd875ae0b8feb08ca2c6544c5f5edd519c9b8f3befd52d329c906f8155976d8beb384186c4bf7d4cee30631547bc64a73b67008e69cd5e5931a6382ab6e4cc58c80493645e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e0cc05ae17ecdf0cd93fa526ce784168e9dcf39e073f5bbd95abd5b04ca7c2b4470c05e3d6194e35bc767d6f90c6d497a9671cbc4aa8dce7c1200053b00369f97578e5b3a4e942f44cbe8fb5951536c97668d3d773ae94883a0c9d2027ec2aaabc9ce96f96c139fa2c5f600e58bef62d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34fc7f111ddce0138b43db74b4448a2b5baf4c1a6413b572729ed60515a1a4079862929d55fd9e824bb2311a9b90f63f1a97e7519b23d28dc0840744bf16969f938259f8db04a7639fb78515e46ebff1b1830cdf200ec1a919bf11d3e83bd65fc9080f82ea81e36d5f2abdebde2014583;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd55e531a6e75d117ebed2198f3dc6786baa4132da5c77d4e5be67d2147c1d457c931f573a1172d0de8a994acde1e43ef7c8143713bfede53010881c137ca37138d798a8ffcf5af93d6587e8011641f139568ef20cb4154f7178d22e84d70165de5d3da70dea299da96338a0bcbfaca64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32969c92b31fd48e4a2db2459d5736cebdec3473fdad644808e172a9ff7ecd2449244fa880e6eaaf98a05989eb4c1d90cc7800699e2292d2fd13201f4d739e4b6fde059761f3dbae486847eed8fe9888ebfc97fa39309a97345702909f88a031384b6cda960490d4a2b83865f266f1118;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfb82e077f15c5f47b4df1d4e679a8619ced11d403feed5d8340ee8207fe74c85b907f33b31a235b1ac7d1ea23cc6ea7b098ab5e2b82000244c0f05ff59e6fe953622af3e556d0a9d2fbf317a06c1e45baa43ba6956b35cf9e16c7f140f801980898373c7798f2a66847f19d7d548a6b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he762d057454207d7bfb4c637314cd21c760cdd4e8795cde60dac014ca7fb459ce24d27f28955affb757cae0fa69e57f782bae7e3ae93fbbd8e0b269548f16aae897123e65a331a472dc3d1794eee54b651e350ac68f38530a070c4d5274352fbf05d18bf4c48b4e64ab5c4515e918f08c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2360b85932e4d31c1676577427c3d80f9ac46bf6d19d526a22ac669ac23f0acbe7e0ebfe9c6b7d40deb0ce9cc3d313b2ee8b8497ee8a360221704576db5c14e273b51d10e41beb1e63db9187fa5c52dffad4b2c654b08c2588a7e75cfc34f08b3ad549ac44ec1345f18a283f436926526;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ea3a316d8465cac958d9378dccb8848670caaf50bbcb976e675df89380231c1f018297873b5d39695611d07a5c38d68dafaaab02d0564811999acb05f64ded3add2192cd095f7147852fb412f1c5f2a298dbbf3f67341e75fcda2ad27a6ae862987e8e745746dda81f27aae4be22a399;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7b16c61e18b3d7bebc3f48a5a70e42de1d624cd0c39a1f2630df3a3f86a82c37c0e0cb013242bc669db7b242974d890b7ea69aca321f755d5050e0112a3cb0aceb0957b1a22f90b90e844174ba37124f033036d7d22c0904ac2f227e2ce6f5626db73fc85e9365c47f916a1e986aa9f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccf28f58808e4b1b787594600a8309377c5b2bd7ab444b26f731e88c5df4e73c0b7407be4b3d65a1046df469d7eb211e5797ef2397b8f045e25d8c11d2d608df124d785b23db28d9a748181fa8095efa7bbb144d8857a26bd8a909f39ae6ba719f6c8ae469c9af59f450682f2d274566c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h373e3cfdd3885d17f625925d2d0a0465a54bf83d9da322283a472bced235d8af6502c288ff3f85a796a16b76920fed83a902522ecbf886b3c280d63f8219d043e21bc6721a52df5f126e591fd183f0822a332fd38c83599f710b688999cfc98544acb94358b833e2907c484223bf80e29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fe494be2636b276a164aa62e3455fd55a628c65727aaa1c5acf06c0b12d8707b20658c76b1094df11e2485461a05117d946f4fc2a4058cd5777bedc80685f7c399d290a973f07348b8c462439fccee6a55942c5eacdac8b2c7ee01ac239f1f2db9184dd6b87c6565aaf7663e73f85623;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc840cb2f6c0d5e7bc62b40bb6685f99316a18ea1d0cee86c55c71bf3317d6f88c780753108fc20ab8235542de24f7a1c54aed5c6c414466ecc56c518c656e9b127da05a220dd65f98fe41828c5361181cbb1c232bd1e91dced9180bf1d204d115d3f123bef3ea22aaf6a3f3bce20b583f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5974cea0e73dab51a60896126b8c13ca0614bf648fff371049d0408a7034438d6e5007c189061dad67e94d79942a18f4f60df42f2a09df2920eaba0efeaf16ff0665d07520845ce4f14f89b32c6b98607b9462f27841d39255694e909dfe3f034f89e2301d4bea9d878e53bee2dd62c80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb64c7c80b5db0648724209a0629ac28fcc77bb0505f070d10b844fa0f0ae65939d48f568ba5c8d03cc00300dcf0f750edadbb7827d7882dd1bb4caf3ea9f2645c715e9f9d78ca70da41e5c9eaeaeca9871e6d9ff3b7dd6c6145c34333d60399382c0ad98876368caba25655b797392ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c200cb2ca928e6fe1d88ecdc3e5edd22e3c3ea3a9eb769aac9bc2a944d935e7edb879313904da310faebfe92597894ce72a5a5ad7d87ac3e57e01803a84c20a4d4ae76762df068f1c3d673bc436934b44f68893f33dacec0ba3efaf004c45f706e1f24416d4e685ee49efaa2733c81a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he38eb83703af1d6d699f44231aeabbc8dfa217c811669e61608d1b523261c438f6f583a2ab4265e4c6ce40249a88c1f573c6333296b6a13ec5d8b3c2da162b97e1bd298870edb8de04617ace503363e0b2ebd14bfe69a066799bf9743edcfc2f2ea6260c8a15d3237e721f61f9626420;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf37ef3048456532a49e2310a20acf6062bfc57d238e63761ac2ddedeab2b3a945c24137785ce331ca91a33e9fc8b3338d21afa4f507c85157fbf9ec09bd369015eaab5e9e6b60b01c1021606f5080d07c637fa2ec5d9fc2a5c06387ffb6abed2296166a13865efdd2da7d38582fca354f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fd65ade3df9ca952d0f62525e623692d1132e3f3bd55f6efccd163de47ff1d6e6d11225f9e7333577e485b636f31682da9c7fa59748f61358af1b7cb02fee83503d2f23cf87aeedb3cb7ec1bba3941235e93b85fe5ddeebb2cf66ad984dc67d82ae95eab1a2bc1646cd2f25c9b3395f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d2e64c5f70c37650e79d49f2b26f128609b4543512f4f2d6046e575b85cb56c85ee21d29742a26b293bd09729e2dfed09dfede972f7755284823edde61419ec95c3652e0cc47529e5cb563d7306a58d4da67cac6764d90549de91f6000cd6e9205b05583760af8edeaea23254dbdf5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70c1e6783b62a2b56e6543069d45aadac89503eb64fded0f75d8e83c0928471ee1adc9d51f72b7ae8017c0b54430188fbaa3caf84de9eb5bbd6abd1227eb5de9c219133d137e3c6bb61c0e9b69463c01ff8bbb1feb8883ad1d0925f4beb9e6bf5774facaec730d11eb0d99c53af3e88c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcab796b4a13a47b5a8d2ed4a41f1e3b6e8d451dc6208646f1370a53bcd4256963986121377340986c9c6488c02657d7edcdc7f3499167bc660ec7370302161c44b72c94cbacd99ab978fc672136c99ad7e3372db6ed616a56014ed4f331f8b1b989d67b21bd5ea0ec7f5c4eed0020f47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h946d610d4184812f0714d817aec7139b5785bb07661afe93ab4a93d027fdbb43036248f3a448bae54cd838f7c0bb65b343d68381febea47c737b1bd62ff223dfe70abc33ac007d9a9a0d88cd8de7923e8fb5b31fb1dda5c10da86948d234b8057e2f6b82a8dcbe8df0daaabf281dfa8d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71b0e8565718fcc8e0d76789a4fb7e483a4e135525da6bb884d9ba2adbd3da3a8e1d3e3c5282e579329db293c11c175ff5bc707e4487d0aae023d51474e6d3c80dcb26088ed8d89175c758869f3545e4519cdbef6186c2460110c8d70a6ebf564bdb62af34f9e63e2624f459b5170b3ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfba2217754f48e3b72d486a77260c3efdbcafe8ed87d67af7f690475f229dcf649b0cf0c9333b7f879f10fc23172681903dd5328fe425098e24efaa18b8557c5d8858230928b6db669c68781121f0f7656325f01119659f936abefc8395f62f215245a9acf63a50a8d32605267c53be3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha49b87ee2af92e18d2cbda322d10a1a5ee2a3161ee91644736df549da0c06b398d6de5cc585d789e97774b62a8dba0f19557e6e63a7ff4845f6f5309da0db6d2a15599c821f91588890a0a5fb6a24e572ead9ad3552a313bff9a82ab85428e52dd1ab4a46ca55376727017f2ca37d429e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bd85da5ded35de0ff2af0a11ce8a48ac367ce55692eb13377ecbf83b56018326e3b89c72faacc7a44613ff335f7730c86cca6c96305f8b96913e56e736c563f66e881888b74dddd4264f094adebc20699883749345a6e267e81f5aaa9d0206196407c0d3544428ca03ac30cedd1570a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c4dc011bd890762c279005928d4e930bae7f9db4221d3b9eb606a80f8daeefea073751638914601fce6e57b9576aadc9668b51da1198cbd7006bc5e0669e5743a9ba19ef79ad4ed63e2996be785894921004dfc7be341e1ee1b4ae90872703763d210e77245059daed8bd9d6dbecf263;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a52f3516314783b041d6dc3d0b264c87905c1700c9b11690f91759abbdb0a1124d57bf8307cae7a6b8d23ca327660ce230daac43ca9f204bbfbef80bc1d33fb14ff0bb2074437acfce1f79ee27eeabd70abd2d456bd5b493fd853a3ca4f60b8986fbae841a83214212556269357940e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ff31c7ec95e6c6472c6c84241321f20257d12fc5a2bceef6240cb00cf9edf665713547461f681f753fee4b1fe38ccbe27c5dacdb246c05ed02797551b43440468ed9437e52361dea1cff23fe19bf19e2cc6ca6bb5263e6821d2067ecaa6a8d8dd89d5bc660cadd5fda518924cf4e3828;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he859099c7cb93001269374b356c69a97f6a231b45f63de36c8825993fbc48834eab50182896f4228ac19389a1a480819786d29ba63f0acbcb2943c4bdb50211ee677f273dca1b96379e1bd06613b0ebad831484c31a564b1811946ed6285ff13ab0399431752a0a0b93571f4b21179b27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93b58881e2fd5a606122886d8af0d051ea8477cf210aed0dd1476b66c4af0503edd41980ab3b65285bfba2ac855abfa635983d2084a25b17e3df1f9b7d3314280d5804f616c184ec11e0b22afd96fb9274ca6f5983f51b8e67d30ca03b31d3a267bfdedb39ff75810dc56b2e6423ee70f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc38d1c2a254b07814d4a38bf6c99324b8d2d2083d67e42ed350cada300ea9b6693059e9bde93db8af193b84c77f4b51384651572ad6b3ec07116fcba2b3135fae1489c43897c16e062703a922b75b1943bbe63a2e4b139796944b4c4fba231e7283f1e58d1d0e5c02f307740ff9262b98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1268b48cd9b9eef112f25cab804cf961cb5818a2d74e3d512d27570aacf481854197e61face38289376b6f65c3507c9069f429826155e5052e01dc9da6f09cc2a37dda53e430e835b3341ddfbefd0221777df50a90f4fb88423bd28ef3b4819cb53892f8bcc1fd0e6273fb2dc23aab14a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5496e00ba2dc21b268533b7da0d6e431440a8b83b91a1baa2a3d2f498f4c5257c94e0257c80b846ce757ab3ddfe71eb485589252c53af8f2f8e3edd698d8c2392946dd66f8774c5ffb843e6b2d2a0dbf2ed4d1c3edf2c9f6c42ae551cdb587fa01f3dbbe9c45ca727bd33e93d42b7f6c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a3b07e5ae5bba571559ded75be481e941a652e093497c15f436387a983cb0925c95569aa224a2643b041f0cfc7d090c02cd6e24e4b2670149e017440285c9c53eb3791f7aa88b0e8507b9a0034066dc6c90857a92010fc6c4d78f9e9ce75d44a2699190f76b6d6532c552af31f6787c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1026e1ad8c9208ca4a548580b276f0afbd5ce3c6d153e416a44950443ca2d4feb8e09b9b8df7c31c1fc4832e8a77c15fe09937af3b0b45a656f560b545f4d277706405959b84e6fe1228fed5fd340fb1dd55a98192c487b909fc7dc8831e4a996157eb5718908cd74bd89468a788e70ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71716dcff6e67e0f212c88085ee6a375eaac5baf2ddee0483abbbe08fde2bbc15044e2ca30b5631d30810ca280949657b6b66256519e2c04aebdb23cea12421469e0ea118fed34a25ba0fdae3af2163c076099f89070800c3c5e316c507ec36990e0cd09eb3ec180ca1eab403de8205e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69a0fec886facb28c00df2e4e26dd40dc5ca690ab6953ba7b799640588e1ebcf925a34e87b4fb598667a463748fe25a976252bc2309560357cab34febb788f1ca5a475cb7feef64b3b27d8316be697c0a0dff128ff185639ccf836fe0d6f9ccfde9f8e3460215a258ff6bb6f9a284dbd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2d8a4744bf4fefba7e7abca237b79bfbf6d6734e05b756f249db7e8cfcfe325c066cd0437ad13300274f71e9aafaa2c3b62419e851c2385d75251d8d1dd19c4b4830e892d5a80b7d29dd02a63ed01f44dd154695fb91cfc0c4a1205595531811a31763f9bb67579cea941dcaa1545c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha25d7f3e725ec5c2054b32a0914f8a9f4ad6a3c3313dbfc62254aea9a8dabb6ea8b46ae6242c951e3c002a263769f7bafd24a9f4d08463cea069b73c2e114b65f07176cbc652fb78505ac01dc362759fd5643b0479d185fe47018e065b9c7d5ae35d3a94bc9a950e5eefa17711db85a40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc97b9d660b9a1e865cedeec022ea86e45071d7c96f5ec9a024b2eb3efc5143b802b9a14ed3fd4b65ab89ce4f7e4ff793110620cf8c3b4c82c5c6437b5b78697ff0b6ab262cd63e56cf495b475321d6d57dd9249f3e2071bb58a75bcd122cad087d21ecf25189f86eb78275cdf1c47fa9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h466499750338949f2cc4347b826f31c434103d5e28131986706f3198fc7f777ef6eeba28fca00787ebf9a0b3077977ef4ecebd8a4e6c6f1340a5aa0c6882de8ae4dc1df6a4b9c9e3c21fc7fc9048eadd7bfdc5b03e254dc3d055f7ec4495209c2316a737982fd17acda0feabb1239c081;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fdf300d7b1b98ee3074f9ec20239b3765db6ae5dc7bca2a8e9fa8394439a922f254d853efbbead8535588052d68d13d476f0d174f4d413329a29a750eaf4442390d0922cc8e31f068c82020fd812407d2448bb04ffcf42c2095e4264fe415941a19615d5ee46ddcd383fe949acb62a60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdad154302e444879c45b1c386a94e4eec4d35a33bc89bc5bc0ee01b2d9ad24753e5f17f45ebff658f032910c5dbe80ee6e4b05ea4179634693f187b621ad22e0f40fb814d31c5cd9d2b148735135aef1f530b64c0d56bb8a40ba14872e5207e1c1d9927153b416e74cc0addf7102cd7b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2a8b4f15aebf0763e41a093192b72deb9d6a2ba222e8c0c7c864fcea54b787396cb3e72bb8b45327227ea9100807fdb47d67e8f92978b6a9764526c3166ffe2639a79b952f430d273582adf55634062e6956db735cf4bb4fdf121d2fd9047d1762ee697aac8390cc264404299aa3c08d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc97a64e3c1f9ad4edcb6176551d33862f0480108dade7cfd13cf12adcf9825880d39e1389d2fdfc5d1677b5213395b415229334d7061fe4cef585ee2c893c6fcfbcf41c2f979c916f7a8943e8fd95a1c42924a417008cf4d9c36f1dc06e62f91af1839214b3c019fa3c3189cb68532113;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e7fd97b310c3b34fe6db4428b24b591941a3c5b876d8557f2e948532fd92d7445858b4f5cb58e0012dc263967811caef4e374c2dce3d731babdaecff2e2ef24c3915fec097dbc5e257648a1a1174bcb8e225342857929376f7e4b20f732459d291f1871be2a9b749c6f02227ce67601e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8339e15c811d6f0804efb9b5733c8e7c9282ef75ff2cc349637355cf28145825ab0c923c679ec4924a31be0da7fed58630a3e9e4d6e6fce2120b18d33244fe5de01c49a61d7d48bf22dbf6b8a652fd3530a73e964c60b74954ebf96ae8c986de54b32d693a3f12ed36c0a8266903628a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h722ce56682b5a6012bacd150921352d647e8dfd386050970dda0c94d5b8e3e2b53144adb7bc08bf07e3860c87b2ca70ca943e56b3d1577bf60cd60c81dd1049d6a99c5629e06c0ba3dc8bc870ae62edd39887235e6f02292f7316b5f00d648fb985b698f9f5474dfeac045b0d09a0dbf5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3cddbb4db777d48f26fc7bfdb66efd8f71256bf3653652ec9e70a22f5eb292b5e20a288f82840a12b44a187a5e6988ddf6938d715dd743f7970e9965d8b504051736cfecb51ff3f3301ef7c987e3d9fb0509b183d0b4dbce679c80938779ec9e59f37aa9b94fd346e07dab264ba71f2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b1cd48a131cd2f68dc6a17f9da1112ee56233becde8b3162c68746f92443fae65cecfad00ced7aa70ce476689d0437e97d3d23733d92f438f9ada812cab0b2e2489aa0bb7f9f0cab569d49eaf4f2ba3a4baf3537761e3e317e48cc7f6e9990b114106e2788e881afa4a14ca34445f225;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4e511757523077e4b3c9f21be9741d351defe9ddc07e5603d8a715e71d022219e5f5024ba032b209ef5614666f4ec2a262e83b3561c967b04cfa09c32b9ac899709e47c53636384c7918b209a1fe2472059643957baa770122e2d5f60710049b94778de0b65b47fd98472c5e566b96b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h435a67190cf99bdad9a4ce7f5faa1bc2733633549e8ef344ba9d2eaae39197fa390c9e311cafa357a60e013a603a8d1f3595d676e930e50da217d94525f9343693a3334cd52fc652a8761d8ceea34656ea0cb3b209bb450eb691c6e5fbb9f19a61d25f2626df5a102baf9428ee2c191d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h923dd1bc997fc36944ac2fe71606ade4a6dba919bfddccbeaf71d8e66f4adaa6dd8811b5cadce2be63ee39967713d3e043f296c24d00fde21cb38e068b870220266dfb19a26aa35981bb265a75c52a5b3ed8214f136c593999cfcff99dc5f7a48f9c886fcb9fe8ae59f92702684d0b284;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42e7fefaaa794ee9d74560c19a8abd160e551f8fb03713e9e554a25f46625e445e28b770059c836bb5e94391832411134952dcd9e4be9ca800a4e0d2c6e45cbd23cab13002944dd1fb20b5dcbda5ca3d0c790d069570e7cf89c34a4d95121bf43b2b48578f6107f17e2d16486df01a984;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b3c3e4cf9af3bd39f11dc3be646f71ea02bd19158cb43ac037cdd71e5b537556a5929a80661fc6734deac1e94b19ca7ef842d1c703ccfe0f2e4ffbcdb4ab8904fe1fda53316b494d231b97870a93e05c891d7818cd99e3de2a61b9e0fac99ae8d1fc39b8052d58686bf89e939c171b8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93e6260cea6c67880a9ee9c7501380defada2b2b9b9046e9a89fd1b22aca2c75eb55ed2dd1f85262d8390edb36bd8cd8978b6b06d82d1f10f66bdec9ea4941464ad1d37fc45e0070b8e36e5cd7119338d30d4aede1f2813a8dc69288fe1caff3d2741a755461e43bb768377bd71ea748b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5c09ed554aaf320124405e1278343f3232073e90f9898665718e6316221362930cd7abce56f80802b64925c96870fe5b64335b3283c9ad7de256b62dea99021bbc5e68677a15bb03a931a9887e4038ad286e426c6c1eddd754315f8f728c00ef2529c926b753d8f05c5fe0c8e722b1dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacd8f45de8dbad7c0df1e3e0cbae68e94eeefdba7d1126fdca2c3e60a9b7c14dc4e3f54a659e742e39db06491052ddf309fe5d9f62a0902022037a7d22a42889b71dd2dc4ff6042b3c00bc69198e943e90aff92e3dae35d49305cc69eae127b769b3b0c0b495f8d6c72395f4a09a02467;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa64bd58ee7c2948477a0f5a24bf4ae8b20c8936ced4a4849209160ab67e96d2edd63f8e3bf3ff1a2438f6ee716163f9c92f0c95b34bda33260dce34a4208abbd7d7185e581ef4cf82d8b42658bad61d94c4c2a79b6b7a9ef3cdbd7ad36b851f5ab1ba89a7ac1d0b74417f306cc36fb39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59c669ef282afeb8e3074055e73bac80ab32a3f289e903d1fe4be569332645513eb811922ebcfc87707647b6dd41baba436450d083cde4541b696b01b6d679b17e4e4c7ccc7b70d092b876eb2c36b974a559529f1facd153729e2c4b3440ea035c118f8d5700de4c4fd588c1834172bc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h659e04616e7dbae71ac0798f7f2bb48a2e76c43353bc929b830ace38b4813f8b802c97e18992d8817e3d3a4d64f43162c11aff34f7277b2bd40b2bb658f4b4a87a8495e0296d33a5577cc5b7422ed0c9e7c782c1a9a9e0fa3bec64b5a7ab6bfffc9f6cb785cd5ada1b298802c3cb609b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83a0368bbc57678273d417b01985739a00416508d5772d656bd09a2f328ee9c1f9b81de22764d7d4ef25ac59a88a078d55a3935dbfa18e77437bd3ba0a329453738e9f6b9b6706e891204212012ed7220f43dea921fd7962e545b174772f9d746c6611c5e3f2b98c061a7335000cd3a02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76ba5efff4eaeb81ccc4909171d4b60f0688592ea4142546b06000b5eb2e044825b11a67bfcc45eb49cbb5caa3179f20ace3e2fb3a70fa5fbafc3670f2a3608251788e46da4f06533e4791def37375c0b4c7ef8c66a8172987b210d6bcdc43b2c567bde7e1c2e094df08c9a7410937573;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb78f1727500c35ad8937f5c41a24e6c878da812c8e87d97797d916e72dc649725beb1f041a38eadd92ba7fa12fa5f68b6a9192ba837059539b8066cd81ed47c3262c98ce8723ba6f90e1ca01a70f2b493298795ce262cb41589ef32d097a327b7cc5297707bbb11769efe9decd12fa450;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eb18d8985048f9be85755bc48ef7a96509b221fe934c191b9706324ea50da899781a4e0dc2d70c52cfd0a73616c46891fcacb3b4dd0ab5d0910c9e6942ac1f250876ff843915308c3e81c021d7c007dd4e568f2eb775901d0b3da692eb359b99ee09696eb6124bfb4fe11b52d5cafe57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he14bc69b016a2bcb3e2dbbc231cbac664acbe0e2044192d37715751b17e34d1da1510413ace5d265394b8971bf495245469dacdd4cffd35e55adffdb0679ff7efc1a67f60f757abe04ed873e95a3d4a29679454a490d3c9b7a36179f2343fc700177d22c7b6f5589c385892c8e4d2d3ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22c33e88b5770c350caba2d0beaa8450675e9eaad0dfd4e1a3ce53626211a7a64a06a8df99903049749233b8045560dcf934a27e876943ef9663c4a93cdbc821fdf17e046c98d7dabc7b607d692d721e80d9e8904ea30ac4d1347204feb75314bf0af6b29d6d41a1835224be8c576313a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88cc93bc14e58ad08ade9700c558e3128cde3e33ba8a67d030e1a68e8c33e100ca9d68fc2c94ab6b53dbf76eac4ed65a4ee523931a08dfca5a86134605b0eea2be6e6a85710b248397838c48d5d33000d51e456bb4312b758fafc0cda07b5fb203f2e0168e40ff976792e1f4052b364c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3383811f06149b6e4984de86e1ca22af98e20a4fd154aff39cf8146a31c226c84927cfeb2df2507bf95d94f9de3d2eb2a49c8e8de932c3f8d1e8c6a93d7427e483d325dd00a9112f4c732cb32ee6afdee505e94382822c642e90c8b6cae2e2b5b0293e7e402a45345b5f1a2273f239ff6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbf5964823e79d0b581cae691aea2fda6ce910e21662336fe8d39761a7614a309d746671ef4d2dde6f4443a61add4bdbdfab6e2cfc2864fabe130a5c134f2fb6eb0a0366bc9f8dd118a76ef8b0438c88a32b8682b9f23f4e92ae21fd707633adf14b02d3bb1ccc048aa1554b43dd9f1fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89b9e20233ddcef6cbb2dc4d2c96d2937ea53b236232e6d512ea85090b4d0830a11db79d6f77f41e2d4d8e43fba4930168a9e4dc1965b87c49bf90ee97c90a0308525f3a9a43e0fe824df31a96f6e736ecfc197c928207ae878237ff1632454a98877772affb66bbb862c731122e3707c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha17ba281230c2c8ab1d43646165d3ce6ae38c72a678126b1df58a29ae340dfccf7d2df1adfc563c5a6ca9e9bf7a2c7f0118e576bb3e9eaba775ae32931f6dffbad669de570f53446918e6261c7f89e854be48ef33d579ce5049669e6c998f856419b17f3f838eadeaffb43b0a1bd6c7f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c678f33a1e1140cb955ec14d9de060f614b7a30e48aea18a72f22fe9f0b2e791668ac215d75ce1bd1c6998bb56f853d3c420670e5bee41c88eb94251d24e49233511d50974a5bea46d4e49ee7193a6243cb727117b16d5f54475c4044317fe6ef555f256b6e6aa687ac55efc9d6d447b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64ada8d9641ed2717477cc4355a222a3286b0db295a550537d4a1f6a41f59764ea13a23df3c5f7312d9ec32631f4f23bc16fa20b3093b218d5d56117caefbcae0a618e0cd289bf3cf3e89cba80ce9cbd07795c2a8d666e156217d08b22a3b0ca594cc740b4556bab263e3a3b5e621425;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a356d2bafcdec9e039ed5a8af4aecfe4d882877ecaed07e67b710b2921ce15b3e1ed67af33c2707d3b67d206ebcbb174f2e7bb6f2d2c81b2488e8f252e66e7faab4da5346344d78dd3e1fd069ef425174d542e309c4d420bd5d182b4156419dd18f58ce59c0c097c0639d70e175d861e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5bae85434cf0031a8a886d94d1751859ad93a29efe20a7fe9de77977424ca477f181c2cb06b870664626c4698954fb818c0a0d24fd4e2815e066b005cf5c36d8701565cd7c19d3c37cc1be3b9a92a65c7c96c894c02bf8de543cfe006bb34796cffd9bdfd309d54cb32f3d767e7d9207;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h771e88720ebfb5ceb9ed7b851aac157e27de766e93f15874980da3950502dbce28ee7d9b3fd0f063a8742f06c9cb5ef947e2d7848b2a22f3bd426db864eb06a98347ad5d23a8a45023aaffe63e683b9553482a73c141238c58f03c220dabd470b96ef5f867d73545e94b81088b76a8382;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf10a0c9b8661ebacf523d3862f092646390733d659b32837c8dabddc88724f9e4617df26589883dfa0b1caa1b4765e1f7de278e89d4943d61c40ced295ed2766a12c34dd1b84b2e49c6a338fa512fc73c05853b8b15633953b4728601e32a330ab13008f0f2d78fb44f81a09fb009d1a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28138abc4b8cd2182cbcf635154f0f722d86b12c53b5723af35312b82f6e571d3117327ca43f87d2bae68a695fa0999aece1273a21e3af6937b2891b2c62d75a3bb764c07a5c4bcd8a6cf1d23c8783d6a9d7149007f38a1015190419fdc746c1fbf51ccb7012993fe87a9de81c5811c23;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc728c5d05d800b5f7752265f0164376b3e1eedb85e4f76619604b1735e95558cab9e1d5b8ff299ee83fb182a4030fa83834331b131af8e87583464ccfd15431f6469cf829657f4902e875c79ed2df90083e8809247f83abdd25db943e3c6e1e2159cb1c3197f0cb856727a46c9b66815f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75317e441eb3ffb1f57fa2328410868a659635b5790f7baa5389e5b301f79cca3c6693fbf3b1a5e5cba1a97c1adcdbd815b292d7bf6d6cd332cd55bc91f9edc3cfbef745aec6e2909da7b131983950814f2017f5850a9993009c266129f0a09b867a06bc167d2dd014f9ba58c3037384f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf156582b8e8d9664136acf6f9067f266f8d85173018020fc3f8b50a451b8c3d14b2aced93ec18ede8ba4dd793eed48bf4b39f99e17e52891c3e3dfcf1d20226a733bf2df19f40eeb8dde1397b3abccda63da41206dda5d455ff9df5a4d7a7cc920db792b3fde1d62729a46ecd20718d55;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28684663bfb362f0c5395825d3acaadff0105f5d5e82ef2938d6e91b34908ffe71e6b5b9741c251a502c9e5a1d74435db165e524e03bed7b27dc1ab6406816b84e883c9c14ea282c2858f04c8f34c8a33c5c9f65ea6e3ff36e3c3f7c66f1f2cce00df4954923542155db8d2aa9e93c925;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha00e66d8218afdf515f979c43c275375481b5c1c7e2ed4de17064346fbe8a049d0fcbb5e7d23b760e281f54b22732058a205034003e82e9007ffc82666babc78a460b31959acf72e355bcbbfc4e37c0a93149adde44fb52deb437ff431a8fa066eb0373de1f8861433729f07ba06721db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56863f31f6d4101bbb9a4b8882d3f70541106f9c7bb0eb5ae536c6c16966930b3a18c4146da76218b8b527867763cc75015810d92b550f83fa499dac3c62ccdf3b16069d1d86a486343c1b51eb2c3ab7a21d2fbca55222593f7b1ca7d7165f48feda8df7cf6ed6f5d2502d3de24579c3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedbb57277598e962c97aabf068428f35aa7563789671065a2c32871edc95fd1c3c9e58638f15a2a1f07bc857c57bcea27f8c2a19359755be91394587a4a73ca8833f97d9a5704e5ed146fb2fbeb3d2b7739cadb9fa0d5fe5e3ea46f52f462299f1c3cf76b4e26cdb74a0f254ba36564be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21b2251ac93335257411c5ae6aa45b0317497e37d8350f1a6c2176545fc1236fd51f80369441e86f373be6c0af5480feb5703937be20656ad57495c2d0d0fadf421dd11a5c6b159b7f699e24640634b523e6081e3c91fa571e1ad5ec2a1cf10709e005db20382d4e79014acff56be65fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacd4f8c29466c4348fc16d35894a28d79cf77baf9fcc136bb294057590b41fe84617555a4da219cb3cbeb84325ec89aa4e8dac2fc995727627d588b3f4b0cf10701d276f951119a6cd7c4e16a89ec2c9ff8da6e27dbdea30a8d642dad84f139d17c3bb903948bb56e2e9d70712d7bb500;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15589310c0db92296029ccf3ba96e0968ff72fe0c3af04d6c338af627a9813aef6a91b08ede6c2648769ffa08c07becd5cdba4052a9720ac3bac66c22e99c345c402107bca513082671af0f4267329bd10838b1f9cbcb8256a3abc48810511e455b8f6382d399b2d8f4495ddc1862b70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc883641b7b3c4afc1fdd10af03b65c07b11cdf4e5a556414f62667f82a97f6ea47a93ad7c3f1b60c44c5dba424c4ecbc17389eb53ba129319ac3730999bb82bb312a28efa4c1398c11f184292b37dc31cc03703500eb5e35ccd0b36478436ee750a5e41d7cee6adbbbe73a65b4e9a1401;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8e53a2fc2c6acf667233c38cf530758aa0763dd408e51ae04c4142ba5d7499ce60f8ca401fa0363d093d62ea07234651fbb91925004f424e3b670f98f9315a7c55f58ab3547efcffc8ebdd57715fe0b322a667f4269b4eab1682fe3074b4061cad70b0bc7315d4e82597cb85a158f9fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6aedc325db045ede895f357fa1d1ac314893ef506a14aaa724b8532cace91a44a08313287e1847fc6e0b57a6859af340559fa3811e949c1cf40dd8463ecf2207fd236ec06b9ec5f28bb9e5c18333050a7d2825d1fc23677dc9670b82e4f039ef997a3d4979ea736075160f4126c818b93;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67c6dcbecc399b93fe8c373281c0857c007bc65a9ee47c328d1675b1888709ad132f5def620b139b177a55e34a4af353919463c1bbc610f2be95e21250250628e6e9e3c8a0608cc2acfe192d3867a44396732c1c5598815c69f1853f56d2af9e5f31ae204cdb05ad0906aab34854f9077;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he33c6ce67ed317b08e9200c520cb5e3cb66d061d86a6bc123d304e47d6375ff9ecb894e52c1f3153ffa64e06abf88555a44780f41b91d153c3c1676da7b68a42048ee1dede6a38af2051b8f0e7c2f7aae0937a09b756a3cb16557ff63978e5fb065254429229f93975ed9e4ecc798b0f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29ae71288109c29dfaf2972a30926dda8052595266c3db92f6b0883b4971b3fb429dd4cdc77c9aa55ff57473698f4bf99c787e86aca1f750788137a282bf1ecb59339ffb25f34477d7d2b271255c3f066ecf2cee5b9f3312e979b13baf937ce80425dfd977b3af4f94586100fb18a6b31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h707f002a98857ad591d9975b5f9ba2b6db39ced561a1ede916cedd2710e472ba6cd38a0f0a789407f32ef859e5845c58d0246ef56f67f7998a658d771fe31dbc8e3d31f0d8111ad06c08c6a0fa4ec34f6be935e591a69ebd2c4d11eb788324d182c4bb975cfd3d170894ff9edd23a5d48;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc4b46ab29725e3675f73db1c65bc5f7643ffff5035f0be947f3e0c97f6feb1defe58dd2d8db073b01d69ca2186ba97d7c49831817fd0677ad68c995fc7a2c017946b1bb7628d535ff0f1be604f3c34df0a00d630c807551073e2cd4f65cd093abc16121031afaa869766fd2c7635bae2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9738542a3e2d6d4db836924c6f79264cdb93bf2db35f59b0c057dc716ab554e8afc04ab684c889704af8f8f08d651d99293b8f0dbacc7e669a910879f368202ceac0190875f51ae106458ebe36711f46a7658ef387521f12aa25eb2330062c89e6d5947e17999c8380332ef544dd3d78a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92d835d6cd8d3932bdde85603deba5672427faa76ce4d66f1d838b952ffd2696efbca13fe6e84cd7bb54dff0ea39e9af4d6cffc9e1206313a2a080058d645b0326b12c747b25dfbb83f63604c1fda89847cd046bbd4b486756a75197e166ba196f6f9d1a17156869dbfebb733996416fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2218b237917e6784c8daf0788106af7df3450089fceead64cac75aa70ed23737448505ad62c34452536d0a226fa19c06a00b2c48815ff89a8bc52cb3cf79ba9e99bfaa09e589eebaa161704df3424ef1a194d9119f707ef97d7b0b7d4990e3a7a97b2c42ff0d496e945063ff7866d2520;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3a98b38045b56b615ea220fefa6a00ead7f3a673b6deddaf87e581d3e10381c71ac59c088277849fc1b2f9fc8b82bd77538b7eaa7b95ce5724bf8a97374515c736ed11456d9f655c8558cd03fbb32856a97d3914876275df075861d3921f26a25f4fea754fb4f9292cc15949586479a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb743be25e500849021b861266634e4b0d1a2cf516cc29a5e059ee8ed0225624444ee0f179a1f13f56a15f11a6d236ccbead522ab57dcbc727d0332f5fe4458486858fd0b79510be7070d604ecde26a0b34da39c17ca32db55e045cafdb8df5f33b95753489f9cfb37c7b0c1f14a6cf58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cf03cdabcb09c9fcb25ea366bc86f0fe114b8accb4d440f35f9037d5f4efcb8de1a4acd4b0caa5594bb9cef843d2cb6a8fe085061713ad03bed8c854b949fbe210326f5ea5f4f520019cc0e53ccb27d36e6b433a7fda5167d4de209e9ba4463ab92de3fce1153761080417bc1a4bfca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79b2a89d4abae6ceef4df2472da878a32e3031c970e576f7af1579efe93fb97999e129b689db8b80ed9d0d42ffc9e5e978d76302cdde0f6f91f7588b6124cab7b71eaafac64f7c37c1525f0ced5c094167f24a8c86edc6e1daad37a4e16d3c3d5893ffb446c11009f05885b3db6ffff51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31440cee77ac9cc3f9275c98843f7599e3703e751dfa2e1c964ba8246cbfbd1e3abd0220f453e4dc1f25c6f0285d92f4ae87b4864bad7c9c8ff4aca9f26c4d186b6bcf0fcc6c9858268dce95fe284c51e26c2b91a5ac2e01a1568d5d83e3302df9daa51f024bad42f636090056eff6a75;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4f61eb6263ce1f97571cfc67e4148420fb40deeb8e19ae14bb9e95fd050caf6dbbda6ae82ab917a5a35c2aebeeaacc2fb9ebdbe00f2f6ea96a281c74eced52ed0fb96339f30ea6a1e7b539b52b6b20377ec2375c0f4f62b2acd17a3ace03f0c4eb0ff7186bc0d8b2428b6830106fb25e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h305cf058afb71f7b02f2510f35a80e2784776aeb8b98ff6cc7408eb0f5af2fed972a881bd5026c0ce5a4179cd28ed26aca9f14bc71d82f8caaed5ed9036d79360a4153525d88ac0f0252dead7900183f8eba81eb0366bd29722b7bd62771b1b42459a2fe873786df92ed8153f35deec6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4740f1b27865a9eb24fb15abf77d17dfb40b856d39be8fcb0db700bf2a2cb18ac6411953fbd95382935c9730af77417eae9d48e05e43a65c210521c59c4e49d760f69fbcd805a69caa48fb2caf89307ff2435516faf09d0a873661ae2913bc7514a142c0130cf5333596a7a0886e5a3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb2e2bc27c5f08ce6a3619104366e23f8117bddda8602c77ff4d13ebafdc98320cd7bb7fbeeec83acd67ab0b81856c49d73bcf76e13db37fd792e88103f71a4e1b03488be0f284814b9db95fb4aad1fcd4005ebc94621ba2beec766d8ec7edbc2d5e54ab024dd25ba0fd8c44b4a429589;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ab7041b69a3467bca7a7c4f83666c3b407a1e93ae17637a2d131589214dab3e50fe6750d354b9812546f3a9908cb46ce8b3fc4edc16ecca91c178626ac429b5845cd58e2422c86669a5ccba9f3f751f89c352be80be4b23b521a4e1165557ddc7b25f62c285a826544354ae6ea6cce84;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49e4ebef09044d0b0afd400ff13f44eb62be989fcd65d5ac92a40de20ec51c63ec584d88cec9190e3cb7e1ff0b1290d2d3fd7fd55da3b9c8cb646b3089a09e42b938eb75850f0756035436e40a4af05e961d3740b43d9da6e5b88d4d70d981181db74f682a9c0224b772defc7744af8a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd82b8c28a6d69d668f247f09fff13a6fb672843354f8c0fb0e36b864f0db52ce780aad034f834561954bfe2d8cbdeac581a5721e51bd780d5a5b99f36b8ecfc30907c3f4d5ecc6a39741a1742d0ec892db33770b4989e44770493bcc12826a99f38c481057650a45a40de3214d14def12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31d8a0abd6de557af4ba5196c0b1c5378590c5d1a2af6a870ba207f3faf216c658ee3982335d8f6a3bdbb84e8245699efd3d97746f65e1dec310ccaeb4e8e057725dce79cac9b033f8805a9eecaf507f2f188f5a1ce46bcf2af802a51b42134309b5b2d7b7ff261cf274984b36b7fbc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2ba9d0a27ce1f27de1833240fcbac95e0475e3b52008929d9db09ab2a4cb6f3e428152a782f8adb1bc0193dab9f2f7a01d41438151b8e5e2fa3fdf1a40729e9b7a7c680c09188e60ec776a67ba7f25e3ffc1cdc4a8f700b32d42fcfea89083cea127355ee6c54f8f9f77c223b303d9ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ebf4e6afee944e28c034915f3154882ce00fedfb1e0873415b0e32f48b00f8e83117f48407c61f41f553fcd1d8820492698114d73a38595ecc6a14863dc4c85e5bdfa60d0a2b14402315aa86efadc7db874a3ea135fca01df441e12e4b5f9f814cf8a904faab34ff3fa31c52ab8e9dc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8f544b3ee2d9d856b3ef953ee135686fabca422c1859a00195a348d459a8b4d4dbb48bdffa105b424296dc5f5a4d2ca406728674e25fe87b4dbf03025093fe4d4de0e514c7b4ebe69121818a7b8df2d88ad94fa89f72b8bbebfcfbd06ed11fd2bbc6c0ca4a5f3b052cad4822e2a78f64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78f48aea2357dfb9974425fcef26b95f1801c8cb5a63a2dfc77d8a01106e69e62e1efe98593e78c6ff02aeaddc49c817236027324c73d09b48bae209a33876c77b08f6b5188949de77e0ec68c34d54a8028b7537b619e832ff60216d7c43679580921e01f1fa097c54cc473f077743b77;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85c06468d82253efe7c0aa91326743e420c8645568e2216db69cc2972c39473336304e1c445995ff20245b3b30395685a1dae2d31fe2ceafd69f4d8fef5b996573998d7e55e15466f7c645763ec14adcfd6617ac14fb9e2d71cca8bcb1be515d3df5bb088e83bfd214fbeb71481228a08;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he53778d1e7cd2d31093edbf936e5088af94f75406de61764d041046a970b735fb7a8c159ec29aff9401cfcfde9c761fac87c734418269b70221abdfe208d41d8dbcda9e3951585351323a1f77aa4c15aaffc9f0ded68109cbb046a10be217f83411f77c2bfa7050d9f82f1b0f0ec49860;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e93719aace1f1a53e065ca67361fbfb79ff349f6e4d79c6fef5a72b3c86fe3d684fd4edbba3bae1e8154cad2bf536b114f7d52bdd6197ebbc5428bd7e5446f05aafc7a0a8f681562ed0d4e00c9fc2f203115e8695f62e604160da202d1a5464a9508619616bbb7c330a5f06af8f89d95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85ea39ff268568bef3f8dc2d5d24189a55d426950103494ba4f28e506256777dc14af61f824be878cf9d534ba21cd6425b639233e558404051b197dc8f65b657b96b22632130c81fde4e98cc12c4b85c69445ced1967cff9bc5e42b6e0fe9f89cc58da88793a4eeb04c70e326252d19ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfecd55b7f916f11e0f35d6e7e947ed9fc38847555a9c02d9533f5c15b2b17d39349fa58043cb22a3bb9714ee9a2d220e77dcd73c9f0775afeb7f949263aba2ab7c6bc9bca6e5814e56b71600a82ac631c3b2b794d4fe1e8471892ecc5e8c1c0204ab5f4ff6a93f29b50d13ca953dcbd65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb440e487ab26a03aa533b8633a68adb36082f94e418a3f145cc9c73e63377aec9a302860cd42b63ceadf54bc197edeb6ee43382dc26edeee34d41a486f1a7e27e4114e16bb0db94a418234861ed6239326cedea3d536f4eb7a823e1022832440c3086d502283b675fd4795b5984ad5643;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33b0462e7320c0b6de87480ca0adebf458729905cefa5180296088dbf361a044d44a351e6b12c3fac7eb7aec98aecca19cccd88f27bd6d517c2df04e069bc5c1c2551a2a582965dce2a5d68ee48ea3b1c153afa219fc1b132f35aa68b8e118b1f066d2e6db953e96007879796768089b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha70bd1952129eb4f73b0470a0de28a9dbd383d8b6589de6e71897cee826841696ff33f4cd03334f55120f9c324718d595279088ee7b23d44cb3a5a0579fbd1c58375e15bc9d6ad24800cd657802e09c7da2638a7d234ee931ca3f62a169c0a25aa415fd4f92425d816d5912edaa2e06fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bd7cceb21c3b37b7cdc90cd859225bf097c59d57d1170584d05ddaadd17889c85df8311f124b863e73d4c18c0057b20a088f122c738fa731de9f7454491f044bc0682dd8b741603e0f95e993664968ae2cc6c08671356540cc284a202d259d448a91b9c6ee4ccb7ac01ca971c5d17fb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb3a57568df3a3ad30b666834b6353971df7cadf2c5e1b7a9d486d96ddb9a3043f2935c03358d8771274d3bf7e86fa4507ab2c6acc572868e700a0590fae58dfe2ae8e2707d1d088ecc6ee3c4e0d65b231747fa7446ce1b2d6be62795bc1dcd5e21a9772dd62e345b2a0de440dd8588e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dd50ac6aa9b95486848e4e1c4f7582f8a73c39ba2b0be13f014bb34d496a86b8f8373d9f62bf9faf09d35a81c8e7bccf4f5aa3ddb53d60de914d05865a35e5b3c9f02515b94b73d1789314523bcfb8ee0f1c8eed781e43d8ad0186c052a9de44170061d6681f5e50895fcc6769b5193b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3983f76bc56cdb4b544967046ae6537455b21d7ef3d51d3326126559e33cc48ec65507edc349a84692f2666410151363a185c713a35f75e05a0bd7f28c820ecb45a94b3306e31078721e4c03a3c6d71430e6f16a28afd81a76aee1e221f477c62b01a1ac53efafcc6de3e16c86dc6f0e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ede816cc3260331f3f7f7039dec564e677d37589e21a9b6ecd412d96541ecd93b1e5b025a314288b54b14c475e3b0c68b512e1f11057d6bced313ef1f49922911f41fb26e2415bd45011192a46884ba621b2f597f1d0c9518b80dbf330427ee8ee879691480b55963f62edf70eee5caf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h740a1775a11e693d95c6d79cb92768c47cdb865cd36dded85153dfc55d251ce813d8c9d62948846df9a9067236922f34811d6bb535cbe20b089752e053148e98ac6003b535f6234f5248c08147401f0c789088fec17ac792be07ab456f177549b3e35d741e1538214079b5b0c7e641a38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae8a8afa4178537d3a03b503690a4fc729e72c643b749e6241f13362411ab079601648676309ad05d6abd30f0393ae5534ebe1727eebf73f742cc0dd7fb7196499a9b97ed198662336f6ac6b98a55d495c941aba7d54e728be0a219a4a1b6fba62c5ad82812d4a751851dbdead3370273;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf62741a0d349cd5598c37bbfa0dbef8c8f2d5b05ed955901ac12974cf3347e63459bae58455d476a631128fd864c46d30b450fbbf67cb73b6e8d501923370d17b51b7bb61385427239f615babfebb2fd84fe375b66d6b425f4a5fd51f8cd61305caef39c47808e5a32de3dd5f2306e4a6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha75eb020c7440894833d65a99535465e12ffc998cd758d827ef8c31929beced5f07b9fba90606d28d567c8ab68b6470ab941b7c0de88deb8790e5469a12602ccfa0464b6cdd58a36469ecd0a9c98f1660bf5c3e8bd20cef2048b36c3be5475832ccd16e52b5c38cd6a3fc697750746482;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h278de1fb05b435e1ad4727bd7a7af535984e5c18af116f4d8abf31eb9a183abb9c9214734f9abda71a89fdee35d905d57a702098e818f1d49c2131dd25dde6bc0cf9feea7dfc6714bb921f60e1fa80620030a3417f1ce4885057a629e24244696c13fe76a9750352f24282c137616699f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h453147491e077556ad3df60221a2a815e5fe62a6027330140878778a661e0f2c8808d1b52d6c9ca6e3e773d4db75c07a320bce3800d9919401739d0357460d2dbeadec09848b56979ae2cda9e085264e129533a9e194369e534f70be5763267b7ded08f789312127ef7bc1e9fe401f576;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2a48c211c1cb67990345ae41b617f33cfb3a379c015a665692a63ff7b879fce44dde28fbed497feb1cf4d0eb048d46c1e4f89c6edd149ba6903788916f76dec66a332753930ae4fa685b815865dc9b11567d69a95af7d0ccbf34e36448fcee9c9ad7bd2f9de57c7dc59a2fb9b4b6ed7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h174d9306a24f5efdcef50b6c9cdfb317530b0ff95ce93880e6fec62832d05244850ba7a71641c073646037e578482ae47ee5e1fc8898d8b549b981bcf13f8bae710dcd3505d66cd676fa58f7ad4658b507722f277c7fa6b9633088be4874b8d8e9e32fd01ea5875375b15cb5512394b01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7315c692e03ff8c0d4c8192516666532fe0cc216ba127d9a92b9933ba928b44582e29eafd52345b3f53565eeb737214ce566ccbe57f54532bfb25cec36ac9344b63e253b699796d168df7d0d186ae83cf1f3b178c0c6b43041e70b61fb8f4f4619b337344065c7e71fd87bc582487e891;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha92d70c87671c419e13e1c6f842a883c9c04076d4f176613a5a96c780f16fcf6aad79d148bba8a582d1caf3790490441b7d2a41d1c3e44e0bae110d950644624758d5d05ba2125393e0baa35629cb484b8d4bc3a5e9b1578524247339d308d5604133dc19530fc22aced214d8f6ba3f37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4922be34c843785e9b9c8789f1b419ccb1701b3a24f342ce6058569b5c45712a2b4c12fffcac5529ef2757c9773b3448d12958abc0e36530646247089d85e55b26fb5f70251c0acc62d5a428879bbcd07f97753dad376de1f8754b77d97b119c8fa37a46b0b647abe596db9c516e5ac90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd96a625e68515642e7ea31971b18f37d949b2b259fd4beea6cef8138c31677c2a684b63c94631dfd064146cdbdb065a8b5b09f0be56d68a0204cb20a985c8882ddd46c093a5a8cfb81594fd640b110172cf3259c05ff0d372d093e762195ab05d07e6ee97b8e3b457800a3866ad4621d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha018e48c247f858b31de41e09c61906df233759c1cb8c880ab91446f90cb1a3dcd880bebd69f54385114bbf3475adcb15f5567a5aab5b8e839fee01c9ffe0463cf2de25567733aba69b335644d5cec5d8d5740cfbfd7f692abb82a7926d865b013c179cc4046fa9588a1910849ab55457;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc9d0dff326d9c1435081ea5b4f852a8934e60a806f6f1a6d1dcccf96831dd0b770fb7a913cff2759b5b67f4a1a42695cbed258567cb1cffa6e28f8f4263e30e808f04c48646b7e745cf7ee84651c7a72d7da893b86d79b652a2831a8f55e7936214821b1bf6457f65f48db0bce5d18d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda5ead7061b01f8f58f84c7ee9a51e598c9628177cef912dda2a8c11862e9cc7b857f03b284cf0db4f95c0f4785bc681a4bc7e41229631c8b7ca772cf983175079a34a2f00a340747ce637cbb70ddd08d8cd2762a88bd6ab68e5e41490ccfb427fc418d286ffc78cb2206fe2610d6d3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a5152fa1b2f88511cba1ca862365c0f7e1989d85b61ef09ddb4f0870f04d3de815beb1f2004f904eafbbbc31149d8d429ea1458b9fe8e0949d5c5b96a8857422b3a6cc31846a0cae95dcfab2a1b22144b414fae18b67bb06735b6ccacd432947edb7148812b8e122d5545f427948d69c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4953923e84b5a6155a8613cd6945ba7f67e2ab3a7d06d0ad07690156db1fa71c55db872be4364acad5546ccdca071537387b93f271f88e7412f4ae8d24603db63fc38de5dd5b5a5e232cace18da26d372c06b62aae13671ab2d72c4893eb518466e0066e58c67d2bca37c965819e99227;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he66aa5b9fae5e324c7328d3d15f637c2bf04164ab83e4d40bff3189be2e87f912e97271fd43050f36ccdefed3a2bb27eb5aefe986de9359b431fcc8bc10b24e6168d624c826ab37c39f1c00a8b8e4c32d7696babe0efea9a320a3eb00408f80ead0d07a3ea7f03e4b89341d6ba7910555;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7938ea2d36ebfb1c32b02d24205f7453abe8d0c83873028275ef8881521df9b3aa26743cd9af2eea1adec9b2a3ed565c9ed9057851d76dd4d57873914c67f9bccc649c40b7f4a53d4d3fcd4ec056111f0892f362372270546f65b96f9f64a97a11ed1df09174361485024a3ee27beaddb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f40a30e7276e55a5a962ae2104c931fd7e99d1a4b59e9681e3659bd1ea53a4e2b0ce3d512d5285880c6e9439f318ce5612f5195b4632e384199adec484634a45e47caa9acc59a06835bc9332a5f6a0311c63053e65a4295bc024354c19528edaafcb758831891cf83cb2e23621fd484e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8ce888418082ab0b773a25eacf627997757f9dd0dc95ae7145646733dacff13a57cde8bfd9797fd090b51e0aea68fc2daa138b9dc0b8b93cbf25ef5bcc0dada48b64678d3ef3f60a7cc9c31564aa399b08cbbf847cd57f0c60ec81e65b549191b505516d839e079b8165fdcf23062458;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f33941f14d3a1db9df92fd5ae682775f623495c8fd2a9a262492eda52b2d279842a95233ac02eda432e771e9616a6dafd776b3001b459d16756a18aed70e7ccb8db5c9be9d641b00a7f9c94bf085f952ca2408a717ece93cd79140d3932c509ff4222815f269acc1508cfb532c31e224;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a8af4465adacb163a8778971fc6102c540fc7402794940a14a943333b51c0f561b2fbbf9f014869ac2419aab8888a8f5474cc9e116be906871219f9d050270bfd76e1536532d12e41095a33be96dd495d86d016b556ff0b16f6f51b14aa3f946cf742e23b9011f856bbff773b0496bef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cf5ff5ec4c952226851cb1ed99054ae19ae4140bacd44e58ed3bccb9ad538c1d4c11cd3ef818f12dc1416aefd7d744e2ae6891cb1dba67eafa7c4fcb7d29d9f2ea43ac560f6912a9630b68bf7334e7ed815b142eb3def610baf8c114d9b0434e98808ffe568ccb83f9ef51eb9fd51084;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cf586a4b832d98dac1e349f8d39118b2557ec07aeff944b73c2d2b42eed9370adcfb19426010a855a735d8c8b2d9698cf89552ac6697bbf38df8f2fb06e8a522d30afc4480eabfec22cae2c1dc2b0352e0951b0612582619cebb04fd61416455ffb698b29c85cf96ef88c65cdc2317a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82fd21d5d8bcee4a89a5bbd7f6afeb8b386bdca19ddb17b1f5a1e8256c3256a3ed919bdbe00738ac24c7357ff516e50d2fcece92c5c547018c9b765a7bc4882f3d9017c7cdce593a75efd752324bea42278419b66f3c8413daf6af21e4dc2fb60427c3776924adb5cb3f5646703e4e398;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87ddf2a8f5f31ae6ac3a949b85782839039a31743b891ff6cd05c2ba47e179fa18e55b34cd751550624264f0928ab1945ea3dff2ddb919ccd65c9b58a85c3331b545d7df51c42b133498c6433f1ee33bec56887166af067fe71b9294377aba251ae1f139aa63c8d8e959934d3fc1606aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d8a4fd01858bf9e17267657d697f18c189c636538e299d18092e2c7b8868c231f04adff5be57876933d490ccba63563ff0d4cc0eebf3098a9fa2a749474f9f4c5513fc36a7d4ff9ba02a732cfa5e9044ebbc11d2caff3b54ece1c6f356a56c7b2fbe7c8dfdad31ce18bc359e2fda76c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h166a9912fed6db25534ec78ddddce92f82f02f10b450032c842bd29db710d424b93236abdabdf716a8057b1d3191b6655bffb959343e1d82f7ed45866a53559a99b4b00bb348cdaca264ef121abcfb30f84c3d22c223bd3c2e06fb68ac43408411b57406f18fd846edbcb014e5fd3ea1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7656ad429b8b1d41e64432d5b9055949643d2f2f80cc23abe4b7d18c0bf0fed56a6cf8da8c0737adb832ab07c6808edb1f293ae8048e0de595b6d72e8b5cbfe957eaaf1ad22e6eaa35bca1e8d64809ac292bfbe6891c33995e7b33c26c6e3ac7b7603d6119586c712cf620a468ff9c842;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h997dd978bb87ae34100d3b0f1d3056557edfe95f58a52961061ed3496bec4d58463c676a4a9cbdf0f72bfad71e7f5fb09f30c0c2d984184de7b8a6acd5e80635c37df91c0d2c4100f6caf3f6489cebf96c0e9e656850ae373aa94ce8504b5a9407225b3d348b82705c9b3fd135eef3ab4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bfebd1a35ffa8fbaa033e553a433209fbbb691a1033060fb526467bcd2b9d7028fff644c84547850a53dcd22307c48818683dfe2287b451454184a2c9c45c237d735403c32e4e75c3112c1bd87c0b68c67ba30bcfda22e3507d07e0e287c2d57b724bd6f0403685f3753cbfc0f4d819b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40c2b051a4a3cf3b9d02e721748c1e5a94481d7cd24567eca892e009646625555d16989dfaf826afaa9cba366ce98fd590035a580ad9a19e1caa935e9d34068d4164da89b32a10ac715d81976faa70142a0781a83c0edce80e8d9d87234d0c9728ffdd7a814c4ca219b0bbbd9941cb1c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4876c7eeba7239390815392860f94f8f39d0daa8cab5aa220663a46196c91108388274ae70776da8f840be70c154af783d0d09fe6cbd9f10e983861c68ec4d19f5364aea9f112a4a7d24eabf8781b19a39f8c226ff9fe0c92e66e635191e2b6d7402040cc36ac5b60019e709045dba2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18ccc683e073c914a0f2fc2bcee3b113126b5802c48dfa228ddab2636231f50daafb6b58702e14f77ce9986c567a6cf87e3867f795393d27d24e15b3896b27be37171384e0112112f82cbd159f89d2e339ed52282208a8198395261a673f4119357575c1cd3b183ae9c245ed4f5eb5fde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48a8399ccae468ac698246a72f00bb48e5639c5277aa7ea7146cafcab5a51e9bc3c8792f7b5bed6c02a791e9220f198093239a03a1cb3c20cd8ac190e481fbe79dd3a4b39b1ca507bd25c1fc5c2f4ea8ca087ea4852c337a438d1af922b1641401d4095f7a2b629f60e6edecf8826bea2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9150df31fd3b5a7f1c45de06a33815b39d505237d785d839a368be4ccad4aa968f62d4b15a5231a03b2f44908fe61b9bb4a5c9c3e978550bcd5f2bbb3797c42ea11c88fcaab7cff68a558f999c5debca81ed7e02add213dd11482262440b1319de6f1516f19e3a6afbfd8daac4ed412f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33f892f197d7a705f46c02a5ca74f99ca4e563497cdae0676d245940aa84d095010f0524ecbc862cff92a685aec4aa08cb9fa60eb2b5dcc81c8369f6638dbc92da3602db1e084940d10ae35fc4e6cb306593e9894dea9555adc82753ae631f0b24ec1d008f575a4932ec3a742005317ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdb637d951d7ea7e023470cd8bdcf60bd60c4871d7b85704c0a91fc050ae9f023f2590a87100f7b78e5c51c1eb785a65afedd20dbed12178e712d6cc4332c78cbc4c142ed3f22f538b49b311aa209f89be44f794c45b9e13f4691ee7b8ec726cbf55a25f6601668f250af70b5b049fdfd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8abc4ec48d5ded2f9fa5950765d21a2b4b62a17c4f6513d7807abd72b5733cb181071aae17db0f89c82aaaa9a95321d8cef44b0f3a845e0939c67dfcb992ba01e842ee43f5d261cd355a3751dafd84601e4656c16164bd9c752790b68ba278829c60c1dca6381c3c81b710b05d201b17f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50238d541d8c419a7bda9f18bffa8cf5740f3a8f37fb90b2db9b1b504370cfce9b8a70acc7df4d3674810ccb446ffbe9a3e68743ffa0da263b3d42b67ffc36fb949af2dd7036dea357dad09865f55228fc98a62fa799f9aabbd7aff2fd5708325c621d413e810b7753a0834982579d298;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48297c4c038a689bf8eadb23de47d9ce3553d6cd8128cea7e4a041bc9810116594cc1a2054dc55f8095326f50a914e89b432e2664075faee7b75231bd185ab3766f4d179654e3af7b1182f0e789d3d071b45df2c2bb4a704ee294225446043c91b77dad9181a123ca35a79c069421e90c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5bad7202718c72734ccc346da78f5d304e8e91d2c47e5d57f0ea6026c1e0cb23715cec3a3f863209909a6c324e6519248c1138b7c2b8b4e998d970211130958815c6fe902dd754930d3dd7c79730d28750fc01c858a17f92577995c50d751cc0f0ed481b11909cde38e19836590f1d41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf01e62a4ed8ba915fd6fc54bc2a91ab98b498faa31008f19b089c0b5f62f9c004631c05c3a4b13de63fda688a9f6048c34dbc53ab30c6ed49c7af4294ba3f9a6fa51aebffbc307852ba774f812ce22a7e0dbe8aa085998f15fd2a4cf4943dbbcf5f0231fe5bec219c6a9b98402b616782;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9505a1572c906847fad36eafeaf5661ff005cfb8fc2af432c5d6b5d9222576797dd55acc9b8c9c03b24ed49cbb1ef3407e568fbee2e3110a997a5d2ba176d8a94a221a2c6ab344b95d4934c825bd0f172b883654c38fbf60706775ce7db399b4890cef037f320321fbfd24e627b7935f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58da1cce8fea0e8660d2490f369a629e7a4db621b13913673bede51c8afa201580e900491a780bc751d2aed5b267643940306e2bb46707161cb1136fccdd115dc14d99771e965926b8657cb56f51215d48da822fa69b578e29d26b8d37ebf14c917707eb66af65fd33a8e5fe6f47e3acf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d8825ded81b00f115e221b3e1c5f31ca0b55dba41592adf6bba6dbd5748ee22c7ae9cea98a3155f95f4df7df0e7dc88cfd63308856b8265c5c7d764d4aef88cdc7602967f33659ac0b211d682817ef60b3ffbcae37871a17a654935ce1a5527f5a9e55ceb2ac6cf2a67f40bb1f94f434;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2b030ff1958f3519d853dca7a7bf9168fa50d431c870f08746d974a8e8fa0368c79bee4bb8b7ab35c78814b87e4a754baee12788d1b19460a885bd9c179d4c13697612a4d56b0ba106e1d6d67ed357eaa1f829edb1daacd88c25fb817e239f9d9e1f38796991201dc501f54482444f11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a79feb0a6e7064f2534c7c71e8697cb2c80d407e6a215ab678a3ecb36d8ce7882906545e670cc68fea3178c02bde738c747f8752220b75eedcd5dbeb0e708756e5154cb2262cba014a94e1d4ca824054cf1aa7a51bee86106d975fd9319a78a14e772ab80ba2063f036f1d748df1a5be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37efc417632949ad653dd524986f9b322eb3781726d329ff7eed3273df331a15557720160dccf5207738d081081b32ece8c34db119ad5bebff8b229c66287f31f9893e4fbc63d71b15de374abce50313ac1bf7d98a21c98998d92a313a5677cd28cd3c8d9c913d8a379a620b219434f7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba089509559f8b463186130c2282e7c35eb7a6d0b99acf98bdee7a200495fc016e26c00e1c4799d41dd3e0034f6e90934e638fa4e71c348855e435327a0d5ee7336e7e0676939c9432a406a0117a5e4bf4b31b6597260f25a66263eca4740c3ee87c4775ec522ba442eeeb8d61032f056;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7fda2ff18c424617951cd93d8ddd5b54eadf51f1a19529ecb25c9053a1779fca1552dbddc7a503a60a4bac462b5c10df756a97c1e482ef256d743ec02fae21c343e735975d452e6c760f77532189f0f8da93b78f311f5be9b1df1918218cc8ea2cb21b6e7e21d57ca1548c7281d2be32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc005eb7f903b4e891fd16075a9d66a2a1f57c92e17e652203b21bdea16b731e11cfc82147089f6c3cb0a44feb7dffe9c32e90f4a4603d69498c41ee08a3308ae0ea67e13adb6aa745014446502b5e3d388418f2844ce8397f21252e968154770786d8499ee1bf8854beec63a4d1c76ffc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac066c99341b4f4ee5803abf58e53f8584141445b5e66f4334a619e75df2334339fd3f1c404e727621e88a29517fbaa381d916bf1d6c4aa6021701a2b0c6612eafa9952501f9438a6973976d61305dcf33935f4cf555db9f7671878c62718579f03015d785e5b4d6b267d5fbf34654620;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e25cdea34c6718762cf1bfc0bd13ac504a1ede37dae536f64435c58b69bf5692b2987fc8c7d453c90e77672157610762bf2e14f746d9b8d7d252c90756c6fb3834fe2cc4d35b3c2890c24b802c56489423d45b7ea0dd133956b65035b8bd8cf6329ac49d4c369893281b5662663b2ec8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h120f22ec293b8e05680aca0c1c5e85bc06634b72ca3530005ce1d4c27198a6de9a19024c991beb8788aad9321108399405cba6597db8235b9ae96d19dfe08d0ccc2c3caa64061ea9228f5ed6852afe2ed12c89c0312f7ac195f6f00b709281d46433b4792f4ddbb9642301a7537bd44e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cc7e7d0710a124d2c041115bcf516cbb7847fc1747e4b7744780990c85bab99c377b75e547d481eb2fa7db4d8f7d8d3db5bf7439c63e64789d88464785769b45e28819922623ef54487a58dff0cfd602ed9c0ff005279e8b9e0fc55ba982ed25f271893a01e39e7e10a7a6d410ec958;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb520f3d5425ee9ec39e4b52673e2c7b28278ade942db8e2adc67c58873f61bbde7b6cc7e5362e1c6f1244b98f8b51c1a5a3f8ce14890752d99b6d6dc869dc882f403f1be646262edd00521aed09d0a3f9b523f9e6d08e7aba6d9cc69ce6fd7a6c08fe0bf1097225fbe9bd991f6d287ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65cf8306adfcda83e86aa92f96163f6aa2b678c45328f589d49a7263bd067897c160cf593ad57c4ee85ed778d7d2f5816689a7940b40f1f7acab73557b379a2dd257798ef6b5c6d57657fca0c17a73e627c23a597a6ba9e3817c85523fc8cc4353f5df183d23f9c915d73b498b0b728ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa4e04e06d721bcf74f57cb163bc93092aa3336a4d23ba99994c348015a1766debc2ebd6911d554a4d05318762d474190a04c570999653d6ae2260de3e5e8cd416368309ad65ea36e8f13b5cc11ff86dfb204a487d617e640542df1e05fc601cfe60af15652f66328fa7574400d5950e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dc1aa94a546515c41a5bd29a45f94f945591e7fd24e61e8fba7ced2288730e3e4bcde7a8655c7a387499d4aa2cab9a05b65c616f2b2f9a8747f322cf0f3276cb8d767a8224d64621d48e5705d9e601f093375548a7305e8168a0cc6aa2dc015a0bab7e23107d6faa07b04c66cfea0e92;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h124997b360e267de5ff7a6cf8863543d186953070a11643daadd1f97367fcf2c0ba0291d9a0edd07bff0055bc46cc28a9a8fd6536dc2f5c0e3e87772155ce7dba7217a128fe3449ec6a509a531e6c45aa1cb5b008398a225a618b654d1cbcdc876418a60b94f4d957c0f644c5079b9246;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ce3bf6d4d8418f00c52fb7ac98167cb76b5b5297f097ae833e91d76e9a93209749718380817a2f8fcb5fef8d943a99864a487534c2cf7ee46cc619253da415012c79af12963a9f96ebf425a36c812156e46ddb0c978fb7ae6ed0421495bd6aa89148f9018f78b5fcf7a19697034131b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5df51e1604a02be6e8efd5eb2b40d48ed9b70a548e15c60bada948a2940a271da342a7ceb981e01ced4280de8e9dfb1236df7b8caf1c3f5b11e21ea824b62d78c0bba74fdc5bf5b55d4ee25cb5325f7560c84b528af59c0dba3f2ef35db54cff633fd0395e483dd26d4fe4c742228fa29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h328e7f61645b6e788045ec03120c934e4c9c9d4ed39931ce08d156149da81aeeaecffa54d22ed954b552983a8ba3daae37aded58bd3a7d86c5ddd3d807c213f822ed88229a0f90068b9faf31e71417d79158e1cddea3d85cb61c505d49666aa4d95c9a75c96fa0dbc67addb6c47e40d36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca648bf0372e4ed67ac1b236eb1d38ea434dec012acb598a7c1ab0a26854c811e1a4cb5e177811bc564900ce560b7e6e503b82c2fe5725eee72de2b9cb193c86990d66dea11e6c432e0b2e5f95dca93a9e51df53d9dc84933ab5e762038ad0114ca1a7e4374bedbd37d50022b69e25d97;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f4efb83f620593efc2f2dd305e56e8832bbf1b01a023115c1dd16285a182a836194c685af3c0fff6a624a90b421b7717e74ce370b5f8e33fc51c66717ae06d854d4d833b5cd7937e3888cfa076dfb9cd51dd0af3cff5ae595fd1b7c96f559cdecedc6bdf5cfb6a1fcecd1b595d4abf45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc859f8a58d76b22b238688fdae2cdc29c74c7ac3d344d4be585ee6af27525cd3c26205bdcecb50866650182c472101351ea00fe961802c65a1d0f5e2cd5b2be09c7ffa7f39967315fb26d0fddd3201377c25331917b26dacabf2f68bced08e6900fc064695732b7f7a8cc6f5f73fe7d43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h266fdbb0f100fe3578a77e20c33cb1bfffa9fbb88468d92c1b8a1e9b453ba40d6baea7af2791ee1e233b27b551b67fdd47ec7760f07c4ad514a0650b545a407745d980727cf663dd273ce19a6c9ae55385d6d5227029ea164dd17fd33289ac089d90dbe170f1dd8c2342da5ff0013f2d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90d9b2f162796e9167403fe3518c4ce9cc387c43c2cb64305eaa317494aeef20daed1b6370808b3cfcea77362d239801856842c0d3068b7d9610137d96b3c37cb6687e744b12a7d363cff1745ce5d0c2f5471cb1dc10c10507c523f46125a8b497777a97c34b3cd1dd2d1cba42a0afd72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee2fda487bfe5e94718fab4ddee3f13253c8a1169ac8c043cef9d548209b41c5a2f18e9d10b2289101f7e733cfcb937004c5148df2c760bc6467b930b063c3e4af84d8cb6f4561a90a2f3dbd885c09874e78d75d9007db836623b1a2ce28fc728c8047c3dcc7b4232c065c42f07b2a02f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8229e2046c9e6d66c6ccea6fcba870f68443d806d3ecbb721c0522d8f7f0b55fe3d507a7b0e0a981746a9d06cfa35e94b52dd8e14e7c0afef5680a289e5f0da5545faaf15424ef728313ca8b6a771b74d5bddab595fa847e5aa1e1d00b91390c42cbbd84e366ab8ce28bc660447f1389e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb553129a68657ae3f8efa6f863ef6534b6ecdf4ae1fee40982e0d71ea8d0f5925491b1664aef66553d492edb7ed5ac1dae685b4ffb39c7000ed40224edc82e70c8f5b045ca61ae9987e23c5cbef20b313100792c266638ec28833ffae973370fc9deeae792732ede37d7ce6661a0554b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc75e093cd1649fafa2b70f3d0ce0a68a6608f20706032c8c83ee74ebb62d21d2834a1a56a331b59dca7bd4806831595a31d2750c708d437664d0c7d9e35e09a751ac39808f5b86542e41c9513433983d96af9e57441b995f4586aa40a480774f5047f6ac4670811e4d61992014fea41ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa00a894f73a0d98a7510d08f607d83035160958bb49f2d5442cfc30e4548adccd9d1d05cf037031137dfc5510fe700ce736c7c833d01b537fd62c7625b20173ec944ed1d38c43807bbae72ad02dcc8c570f5a9f76b952e57c52b866e19bb8d583a519c6955a4e31d5a5bd32544dbbfd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1d15908bef7d0ffe36c517d83ee01468f8a56ebfc093f76e15540b1a921166bc131365f13944107bff0c1397faa5dad853eb0eecbc5d0d7a90f1b62ce50071352b8f90f80ebab45534c69f29fe5d4fba5164c862e387c18a15a33b27a6c3f7548ba76912c17b594cbc30f38c2eadf754;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee2cba88dc9bf98489e5519c2caae69dafe18626dcd927f14efc16db90133c9ff5bd387ce9be05ca5bdff32b17e050145299b205b9996eddb3e49c4b3b6dddc8bf5cde16c5e7b24da23ddd408988c03001fc80c787a631276d6d2e6f1a465344fed05a7f8a206bb5ef174c7b2d439e95a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf19732c7f5980ab4170303f86d59bfaa5c1644449cdad06e20ac2bafe46717e804b2f76b6c8295333eb1badaa313cce57e1d7640b3a1c13b87597d3ee1c6616d9a523454604639141df2e8966b5f79d90029be7ed0203fe181cd7fa4aeb69d8d588abf59e938bb11c3a4d24560f47ce2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h519507ccc2aaa9967dba1943466f7cc6099056f13c2ab9853fe10a1da4f3e5b84ae188c9972cf8cfaef965c9c52326849c1070135db95ff33dd540c146423937612ae17a6644b09bfd113f55218b06b6f8c4e49bcd59fac3fc7c0b7e407a7828b487aeb0f87d15769ae20621870e81320;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he619feb9ca7988512d7a408e789ebbd896164041914db3ef286bb7eedecfb89474f38996d1ed7d641d71122dadc72a1f38ecfb36ac742ad5bc15698c087ed820e4caa68932d0dc835663990081f9356dc4af9f7fc9906760bb735573a556a38cc7836bcf648211a3a4139cd0a40385f3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37ee6ef334cb22ee188c17e8e73bf4997e8c670dbc80513d91793a4b6c3f5dfaf638e61100c6cf7f600f3dd33c61df4a9c9bad126b6646c6723fc677096f7061c14d59be51bb6b7c02bc7eb52aa9c890796bc29606b2062e53fda2f22d9ef8dd6f84a27eab820ccab9c55511c8223154c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0c6a4294775b23974f57f97a6e84ec1bcc65ed028e54249dd77251fa7d3e3d71465212eb53e64ab78c745061cb9fe17ec6ab16e62c0bfc175213162fa5dbaea576ed2d9846ae4e135683a027f151857a2e207c272002a7e96e33b807bf8076f7fa0a21010ca087951bbb5c5b1faa5cc0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e06577ffb4e8b5b10d3c535f45909fef4aa0188702eda23aacb0b945bca3489b7e151156e3ec0c62327a5862711a49399337c687aefc66e9b9b045f6732656457b432776aa7089950c63ece4ce155be5217314b799425e0c92a5d4c0314138ed68afab9ab85d5cd495d4fb7de5c0abf0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467b3b794536773218b56ebadb998cd098c8bcaa16ccd0aaf230aa7c6241a1986f75a82eefc6d45538587cff1c118696e08825b5d17690168a2d02b1842e33ba0f6808eb2936c7833c9a7da09e10417baafb485ffcfa99a7dda29ff89a5a845ca882dba339d9930c3cf974a311184b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cbdfd6f6688db79e46650022bb79fa3c5e6bdeafa75ed7066a59788819980b65d94c375ae3132816c2dabb2a9f3d5df1f7ef8562fff14066085b22204e020e279091245f639b90762e88659f2428814e37089c0e99a9b57b90d4e411a12915745c275422f752474d92bf71e3c95ff4e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h296d1303270b7545cbe1470da50010490780437e0bb3b292a8c5651ccaba27b5c942f96310d078dba7d764551a5faac3740ab7fd1cd1b2ff8c2ba1dd8f7bed82841dc8d35b0bad39fe70af2f1a26c93e605c4e1558c79a53dfb6d3ff57be7226664763bc9468378817e7ec46165265a15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c430c499812aaa995fe6b0b8380af2efa41a300986333442442d29f44be1fa93367ba7cfc14dbc93b8a36251fb172c05db5ae80d3a6c778b0550318f56882d843c0791e8f1e40a215a87d503d64186c58382ef1e23991638a65382924b909e1f5b8e612191c99528bdb95f8e77863cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81f6e722d48ee27a34c66584839bc182dcc8ea667905e6f0e7f840250cf3848cb7eb9d3ae741e0f19bc45c695c39f4ed6d0711d2816f02ad6f2dc7b9f511f5f480b0241a86ed55fb6cc4afdcf94716ae3ea3e2525d94ef8300e26b0da295ba3bb1db376bb4f3aaae87ff465a6d7191b12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69b7bb0e473a44d120562ccec44ee7a8328ca04afeed77025e9a9ce9d0788b874e43c63064c85199519e580d977bb6a65a0d187d06e4274897aa3c30d5b3a7ca5fe34879553c270fdcba4c32d34a4a4e4c42fa98709a5fa5044db604eb446562ab4f2acdf18c9fbca61fde2d3eadba88e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebaed86be5e7143ccfd5e01932a9e9c1f687b32738d71418bf909dfdb5b8a6d86644069808f0f1278b5417019abb23b5adf8c412d153fc2ce4b43b5d56fc390c475ee7dfd091c0c8db9008052e709734ab17878d3f780b9588f2ade06ccc1e450fc2692469341393071dac4e6d1ce8b1a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd0ea86dfea04a0dbe5682e53b5d5e85cf7a6fa5f91f3abdabaca80d6a2c8a706acfc16db613add65c29f9c7af80bd1511bd90cd1b7d515247ed77a378e6db6b13e333a0f894de5108528a02343338b9c0d9ee611414b6e8f7601aa0c1dbae08b313f2e33b50e083507d58c577784aad4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c062951e3efc8f3244b8369346c01a4e1d29251e758a7c22f5fc261557317eee2386b84a40dacc6b4d49b34e29da77e09631dbf4f836c410756719f6ed6dc46a6129f6797ea5fa1ce428b68d6c02285662ffc4d3bb436cf3537b0e13ef4b683912822a27cb011ceb951e249a08190a4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a321d2287ca93811db7ec0c07dd2d581b8e2379148f23360c1f9e15b7b88d71ecbd3e116f029641d0ddf89821dbcd8dadd9f44861fcb9e6234acbdb0067d8097db612b2078075a99d19926e81dd8cf02205bb99a1ffc5c1e4027834050ee716d988d73ec1affaa3c1540aedc6118477d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b33e2b1fd57e80a0071755bfc8ecf87009b1cdf648189d7ca2ca9e54d3ff1ecf5e951703d8136040792a00da1b3f8a99144dd7176e2957289cd2ee08ca9887612b9047746999b22bbacd7c462a5a41c17ac7920174ae812ebee46970a1a542e6a42e399c5303a52e2e93df6959c093b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ce98cfa42b71137a5f17ef4f7dce91de3e6b4b91d0f4db7e2bf7cdb3095ce6cd230b764785d86dbc6304c7c91a688e85ce50e506d0c40778cb2604c12c31cceb2713046618a1555bc9db9f7b6768dafb9287d80725c35fb227987174515099ef528c83c9da9f1fdc0efe560a000fb3dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7810cb195d844fad872ebc22e808d7158e3f64c983c6f5b632e9213f9ed0621ebaf1b93ddbbefbb2184e32d9a34406395da3e55878658a553ea8eab844c0d75307aa565edcc99a913feff2af3b5126952155a1448bdce42c08158b0c9a539fba7229a44f30db964b6ee42b0ff996f8845;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12ba693665fd695ec923034af6a5cc40e603fa5e7ad43ced2ecc50261e379dd263a429d9f949a6e6cee4520f3e236678658d275aaacade01490c6d39be3986053ec6aaa78a65e4b221c374c6c06a1eda0c344daf119877a5fd391163dcf2f41818a3283581b3e42c4b7a213df305e4752;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1e33475ad69157d6c7cf09247c7a9f9acaf08fe32a626f74034c8a6425b15bc598e0c1b37e58a720be65f6e4447ebdff8eac58d53287a4dbd6ca24d53752bb09f35078c7eec2886a560fa0421c20cdb530011f92b29cd4b1ea9b6cacaa2ec567ac751f8b56a1e9937e69f8889c4b1a32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2de97e58251b7509636ce98fd56335d43dffe5c3766e622b892fbef1da1cfef75a88fdf71c6e9c4989b7d8dd5079ed9a45fd78468d4a36d9701662740cc9086c9b60dbdb039274b670e053efe1a33919f432431815ce677d0719a922afb8a8d03959543397d060da3b31fc1e536c6eaba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcad5222ddee8e99d84ab01da763819f73642994f1943c0749937f6f6fbb683750b5a3e3e4723c3b55b614cd98591ba02c2efb40045f9d794ce40d52661459c109a16f8adfee4b010e9d01033c8ec8733784bac75c1cb0369133a16f2475dcca9d0beffc7baf707a0647299b9b02382670;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3cc614934e0ab9c5a8e17ca33d2e201ea76cdb16ec93371327a344a175d58f8c46fcfeb424bc9ec27078f5ccbe06ea0dfa961714b28828ba8745f4e847bfe8999dc5e0f0ca27b2dc09c3181f08fb6b665d00d07fa2c0d82f8a0b20a37c03b689234316703a3c16b0ef2773cdbba3a74c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfab78902c9b0d6efc98971204254589d18d3c670ece7aadaa57cef0b33f6be26e19d55c67c4f1703dfec02680d29e6d1b046b3c65061e543e69463b6602feeea1d823df74a8bf51b2a5d81d55929a5a299d9a3657d9e1a5ecad1c8267c995384d7e8589712a363ea3ce66af11548d837d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7120510bd0c7d78963f718b52ef232ab9a883885c885bbc1a6f7ba8132daf17f4f72de922293c45fb8cd3dbfff9214a3ed7eda753e2d9790137fbc5516dbdfc0aee194f2ce61cfd4f0c3d088a88bdae741d70fce3c7e50e32e09131ba8f06c98b004b179fc45f8cfa19d554e7a3738ae6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e3c0331ef08f057bd5831038542867f89832c536eb27b662e9eca711f0545c5cde5c56690317ecf091c60bbcf5b802e0e3b8da42f55ac0388fa9b39b628e3dce328c90dd0da1161d7ce309a95cde38c6fd3a6bb667b23abab9800d0284289407259bd0288cd21d7c88eee455bad6acc9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70cf89d8022b18ae701f2a8f51f23fe93540fb117e53ad1c4d54fa0cabb932fce053ba6965d987a8c1444abbaf3407bc7c71096fe61c05ed161db2ef0d75a5f31a4fa573009b337495c3c826cdeb6a44a66b896fe96e08a60f8f37193ac103f01ed3a3f1fc9ac7d3afb24a3248bf86f20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h684e32f993647bd98dc50f2f710246c2e9e4110719bf00a5c2e5a77da7674a59991c6f8697a8faacd3d46550462cb9f90059173c89b7fb095d149b9f2973841c6570215a042e6b969621b5f679d2841413cd1bb1df147ff912350ce3dd9f454809a4f055c648a1cb3629f6bcabe6c8347;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45130de5742b6dab6feac3cbd8cdb481953a96371aa00abc04b696bddd3bbffdc78eceeecd9938c0bfe55075640cae21b35bae4c8c27362a853bb20319ee595150e6913415f0d4872b4103d0310a5794402281cb91a6e9ed2b91cc7a30ef62d8bd5e608d9efdbd7199002da3280c0d84d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heef5c28b39808d49f7f6ec74b92a0c7c1e4f6bf7744da4cae4c9ad702255549965b3c84ebf9beec60bf47406fa6c67f6eff3ef59fed8774947eb2a3bc8941d5d388e778fbd067232dd76aa3b8c82c048e0ce7b41530e858ec0b11994d92331a5a52d69b28765a9c5fa56b4549aa0c5dae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70bf350408039bef81d7b72faacd9aa87e051b4fb78683df3b452975ffc543b5efbbe6c31209ba2c4fa7d69dea4796e5a564476fb709c6d6f09b01ba3b9e07793de4a0810cd0f6517fa0d56f66dffca94603c918c6e12e347d66b050f4f0aea69e0a777c5522bde351d5382f5652cef2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde0a092fc6fd5dbf453fed078080c8bad3a04779c43601ed671670d345d23d052e979d49b61068a3c588086b1dece04fbc6a2eb6161959767fd26589f462d0b7cdddf1dece091c323a7d3defcbad95d30f1a8139410e34cc311060c856dacbac611ccc6eaf253cc0a697562a4ebc6496e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d2a931a3034a4e635e14857515df03071b1e63a1c00b2d407832042723f7ffdd1cb61105e1ebfb094c53d74e8e29896d8dc150646db8aec76cc1d2a96b7c54a7ce6892ed497511f2049d01b94e9847dcd45e4282e8529f789e8190d978e8b4a40fe1f2c026538ed610568feab5def61f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2205f721dda78a2ce96ad66036be6f267f14aeaba07cbd2d745962b1f2f49d22848279d97621c8fcb5907e2d0854649dc1f76f134ffa0c7cea5030aebe46c33dc5aebf7eb9b89934b8ad17fde4680a3e830eed2f24c45613927a201f1357712ead29b38d159b0e5af72bdd40fe97ec058;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5e9c506ad53c994f1a94c181feef27b8ed89a692c4b60c69c4b6c53a4ee0a3a04c45b28abdd4c9f111d00918481b8eccbdb28706d38854945e3e78431944c8626b4c0a9710117d66574c18954b6d01793260470c0ea90ded894bfbdbbac03008fe919f80d30620ad59095adb0bbe5a1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h670425855dbe4b21568101434bfff7c439d6b39edab1898d661435db0ebd1e79613dbf95ed84dfb3116e45449ec1ba092a5c35d7015f4fa714583d1fd0579557c292d2a5612f85db537773dfea738b744e13a854798222ff86c11d1bd2ab0327ef59b719508ff02ab15d0a6e62de8c5d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h644c14f7f07e793c37f2b447e1a5d2daab3d38e6d687edae9f9e31323ca4dca20f527325d2dcef9e27c00bd53105edc6cd905b0df20c816f045c2bef89f17536bf4811a6abf8f7522958476aa2b1d2e81c72dcddabb0f01454a2782805bee92dc4920bb7589c9983a1baec38d52fbb1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7330b75697638e5121b5db14acbbfb77415e0d533b15635aeec83c2f14fccfa6ae236ff82e48ee580cd5c4f6fd02507cb9819bf363fc5a54b3cea7e5249cf006f6ce11b06ab589bd312227153a264a683d8e660b2557938dd499ad0d4a647d98bebb891fa21af5e43268747be4ecbd75e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb088afbfb5076387a29ef3b7cbf5ce060d0efef1bbd4365d75ddc3cdccccc5ca56a730395d1f73ba307c64f0a7b13d536c1d19327b224b844a2f7364c6c475f42f357dc61ec5d6df5f9fd2043ca3c854e0ebb1cf82e56626378af9482a5e3afe0b7c564e6f3d07ae4bd8cbcdf0b920d30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26d0b39cea11d63f251cae7e8e428bda63f7496380285799823e592b4ea1574cb59aed6bfee362a36b3b67356c9e4a8f0fc9420c3fd1b76b2001c38230dcf00b9804e19d91669397987cce8155b77ec0fe93de51eeec9245054ccb87691bc992f5c9991a8a597d4c1caf00f7167d5cf22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc88fa97ec58f3f7d0c5b4bd93f006a18297b13ee453bf96596bcddd6cf12f9686d21db083e2f9795858b918d5f6a897722e6ccf1491fff2d2376261c72ee91f5da2e8924466e24255a325093b0c967759d53fd8c5de52049f9105df8986489f3bed1ac918b11112e64ea5092becf24ff3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb83eefb604ec30ad0ed3934c67a7ec07f75e50c1d3292c3c07b7b997a14f8eac62dbfb66d9a535832ef10109608826fe3ed284ce3df2e1b76418cf015a08106b1c9d139c6456804c34371a946c6fa7681d9bc74bbb7753c9ff530cca39a52de8a0a9d145176f74ee38f2ed6d0effb193a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c3b4bbb4db4ebcfb238ff3cbc480e1accf8b8f119cf1d2537678b344c71f1d7b7be870ca8e877b549c1b84ef53bfbbc1b12f41021e74a9028e8567b42835a7b2489ebb9c9697040f7382244a6a025bdd32cb604272e85b359d5185e3caf175c787150d806d6440a5dbd748b4399f36c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9802fd6eb3d9be3c69c1d7948abd5e6b243a50dde5443b79b98141d48a7a284cd1c740ba37b28de3c5f5d5c621e6108b6a7aec717df1bc155da25a3c36c920af97c73c3102e735cd2c293b768bcea82f338895c3c167831112aab10c313d84ed5c94bfb5dfd6b712d61ed48072682823;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20b63980e080cac06008d654bd8471b042ea7972c6c789a98c5d36dfd749d8171d37075875415c93f4863c1ee07fed869d976ef52ea0058a8cb693435d0e9a1837d2d3256c9a2ade393474bd40110b7a7e1c18c9c1483dff6cf41ac35c78d70354b6fbf5cf89e527d7c990a3c06c9da31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57669e6ccbd3fb07fbc69096ce713d3b0dd89a39995cea8b8ba2fb377aa7cb9931402ad26406df89d9162ab77dd9db1b42706bd9a99b4c3bd85b1a9b7edd8a7f660e27662d206a53bd13adf9367b412186c233b8d17410042700d0069aa338070dbd6f7c7e256675a32810962e4ab856b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h746a7974cf6a3c71bb1df46182ddeecb5a8720273e85a76a9590a0a9beb60a6377b585845a9b267819958213e097f337e9d02125a42ca295d8a0493a7c86e5edd6689f2f57c6ea1279b8f75d66fb4b65752a53e78e3a7e96ca1832539590f3e4678125e040b05df6f427fa0c8073281c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3753d8c274ab4f1162d9197a3053747719d8b847cc599f21aaf94b1104f8067646852793c1afab865ea58b6acb2bef0c8466c764a5833c284d2071d61618d1fd0bf48e35fabe29bcf78cb9667b42a77790dea4aa6fd2c48db278be5f2bca9a2cdd49f845f5beb1e03a08324fb8b5077da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b4e07c8ae9a1785eb23a3bae5fa91ef66ab71a0824f6eb38427abff4b21fb01f63e9c7f70e80eb9ba47ce7f7a1dc6911465a6cef0d6171f2e88edd9da5a6ac88ba0a66505c0cf2ffc0fc383b9f0efe51596b5574220d4b99bccdef49135505f91e8d9c49095b796239b0f934993eb0d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b28d5de5bbfe7a3443c312b026829e9a52d5be872a764a344284189ce779c06530ac6a62f8111ff42eca08bd3a9e861febbee188551a57adebd42d61baeb1d2f1b7dc9ace17e8c3ccfdfcbb3df7b1164e502de5cd9715eba9a5c05af05b8887a87a288a63c39ebf95d61c500a850d2ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h524c4a8d46806132b7299252df609d69b8fac7e0e6df8cb8284fe6edd0f392367536f1311db27e78e1bd679e71789b885a3bc8254fbab2ccee6d6d52f1a004e2924e2cf4e612e07b378e01eb865f04bc0b51203c845a7dd544a6d16a25f18cf6fcb1bcd9a5dd55b25b9d75c1dab44d3eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef56c60376ad1277a920c666d56fcf79503fd9c1be5eb8f2c4fe966043d68ead86ebfd077d4adc121e4e196eb6a6637bdfea8e6ef374d90151c55daee8b6c797735d5ab101b872fc7277aa703e95420c8260337a141cfcdd105ed85208f56f5d794eeda9b2c0f3ae1d129c9b41ff2230f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e54076a323fbaa9d12af31cddbdce2bdf3f66ea9f53c5e6613835d58de279254eba053d2f2ab494293a1c1cfc89d89d2d63c1bd23092e20f8eb877303b92079cd184aafb569fdcf53f80cc6715689414a42695414eb8a7d5e7dd1145ff45c9180b2bf4c2dacd24b88b6b31e5b3d41d9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa4c2708f40397ad9621943472725e200732066f926c727d51c87be6230f170b5d51a526e459d95c0df824e5512019dd29cc43797701a6b50573075a4ce0bd9b27cd226e419e58c82defc933477387eb0d571980d5aed3491813987979a385da90ac944df1d677af3e6a56e9ec0b036e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc86a491f75be074cf82a82e9af776c362b5f0488f900486d51dffed237517fc2538a273833b98532122844f5e13f0bcfad639db2ae551939fcc67bb03d5b3ab00833d644d56c8f5b27ede82f1e1aa79908035b4f9150d19ef977ade86b8645175414ff661b12b2912613d31c2d61e8640;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf741a18031cafb1f8ffe03e23667d9e3fc131f3d84406c19e0061acd4bfd08b531f2fa61d827b5404176b4adc01390b97e2cffa195d5032ec6eff4a61d218b6f7205353720efe304e5b6ead9ee712fe741b097c2d458e19029539028ae18ec2d3eeb716e438ffa4650a68033af422615d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6748fec9d286f4008940b10414446661e2022ec6a88c435a8076deada385317b7e775c54707d0b950f762165cb7ed7507f7b962630f5a84709a98314194ada508cd5252542e40adc41e4eef78021645fe3f8ce5a9ea45cc7a25ff3de024a21aafb29c133e5ee7e1676a4f194e067772e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf47e323076e67e5ad38cb1ec757d6dfa4c26ea6a8003a8e9b65428e33cd0eea76377bbeddb14b02e155b694e1f50a64ca8626d5de1dd689a8afdbeb0f197965d83b53c2cd5507fbcfe78a2d459b0afa46b2550f7f51a3569ea659b732277e7a8644b563f602d0e1c2129769225ed918fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4befe5a38bd9a2ae64fc153081fe9040d685a980184ad22cfc9fb64ddc8703eef1667b2f65589e79f9ef31fa716ff5ca089ce6925d75d3d53da3eb1d8a505b7ffec082b2aacd26f6cdc8a1f95fe2f14797d4e05a618801dcfddb17f309698bf25e33b153792b9f80d43991833f7b5d07c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91570afc19ac594026f1a2bf72fb4387933a62d516cac102d9a25f730a33f1d8dc0590ca619a38bb09b28041abb0fee5c0c2bbf2bc3afde524e67356b98ca4bff656059ef800c7dda19d7b13eb5c9e223f2ee4671c31d938b421bbd2ab62681d06b8365a34cdc5c8652fd59fa35e48e5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8afc1ad97017aef0792187cbe57cc5031fe5739323f0bd5be79fea6feddec11c6c644a2895b592a495a7bccb19b08fefb288ad6873efecd8e5445f864e901002b375384029a4a75d1415bb096e9d1aafca69fcb452e25f0f98592c5a519ed2ae7a840786b59633ac1625b55fae4e477e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcadb33713fe1fa47d4bd2a21b61a03cbb4d708111475551158b3bb70d5ea24f5de07f0a70bbfda1e5700895354f23bcce5ec9c21ff5c573e958a485bbc6b263c1c75f55725cc39c478bfff3796385c695f9b02795d7a06f51ed41b85e54e43ae3c1b1d5692788e3e2183507fd143febcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42622ba5802f713679c5e0b32c616df52499da40aecb735c00cac1ab86c334ef3e2e4cf0cca007064957c6948416c0117f9e8edc51bc42d68dd035d477da977c58a9a94c201d0b04aa973a39c1ed71ed5a465b7c25f06f286dae5682a974be75869a1ff5d56e156151b7a2c746d65918e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93db1f7ab7d71a9b072eefa0c3ccdffe85d0baed15b2367113ba03d2efcbdb4892ccba6993b5b3d9c2d087741690ffec8ea9c4229acbbac5c59f27ac6b999231c4681c2b6e8622d35fd39bbd31fc1291c3d49c852e6fd9e0aab12788330270b363a0abf13205f9ae081b6860a61d0a0b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3449b2cbdf57b06decb35c2535758dbf869fd58b763ce63e78b1fdfd60ff6425369918d9d303fdc53ba26e74f0c40f3bd48bef511d980b74e7005885f8376cc7a1c3174fb62ed8620a81e5af4b1a3785795b3d78f499e71578b242ac4f8cd7697c2363e6fc2cce5148030c33d08e45b2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd1c64b7aec4bec33a6cdbe14d0257d47db7dbf8d1bdcf6b2d47dae97ad5f0e1553fd805a5e9f04b4e2061ad72519ce9e26f69b5d0924e8ba99bae2c3c73477e0108e69f3699c4cbc05e40b5b86d6c1bd5165240e23ace53529475d1d634841f354b1e9551be352eae191260e452d2fac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9dda82ca911e665b8529557f01066e82a5f1e0ab2554d93fc1b2b828597c898a3e3ddda1b4362170e7fe941423583c808691f742360878e748ef04c9826401b100fc9bc0681914274dd07e190f76bb58b2e737e4489f944266942a738c08910c06e6ee5bccdf87132dc19b4e026da765;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70ba4d1649b635b4efdca2870d4a0fccb9523be9f206d4864cf513479badf8d6cf609174ba44d5e4f723458facdc7f73f26ac025252a8cab9973e88b4e5f9bd4ea0f8d06453297ca6d1bfa1b0609454f8b55c625f99199fabfea922778ab1fe8557353baeca0c740fb3f1bbf0bcaf34b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdfad2085a029cfb81b05725e015f8e2b9e9c0317e451462d1e866e730ba34308954aa3d1adcbe06f80db2dd75569b2bde98b209203f28817628e18259825594455d32a7022bd6ef5cba618174807d7dca1a0a940e685787909d31235eccb3be32b72c02ebdd53b95cbbb553baa8beb7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc32731fbab2f65738e6cca9d06add49ed8c08fa3528b363ea841fcdcc2db9f23ad3177e16485c45910fc9f32bd3928966dba9b648c94a9501d570db24a11d71a930721e415facc03c2af17702ad2085c1d5f684b171c907814ce073fa9a4d16c6d726593f32d49f13d96094aee213bb85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b89322e4c90a64b918cd9619a50f6dd8b1a24c54982fb079de4bf089e8792cc7da7d1bb6bfe43e632278e72e20eca06b6b237be9bcaedc4f001b7172fc854c81189d33e5c8a1e0bb96fe4b6d6d79b82ae839eb601ad758147bbc49ee22a9bbc9919d5ff6f5b8f9b6f98b9f78c126fda7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4884637ac2f2aae3314c408dc7a2475820821378d487d63c07149b75868ed5305898c7333d5ca4eca75736de55e2f6a4209e9559d3bece920f5197807fef1c5af5babeb17c55558fed064756683f6836c79c3d74cc66de3ec54f25cb321ac39ca4a775925bd7602c1eb09dcf4eac5056;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdaa0bc9cdc1040172fe9d7810be66d4bec5cbbee567c1a80f8678a7844ef8925751a370b7edcf91d19db8c79a3e51b2dd6fc6ea3e7541632c485e98aa465ed8cbddb3529933583314fa55f78bcf2d70963ae5509b8d821a080ebe3ccd2aa7cd3150a83b13f4d8822099c751dab7e155a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26c35fae1e4d4c28c0f2a7abc9f9f750290f2cdd8b1259047ecd4ceadc73012a6ddee16daf03f69d60cd7a1e2e082d0ef0a78bb16a264ab99af307f2a61015984a24128e4d3e166496721acf52203d207e2d77adf0928a69d1cbbfffec089e1259846e1680f55e88c1a146e20e22ac07b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92e2f98a417ca7c5f498d240bcf0c12e8749b182dcbd7450acf0113f27e21c471d0d8bd07f7fb66d4bbaea411393ec8a6d1cc9d10ed975a6c03656d2cbb6a39cb0963576503088bf863ed5c7dd8737057efe2032796328d0e514d31ffa606a480f8cf507c185f01fb7cf7cd730c8aa575;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec1d4041044da145bbfcaa4a90b9dcbdd26ea0c273ea549ff1a16d90a712e341245e7546ffe970f6a6af21195d88ea9fb4e151d80e79ea44eb1a0747f804b07f36a4b1b38b8a318842113cbdd648dc03773c2f3fd208c36d6b658cb5f97a9c7e8bec541e408521046b631322ef96a3705;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c8f74fce2355888fe92a84e33900797fb0f3305bab23f26a52118226f4ba9ccd4f67592dba8ef641ed9d0b8990c7660a864c711c15364709129dce338a6c892a322265fc34e8847a4e183f19a582e3c963c4dca42c839e07b37a07bff70dbae7c5e5daf4831e4c2a9bf90e216d2caee3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h254c55594d6233b00a3a423745543a826ae3e812b771e1a16c70ef4e1d306a29fb69522b38262a76eaf8bd9f894a33413574a089109e3d40cb308a3d8e33223284a8f64981ccb76f7fc85a7f78aafc2bfd8b94a3faf05f6de50ed93b7628597648d1cfa6b0cf50b70239b831ded366e1a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75775ee0bdbcb774a2ef2ccf732242ebc5febefe86d2c4bd6c31dd32967167b9e8a4fde019ed6f50ac9ce215713d9acfffcd6bb76ea40e0d3311a8d716ade53db322ebe26ecc1f97f37158ad54e0ab4ce34391f2c3e4afa620870fb0b6784d8b1f54f1acc5bb23cc1c7624e414e785088;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ccfb4b39758591f4b6f082ea9ca26acd76a073849d6c274cee4506d1cdd24767742200f758a30ce759196ec628a14f337cab71b0f26ebc296417b3a5b1fb765fbd47ca2251db143fc72fe835b1ba5a5bf2c89d941f585c16a0d8da796de41782f0f4d3a062d8bbad906c801e51a98bf0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd13d19e937e4cb52f6f168c5e83cc8f5d0477b710269cac714a58de78ad39db8a779e681f0a5612f1dcb536085c305a2f5d27a3d8d31281d4cb999b98a5e3aff1e064bb832f6c27aeaab91969f5ca0211017324b083474a6f3d4e5d15da96b986f26ea87790c10a47c06acc8a19d8ff3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29516b63ff4a5c9249f885bc7a6823a1dfb554821b49a620e1f5b8f40e236a4a9ef98c76abfcbb5a5a12b8ac00010c1a30f8cf305828be4ffedb519ef13c851f2d77dc20f27d0cd77a74040e0b23199e3e84bf3cd9cf408c6e6c1576768e83ea3dc096f95f4013fa5c7f0ff05eae26d4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ee65703d40acd9978f99d6177f3ab093d74a82cb76f202dd8eecd504341cb04626f1be85d41d2afe1d941a1f863b59d97c5144db80e7fe92b622019699b8aac08c4e99b5e23607cc2f6f7f03ccf9e4a3a275b3472c7e1e37a8a18a20394de6b62669b9f3bc9720c3e64b4d8626d7679d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24d84fd5611bba02a75c3ff9b7004b491fe01df3a46e07b3e96cbbb794fd94272c8e5cf314374bcfc060145b9cdd674d8a50801d14aec7d9dbc501c348bf1c72f4072df079da64e47f5e433dba6a20a7d910dc96494cc22302443c0d6bb31d354d29c1947124194382f97bccfacb9b1ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84a4825661f3a0d82cbbcc955e4c6eef4ab0d84b905c1f94a587d0d5fdd22309127ef0c448cccde8624b9c4d0a37d1e93067c3260fe6d4d37127dfd2ae7497ef538b81ee53be93a409f00117f6c975f8d53d05e9f12f669eedb9c282fab6c74e1918159acc41405c4668091357f2ec8ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91ae63f7ab8f53d7c4972ab21ddad24d0e909592c5224ca240c03612d70553b649fcd61936eaa13d23413ea86490abc8907b08231d68465b8b2cb98c334f047eccbf2661bd07dc7a0947b93289d4705963380a68d06066edf626ba7bd763133dc9ff4b25ef2e1c67c231f6c9a06518b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56679ce4db2fc0d36de68bd83c03937f13f94b24349d5173fdce655381869810befd4231e3f1d3176ef46f1b3cf8f5d16a78b90191de8aa6bd93e84ab806b826b5595a0438f48b075d327658611a7bc0c7476c4d8543369b6086f1b4c4b39120834d829b195baab96a62913da7069672b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb67d9a05b4c51be633eb15b13430557268e93e98eebb6a9154a7e0523a8cb2662b00ab3fc6221cf38821a1408eff9e05126b4ac215841ae0e9b102fb40ca569e1e03cdd6baf5f0c1d07a07a9c6379dc3265a6d21ec77ea37b23926d9e8a28d354e6cef36633011caaddc379bf7221082;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d60d8513d7a56e5b33dc14139babadd5eb276a2275e02498e24916c1ac92954d0684e6af33cd5514d870f9d1b00b7bd7eb9806fcab96010f3436d1c277db87a58de873fda1e90bf2323f95fddf1b29b256219d7eecf01691e876db4989a07db057b7b8d5fe9a01c05ec5d3cf374893d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h398bd6c322fa8537a753d5215bac93f483355f4b2e1d100b778bce0bb2b05ac774489c02d5ab002f39ca28e5051bef33f52e5a8745d85373847e4e2bec83180ef28a42708bb7e6d0ff8320044f7ecadf476f53271a20c43c7146dd280f0155ce474afeb99860da8d9ae1b3d4d2309e339;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55d5df5014c2137f4efb63d42b7f15d7414beacbe66ddccc2aaa88ab235c18191d3f9ff03b36aa5d465081f4e7fa441be8366dc44162aac23635429bc93dfec63bc11e175cf68df684d263924a3baf2268e7e3a5d20c61685c4f1efce4b2a17cffe7cb09e9d7ec60aef857bdc7a3332ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce4dfda0aeccbe1243b03447e75536dbbe6fc8500e9ca06543284fad3c416fce8acb98bbad7415a67f2e9f3e600e43bcbd55f26bb269b6887e67917e25d08dc8058adbdd2fa7c72ec4ef9a6c4f665ee51db2155af1f23033e90d8e483aa1b9f474e12f62407f4f90ab5f4ef53c08aa9b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8edee247ebe617461f60ff1d830a88ce50a00e96cd24a0ddf2361ba13b6c9e81a107f99b7e4640eb6e004e87cc9418005652c889d4d82ea0506b4974459277343440051388a39e98277e9fa64129a7471e3009be76f86a84f0a4a36dad6f29eaa73fb772e6d0c418183a07f82445223ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fd4196cd3b5500fcd84b1234e92ad9d422d1dc6559550130f036ec056f227a9da94fc8788b160b454057e55200c358c9aaf97459a5fdfd3366658c9948e1d9862ac6086242f7884b290bf0de5555ac149d208151e0327dcd9566e2357d5ab8bed2236c70bcc3b218be546e42ae5ffa6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d6ad54d28acfa92449bc06454b1d2303d456144943015597323dcac36fa5ea3d912af94e34e8499c272f257fd32eb3d870aef41396d1b7c385de6b376971fabad4a10993486b4c79afc9da2bafc671c81219ae80dae2a989d6afbe056bfc6c991b8bb5db301351cb78bc88c3ec168780;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e845b56d075c4a3cd0d2f63080dcaa28f48439866aa3a688f1fe2ed52e21d61601af4fe0f214a3a7c729c20ac3a6ccbb1ece5e1de293beaaa8e22663cc4ca694ca90ca74c6f11eac04871048eaa21d4099842c29df02439ca9b9afdfc5b93a907772650d33b2349e75e6a65065a51c1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fb749699843d59331215f611166d62dd9203bf0908deb0256a7c3eff24860281e3eab712385b1422610453bc21cb9b9a32acf67936001f09e9a8c5b365912c9c2da1a6e98e290c739c39ce204a3c506f7cbd7fb08dee742c3db12b56bd9cb130a3828f5e8c6859de96e58a5099bbdaf5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ba0a6fcfba001d04a184699ef8a8390b49a184e38470f49b49ff37119d692d6bc9c2b16bf26dd095b11424db960449e6bb3e444649e56656d1855ac9b45d8c890f063ab10a45670104082b27123f81f1bec8c33101457f5f57afd64f1d01af72949fa04955d6b288582c7bd12b0fa664;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8460d1c4d4800992d33553e447b6a827eb01d7c1a9dddab86cc77416a33c2bccb9ce62804f6397482e6d003b8dd9c4a955ef220aca21d9bae48d95240216fdc42c19c560a451f8985a0873593ca62dd19a881028d848c0a3a53fdff1b925dba012692004d64e292fd4a3555c51cfdec65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd498f38494d44e47a9bed76bad3a4adc0ac06633677fb4ebcfd6e8637aa763cb67da2834e14229cde0038fc53c329485f5d0e9069a6b211a2637c776eb1c5d6ff8b431a649587e8b160fbdcd72cc403d163b53661082d702909e69d8c8e248ab36d1bac47702f7eedb85368b719416b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ffbf13aa414a8a21dd3c9b79009afe95bc9dbed91263c59eec93ac015adca81711181e13cb6c7bc2bbe03b713853becdda0321b41d0d6a3868494bd4dbde25baaae20f7a582a0ae4ce7e15beff82212b0bf322ec21ef6ead41cd62b1a679a85c5df5957db944883c049bb3085232b68c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde319971bf83085792cadda12f9a8971979c1a9c927793e6a59d95dc6c1182df16ffeb9a5922b54ebf76ebc45c508cce7bbc8a4e8102a39e59d106037ceb08e8e6cc37846509514e8d415a0b76bfa71643daa9e365ab7f0aedae61b2148b1d763f636d0ee2d099e0b6ff62cb3fa542f3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3a1b33f612486edabf23141911200aefd25488a3b38d6671b46286f0c772850dc4e8861ec242722f76e27c55c5a53c3ff7588325b51bd8238d5ab9050d8145f2bbcfa8e20f6aebedc29c432dac02fadbd76eba889db8c2c108cb5658b74953eb38ac2a30ce70b1d4f6d43fa6d66e80d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d924cd489df2e3dd02057def03599a0880e26e93db83ce09b51c943b874a9d82d38b4619cf7226295d22beaa0454e58759dfb73aca6df3e057cd7f61dce6e78d85c5d6e2fcbb612b40e7c70f2e24ccd34932ca66dd82aa3f92cf530a9e7c10a412cdea7be2cfcada69b1c30bb095fbfb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15e19e7cb8803dfdb3aa67dd801415b36db6355319fbd6eb720c9faa3effd6534929bf74d8bf661c7e784f9a8782bf8afbe359fe47a5ec4138dd04dafb3877d0c87dcae5447c8b400178d8b886f73168b306437f3c906010cb5fddddfcc30fcaca8762fd863da36367fb0ca93b84e2766;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e3628c3b828bc8dfba958418842c033520b005faa0ae524d59c44d4121a135f4970646ac9abf3481dec650df4c687f2ef5a9afa3a8dbd48f6450bef3377903f89e310cd8d04ba153d30e35cad1cc324954e7014e59a50fd67b097ee6b8f39ee0a1699cc177c4697609abc9b76d13efe2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4768168006b44168d8abcbdb38758c48ec40ae4a416c6d5f25bd081d45799135ca5b0342ef14d2ab7b04ddc907ef624efd08250c61272584acb77bf6b0082e5d5d370420b59e8761aa7af68f806b51367fc7e9a945601a12c74cb29b2ae68de011517c4f4b74ab2f1c4108f30740bff21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7e980f8bd9acf7b73cf495937f38d6e5cd89897504abed4b61339f64bfe8d07a00d9cde287863b87f6654ad5c64947abaca687591b3bbe0c41d5d22f46c9d72078c24e1e841e41b57c6502000baccc4ef758469a3528800fd41135c2fac033283abe8dc2c2e235b79595baed6cc5fb8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc037423e102cb3cdeabc58a1d4b8a11715dfdc5a63d3dd80cf41a72f9fa1804218bdbc5f36fdca71a4befcc7794150b7c0b3caab32a6c120a57a7b2e630b3e0ec65c299b5a74f819dd89dc036d2d906e9bdf277085b643e33584a25c72317354e23864fa12e187e5b66ff351449d72c25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbdffe6bb93acc5e6d186cdbb0a74a33f1c33759f3fc98c91b27f8cbd91cdff02274e72565156260133d2ff6f463e5e1d7cabd112bc0eed434e831e15c6d5d274d5c6f4ce4d16fcb38a0062a097c84990f987ce0db090190e777ef48f001324406381e95ddb12037cc4ec2777d7b3b585;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb087101b1367f5ebc888fc343d613065aa127172696d1bb4d43cb2e5f97508b9a12937d048bd741270bfedf0243bd751c772d7280d7e22e4f190be4098cc0e768bb98ea01be86834197154e26c969909ec90aa464e7e6535da7e55744979fbbeeb5f13b86580c7c5395d91113812ffcd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9d5a3f84263cee4a7199c03382e5f56d1a5ec2f1f739051c61d01d7c3d435efa3e1b4efdea273c5a7a9a378594e011879c42c3145673eeee47cb3afb41a47e7091fab609235229cf79f00abd30fee6b599b3be5d94493cce2af58cbfa264d705357fa0daf30ab42bfa9fe42dc6bd6c7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49296acba626cc45f2b7183a7a372001e2bc2affc219ac273b21f45b7fcc35bf2bc585cc89be00e7fb6885129e037391075df4748470aec989416945a897102f71d6e5198344bf0f74499819d68a69aa6fd400f189d9f6bd82f62fd38e5e1b485aeaeb0372832540f86204e165d9b562d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e86086445dbe4cf4f6181e106a103fe61373965e4d5ef17b812fb9f68e0e08b3b50d472e0865433ddd5aaf1464715d3e323e311d2c8f38b3d6ee9ff747683100533b077321f050d96a341ef7262ec28cfb166095f057c41365122740031abbac70c8ad25a8bb039e97237d6789cba0f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbee7584fbaa662755bc85ac54749f1b868360b64fe169af12b80e45b8863abc0ffe3a14c319de52b1b78405f3dccd317bf5e1305edc11c81a44a0d879998b76191df0f0b61dcb6bbc3ce127c5d7f85642c5415c5e7a4c4525511e9702b85a40d2dac840d60d62eb37773bf5b83a2f759a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4930a754130ca6037df794b2d76003727a06c40ab933469f443c070b892757de4d0e6548c9f3d87c47d70a73b83ff3855de784b3b1971b4d00eb74cf728476da122bf216f8ff5ad5b59e02b84d761d34ca7c47b6d2b0d24ea8029fe53d0c9772b6488539555ffed9cbc97f86c5612abaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ea6e81c227bc88885e05b90cc5d6d17fbda7386279caf5b36e784c2c34efb05d84fe51320fa391e0129d71b3a53900083593afc74e5973b684b12a72e14b2b9be068058fed74383433bd01737fd1b5d7c8132accb766ebdfac1de37aabccab19164517abb9970e144da1aedb3d61802;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8b0e6d262a1d67f528b9c63794d517ec9ce8eab4a586e8404369cb490b1667644bf2ebb1821b9ce9a0eea160fa52f956cba7fb8c8c985fe5170dd5aa4e681c17a30aebb931083032bfa6886f8571c0c6a090256831bc0084093e8899d5484557a7a03254f3f9f099b6d7c500573cecd5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99a3e48e26644beb241ab5d26995e1e309713591e92a37663d7ca5ecd4e538eb9c6e7a069322e44e900fdc1eea81badfc6a1e1ba2b88f5b678aa96c5b72327c287e7761e4a197e2ebeef132d57088918085262407a98154e25ac754f12204290fb71e151ca8359f686d13ade94edfd06a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a9701941f45766c4780e1d961a5d1e7bdfc2895b4b71002daaa9de3d7f76f1140d580d232938f507823ffa95508871201c5de5bcc945f08e23a2a9e974f692b20f9d7b92c7cec5afdf94d3febca8271e062999db138baaa107d417953e360bd343dc14526c3a32cd511374af7f3724d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6952eb899314a43af8a03c304054da8cfcd55d1528aae7033d91057ce8cd8ea3c4c661b382ed708c07c70d6e39b6d4f5ff6b0161512a47bc0b393d8f0acdefbffd0feb985dfbff202ecea42dd5218ca292a9feb7a1d517e5478f0189e403e5bbe4462b5c8c368309e80cb357baef61580;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h393d5c832d9178f95c51147b1998e1d9fff89a9324d580f4c272dd865472bbdcb6d19e0d4c55c1948d8e481b55a7c76822207239bdd994976cf31f1f2e86c5260e702453c73445976efb6c8b7d38700997e0e7b562cc6d66e1b3e2a68ecf6dbd11956c6c970412c1a8bc2a11c2112f0d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48d20f56379b043baa7fb8d41b94433b02e8a127f3f03159beaee4fbc7784a8a760fc4e8c8aa97fb482bd8ec58863df8683b75bc215be028ae0a7047b89a244d84cecfe58fa430bce917d52fa88517f19fe24aa331fd6f1ddb67d16b059c32d253d4734387fc933bfc9a2da9cb7da1ad2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha648fc165366372e7f24c49cc0ce2b12dba0f76fa13337e1317eed338065f632ae7714a26ea59a2fbfba8301656a14e410a481304a5415929a9553f2baee298ea44603b49ee4bf2e907fa12a482be8bd6c2fe42e552d05a7142470a21f2724f5cd10cd61feb01d848ac4e8647f1d68ddf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88075a60b754f5c1763f9f563d9678164374270f1eafae732edb9e3c67cb05bd887f9cfe2227add37c65c12b034503d19e61ca9b66bd7e9ef0ae72ac02caf1fc5ea850f012b7b76d2cd4a1600a1a3f849313103b4788e5f1fc190a44bbe5094774392fec88c7407a817bb3da38338570f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25b799818f1cbabba8f94611b4289bfe5b9ba6ff8072fb9854b3e16f8ceb0d1386965df433f3d600d6aa3cf5506da86e19891da929026b2396db806bb49bf5a3035235d978a4ad9b57ba5cff91d4abfd49f20e4a43b181f0e10bb84ab98bea9bcc3e581587e2131fc8eefc1e7ccd09a06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h416763bc9fade547c5d5c379794c7c5646c6a4559ff1a8215ed004a5bf8abd7eeb9f718b1b814657845983900e67512cc357ad5db08ec2ec406ba185aa73bc53b4dec8956efe8f16fb06e4107a554b3df980987a6c71e46c2c04bfb9779230e0fcb8d23d5b0ab0497df05c06f6a51469a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9a74c8413f3e2e10ac13bfa8c827a443b6df0eb9b156478f04255472f0abf2fbf6a868c53dac9e2ef4277d6294e615f56297174c8dbfa3806cd05f04151e00d655a4d78707cdb890a56776d9660ff7df92569fbc9a0662eb14784ad0ecb09526cfa78913ed3a4bd0da3fd3c62d0dad9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had851e6fd19d96c5a0038dd39d669dd604b2feee999cc719c310b5469eef0e5d686e3dd2de3f70fa5c58e4ad85a966ee9578afe82143298d9c999e44b8a6c4631064d32f0f71c2c2e1155ad548841dcebb7e3c0337ff03287451040b285ea9734976771ca2bdc21d2bd730d1af184c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13f6c765e0ae24bfcd06e6b00d7a3746cf29d1e0c44456bb0ea7918e905c173c77fa59737333ed9ffcb8f92064470ad928e802739d4f7e892b9c0eb46fe513c1882c3e76fa942473e99054a345df394bf5c9db28f5db751d8edc3662ebc9af6a746fb6768111ec402727cc003dfd3de35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha496a62b2db8f1418cd8872377e1f7877448ee07597fbe8a95fb71733f0293ef9ac3e1fdf4f460684a030020e14e5cd45402476a806e04bf2479c38c15eeaf82ea0c8d5dbcf868bdcc508c3f5c27bfd88b4d3bd6e8a5cf744ee54e4b7319b246fb3bc68931947fc02b2123dc72d520704;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d8dfedda02b6b695b051b983ac41989b937d40921ebe9dc863a355740f1324abe0e69dfe982e4c9c6a9cf7de548d71fb1fc57eb90da86d703f9bc7765f88ffbe122c5ff52f074472ef14932c24da24219779914aa683556a4a802d184de455e4f75755214123a728389b3d12eb9910fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb159bd1b28adf4e8edcdaa35d9d86445d8d09d620409fd44d4703a22d66d50fa6381d597c03059c1f8052f5b53f699ffa51c63193a83a1f32fb9fc816b2341f9fe118c6295125b5919a5b7c90128808f57ae41f333495418629cdecc3565bbf1f1853447624c98fff22714983e3eb7325;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a33f23afd179ee50f721147790cf906707d2bf2a46828cb4fcc4aa433e8d7d0be649467fa21ea28400d3f4616e05f5acf33d858cc96ec80c9da35f99785156549293531880d653cc6e63c74402812cd3332845afd04d88b4484a407cf760ec9f308160c2cbb72eb685a76ce4d79e6795;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8a0f8b90968fb2af5f48759f4e39685e8b55d750cf61fdae672c9baba9b73780f2ebadeaa9128a48cd322dab92a21f9d5131e261ef334f6fd4236fcdcc0b03cb44b99b315591fd6b3bb6a9e55db54350ada6153a1c47c1b7c0b75a2d9167d1aadb403dbf4e2ac9d46bc87b2bd5c37cf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98fa52809e1d9327f9a7fe2223071ea26832c8115618072eca776c37562182e497003ae1e1bc6676b99c80a0551e3e4bbcb725bb348d708a7df6e592a0fe23da6b2da6d4a2bae3dad16feda9f41cb811bd8851e9b439b80c569df5061cce2a9fc19914f0e17f11e39f0b4b3e1635ba135;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb03436a49bc207507d095c43212973c202caa2177772753a7871c5ebf965fa79c1fec9ee9f174e3232498cc0d83ca70f86deb08be4e8a89522c25d9a3992289a028b4075f6b0f5256ddf111074b1068542940cba450f21e489e0fd72becc366349c41d335ced58b0dbc38987276527b04;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1194af76f543b2f96ebe3384767b93f5b86f850e15294b0fbfcd1d59b8fefe6768e634431d9b171087c1c0d0a86ab92116eec8616006b0ad6b9fdaf0e3970465f70c834d5ebecefbdef2817c0d0cda5884829be8d33aaf40e9cbec1e42a3ec763ac4abff8d407a3b7554f6ee951f4d7cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ee619bb4b8125738906da705aa16132e21a1ced7af3b61631af401d8af052ef56e98a4b7e96e95570a340f709e8a1e459037fb6afc6cbbaa9fb2b608ef4f7caf0689e172e389514ff5a68b64c92910e4557a2a25e3c57db56004df6b7381d1c8d605c66bd096e214f5ca3ab331a8bc1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7440e66286f269e8b45533b861e81b23d5ebaefa252e277ce32f4d2e535a29677906c86b9d0b927a6b1409fa58c49df8ab9d19ec47262467507caed76cda55c0003f961fd4e104c11f35cd9163840f8279bb3ee93481ae890fd9cb0969f49c7974cc63bd57c54aa51fb0388a414f567e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he278c675698f797dbd1a10fe9b257bfdea125344db88ad9e7fe5b049f8482d9eb8fe1865cff2d95ce33ef3eb7e40c87fcad8f63b4e1322aeeeefbf46661547d662814bb43291d0cdd13b106c624e68243154ce13d02af63f9aeb4facad568fe1a27cd1daa532782c9e0736cbf6bc6b122;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdf16380344fae320b5916f18b0898b6b3b3a016f3df68ff3d0f063c779937faab42a67d6b3d31722e1c73b542a7dd3be48ba6c6982f26a3674c078330a9ec1f40522a73a4af3b909747d9ea163aefa08064fb206e0777b7dddc28841a4dcdbbd764c8feaecfed3ffd8ef97041fdb2672;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e54d42b6efafc664c2ba772a6247f0813fa2a476d269559c3fa2ecc6000df867b4409f1e887a5dbff296040c934eca0469e2bdd3092f309c46381bad378875d3895d9dbfd0ea1c380d673c6c2871dcdb027f9fa6ba10f80c05b1b030c4a223fe87bd67f6511d4ea99f0f3cdffd1c2f63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45aba41b93c45590cc07d38a38e460bca4e4e4c914b058e13573b2da71af8e9a014da28abe24c362104ab4c9293100de997c0a6556c44ddebdeafc98a3b3a9a8cbce87454ac83ff75acffeccf6baa6b311f76803c039f172cf60ae84dd77844833947990d0d909ec3f89d33d634231a83;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h729819950e8d35bc9686ba316179a34859adf7d48ba22ca6208720628083ecdef34a8584f5e5dc4c0e16929f92e20046b654aed9cc1fad90bf57ea6e811575e0f6b88ac6f757d76afe444d330f2cd077899caabd8af88eddeca4034252d60ea8281ea53b6a69d3f8ba3bcafea14336bd2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2c9515cf25484943961d4f38c3732c36cdc0983931306d5bc1fe6249f4bb929b118818b7dfb609f9b877d08e8a8e3970232c65df3e420faa324418e37d47aed02736907bf48bbba60d30f9070a7682d41654e74fca083724668247fdb4606e8d4bc13b9f4747234404eb64249cfe6fe3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4417c38c5eb8e0ad6c099f209018934cc9cc4c0c4dca6b1f743d1679781af712744b608d9ab1ad9faaf31ae280cc7515298a91affc0d065f238ea37d7e1ef9152f0da3d32924af0cd8982ce2623e60c34ed19104cf77b2b7f991236463d635d0a3dfda18f68380d623b19af651155544;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had2e0a584d751d275f8377f06f8462b7718f5da6da0fb137ffd4e40ee5ccdb4bdc516f38cdef76573422bbb7b8371fd6ebd1b469fc08e1e12d800a2a792f0cee715cec9058d8a295e6c13a04abf66428e1422c718aeee26b11e4bb0392db17a4ad3aafa6b9d903b022d06d74499ac1eb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d6bb81e42b65e9f6d4d2ae0d2b78395b9dd7ca35830027179108daade29eb73153d7cc25c84eacfa78c2c14b6fc582c72ee5d3d446a50c5509aa2584c8071b1951326628e0e3ab62fc5e89f4e5b1e922ab1ada968fd31a45676e72cf352ed92c263d652981631e1b0f721fac591b3702;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a39b841a6eb6c72958d7f9a67e91ebd09817296d7410a63c4885ace14d35bb967fd04e2f87e20642eed036a52e5f91c82a905eef911fa81a4236f9d3cd95ec68e96ece0e84e7b23d9fd6a7cc8f88d237c2c2fc80962da516572809637579bc48579399ea3938d19156a903365d3e6ead;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56ff4f197b895d9979fa89c80578a4934a29511f2bee12d20f036296eead2775600d58c40f4cb6a3ab410d1a8ae65f30b9a5297a0d1144026352f5c0765d83479d5f786ec4a8781a08f2d39b828724535a306750632e2d93509ae2e8c66e70996322fe6ebc80ba55890adc8fef0c4afaf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h885b85f3ca127e7e067a3d8f24a9d65b9a1e546f3d2c504b62f0d62105ca76f999f6ffff6c1926842968b87bcb63a9a4b333e90ddea0e3d2b5cfb02f269ee121dabf81c61c5b95db65822ff50e9bf010fdf76c13f29bc6a824631034ee7401a92401e7c6c4a633208b14d8a6b23e08508;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e62f8ec5266be147d6581e2f39f58b65fa1e86f7a905f70b1e397d7eb6a5e1ae1ff3763e0b1102122e101cf206d77882b3a5ec20b69da03643a7bdc05bb8ba5cc5e6795a6674e93b0bb287c131fe1433f3576d219f8d6b0a65011ce45fab54fc47a89ffa2075092ab103c2ded892af6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he83a7d9b258b279a96828bc4b2d19473a1feb6a5362b47d1d672975f04bcbaad26fa645941bc8ba2e46cb6c04004df9e2947cb697ce9ccc97d88d136f95338b94a260d0b66588a77baad77c9bb258804891059ade6df2c5bacc1bbc755666b0bbb81100bf2ff9fbe08e1853583a7df073;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd42fede4da174eeb98b5f6d843687ab34f19d41c56da2e0533710c8456cc5bc70986b10cdd8e5122456b8cb742fd8667bc22f279d21ab03fad1426866ccd79deaadebeb4d75489d6278ccb61761473d3da4fc0e6305bb204c4a4aa50ccb9a6b678f269b91d601b5616d3fcebb769c9e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65dc40065f119754ac8b9843cb51b18a99c6ce033caa25c990b24ba0fcfb4f7a36dc3185ce53abe366e2818346797fd945f7f2469b9b976b29259e6d635e8607eeb1cdc067e9bb7c54f2bbeded2b988e69f58e1713d0935922fdea045fa8b14099beaf1540cb3972d643f2dba0a934e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4406191afa1096bd5a1b328c959310f29608b0b6c3fb6a9996ad77e5e44ef877243ee9722dd9c7c69d8abbc4806084c219e8e4ac198970b7496f7264c1d744cd34d2df9c298a6540fa864eef456f6da0c240e5b4b1c6e530c47c015799554f8c4bd9d0746588e30796319e044ff91448;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8ec7107f11593006ecd67436ad20033a2ef298287b6f6714ad7021863743e02dd990e56ed5a8cc0abf477e0df4a363a69db3dd29e346ab1de9b07d7045cb2ec917969cadcc26d994b4aaaaf9e5cd15b8830e1d0c89aba8cd0a89a68b7f6858f29c970d24df92df905540496e9c11d4b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c40b857776dc4c70f39fe4e3a522fa7821ba3543de2cbeb4c5dc1b1f43c208ab46df47a50979de348f987e6833b029951ef49ddbc6e9abe02b1a62393027f427fb06ffc7dcea393459165c4d2c1dde74f17d0d3bcc4b116f091da3ae3015dc90b6131d317946b596fb176a7b6b7fde4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h416f5050440fcc0f843851aebd9ffd9aace23609f8a3c020f396b9b6c7b7183552235792dbaf643fc6f7b1593d540637a8278a367ae9b8d425b0702e3ca5b188e5455878506c4b11685cec6764151ed3a7487ffce31636989e819c9d68ef02f5dabdf8be2daa23b54f5650f2bd7b20856;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbebd614202855646dd9959d1003149a6ff5c3bfaa1ae55bbc930e05f55bc543197cd7d4bde2563b885bab13147f59fb2faef63f9bfa8d937a64f7bf281dbc8024e393cf91e41bbf435563f0f8019436dda6f26878d776dcc387c149cfaea896cac059b157b221191d91685e5504184cab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa4d640a7ee1b4756915003d166cc3759f61829a187edbfc262b5d59cbaa64ca6cbe9413078817a07d323dce62bb19a586466973f3a96c631b29cab872b0dc973a0fa2a0ae04d3a1fc32ba357628fe603532475d472cb402f5c6af4947b7606d74913ed0199e1e57f69cd691ac364dcb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa06c3630efb033d5c9652019a4b85cf0ffbbe55a69aa57b875e520969bd82e6a7a02bd3a5e53ac03455107b86c284bcadbfd3c9c08db9586b27b51066234bbcd3cd6634f4ae746940687081c36570e96d4de34b9773ba8d877a5a01884310c7c8dbd6da81092e7dfc191e0534acc0b64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6daa8ee9c11df44b3a3c58765e3abe1bd7e85dbce372420daa02392d75896d9215ade2a3ff66d2ece5b8924acb137561d798ff8edaa401f41b8eab7ac81c6e499ea93f4d9a0305f606991314b3556bfd771be605ca41d0869435482394a34f8a96efcb1e5dc9f13fc74eef9f14cdfe0d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cedf3714b5ddf3c34dc3abdf619676617ca38ef5c31c0eeb922609004972901f40e3e63ac8bc249d2b28593afc83aa5e27d05649baae0a9216b9a349af23438332c8aa5bb9dfea2d9aaf909955e25a06c5f0137b08cf527e9007297cf7a9f679a4f62148b0f13aaeaa9dde39ceda9b5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79fc032b62a737bf58d052a4b5edac255546a2fe49b73382f7e24ba442cb2ea95277a2fd1d50bc09f25a3f7da9ab0dbf9b6a07b9fd6a35efe044c8304b21d1da84d4771ced42b18d03b5582c19f2ca2e74aeaf8dd95b6944264ce31b9e122e59f8c96feb3e3f669d487bdce2bd9db9c88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2290d6c370d9f17da16cc830914c4b22f784bfbef9f0b94a4d3133e27e741c4147a0659dbf4b78c6b8c4298fecb975a21f6a64e843117067189808f8b662e113da8ed8621c65e09d6d105d201b64dc05c4b867f77cb6ec6fd07b17af8f29762b013c971b96fe7f1ddb6624fb5fb09d056;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1556c219b1a625bf6c4fd9737266cff2ddfca289aa9e950f12e51bd8bad1345796f0a1ff8411134878088ccf045ccefdead9c59a7df5fe5040178190cbffe9800b23c67de33ed9ecc4a1a663134fffc10f4ee212b4a618a23204303176eb1221a77178bf5eaaef30cbef55d79c94b3de3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda33b4635fefafa317463206b59c91bd98f6c5e2a57dbebb4cef23e4907012ad40a971c9cf840413834a2bd77edcacf62c8d41adb54a63eee13ed8c675fd5bc23ff2e0821b791d9c8a21612032b3e11ef724af5c158fb63dd9ec81fcdd853b150874b9ab88f5579a5c79cfbfaf87d90a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h903f824cf14495a4828e1e200da157794550df066c53087e960f61c37f6e02f35e9eac638b33118fb22246f1a58766feaa77ac530d2ad206cdc9851bfaab0de741e3d6faec7e31165fe9d34f5de7d350d60306f74f16a029b0e560961d1305dc2bcaf777cf7a5d723dc004899b498f492;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ff82c83a12447fb99954a9304bb578a304ef2b4c08b5336a87b01d025be0a5074b407cc6bb3bfaec6774d534dd5566ec4b1e4b9c080e44b7365a51dddd18dc0630502b15e47eb9136420d930bab2ab25290f644605800863b913a588ba7244733dd46d33e09ff0f68d9a2f9a95effc8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a6bb550905b76028c9c7b52adc85ebd89c0fb3e819749b881a8b20862a348083120afff44e7409b971e42d375b61aef39fef17c0ece41b2dc33b2c18fd8bddd9cc2ff725ecb918cfa97f82c1e0c38cd90297ed1abe2ad1c2ddec81bed7a8d633b123522e983f28b69e01257a1316b724;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ff2d8f31874823333ff31cb2e4cdc2c79bb7e79caea9c83ab362f131ef2f36cd3798eb17b5bb3e833ecbfbdb82c016ecfbf591344982786e74c887edb3c4c209d0f061ad6161c2620f8fb4e5f445d1aeae1886f2147613572627494a7f6c3be1b741b83158592030984e85ddd866ebc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80b98544653d39e1140713634a7b7ba5f4ee8d2ddcde64e18176f075d7eeb22a253af80ad266d92d11dceff6e06ae7141b43b2501a90358d6f915361c26b83cf11d61792052cabb979825f77250276a0fb38ab121be5a92a4cc9c0285768aee41f3a869503bb7cf60a5a16c983e107968;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a25129796a8982e2adcae8ac2f05ff150b5909c75e5a06cffba4684f416b058361f13682dea193ce3989bd7d0a53bff78a7a8a2033fbb00a1a902c8b0c0b51175c3eed8abc27271b51f5b413dc111a69cd6d1c36a537c95bcf4fbd6ed6e5480478c9b1218d3c3ba78a783802ee2cffcc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb30168e61c65c655ab7eff57f321fddd0914fb92a6af994a5725d75662f134d96620602b98551a278eea54b43b91394077757eccfa16933326f1655a81e8739d46e9b6243ca3b27bcc7a8ed78cc00af11842398212fc9ebc4133a70c59a6a0eb67c5402974696cdd6c523f562f220dffc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75f5772b557f29ce30bb5cb5549fef15370a0e63340cbd721c378878af43e0565e8d587e4b4a64821a90886d8e67063e8dd879bc1ed040289aba2ef22b750a8484c273a40da85611922deb1c8988734498c47b3e33266d551ced6e39ff7357e5ea0e0603b2a126f9cc8b8b00795759416;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6c5c44455b0aa4017ebd221c72eae2831cd5beff18f71c784e3e0cc70be0bae96af4c9d9ce5caea5eb5d5db9aae55e68775f20a2992bd1cf28c431dac3374e1eefc864b0f8d1cf8b1609668c4fdbb62b3b8a13031313303e84f5546369b6d7cd1564026fc166f22893716f089f63e218;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd50c081261ca36518710a9402874146de93d63cc84f6cf587d191c5e4e3cce6b08bca5f169a82f13687d377bba631871034d8b0aa29a34b9a2cab89d62d3b30536b62ce291df5e295b4d9f9637140ab4e3d61552dad6e0e99d288c919f99be28bbf830d1e93f178a81daa10387f003a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d3710d10a18b2457286d62d4e6e2859439a25eb568338f0e32dddd56ba39068a8107203faa8f15cf39c63bdf28a9a372cd59c60c36b1c5ce60ddde7a7b9c854164acd69abdbdf554e9cdf5492e8fd2fc87e3ca737dc7148b2d2eedcde01fdd771aafe4cb5bfb0c6840945e751ebe3206;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7db1a26ecebbf8c8169a0c9a9d9f663ed31cb43d140880311aaa5746c50910c3dad7acb03d9685a78d2de7db4194697fa2748c7e2250dd8e34209c2ffb690b9eaadd168cad83aac2336ce8b04f3cfd40cd5c10b8cb6f557b3e6678ba482ebc764a8cc8436b7e3284bcc27de58992b16b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30e41685de42d872a5dd9a88101af1d84ca7e74956ed2c13d6ccf492816f9011646de44b97a13b64dbe945a8fac89d0e56156daa07a39d83b7e0fb9eb30824452e66e80e4c770723aa39b90978b983f6517fe968cd3be12b3a91ad4d1cec26a4844b2f6191c39874be2526e8b91148ba2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17cb04e9b507c970b759bc08498a6e021c9c22f10d0f8fc537f1d038b95952b899f3ebfc0b7bb622c4438b3b0679557c667604a9c42f942f389dcd9b9a0702ff722eafbf3ff8a5a7a8a470eecf158041feaf0b172a9ab81b44a5a24de1f2fd265b37265bf8ebd7fb7a256f8c168b29ef5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had844fe77ff3673e369400e4f5161f9c613f7f58db86fc5aea50b41df87cc3cdec71dd4f6aea6afde89bf76a5225f11883a6736e778dec5c40d0eb9c1e67d0968c278a3795b8d60e1565421b1b057565130b4a88d129bee948924aa14d8962e864fed3d637a0295ccfb4bc87259dfd34b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e87d583a942f3a6a5d7b2bd9733a7ab541780da0ef4d632828dc760c0242ef61ba3bbd40eb57320730fa6a930ce4fe80abccdf82c8e4f29c2b81559764d16aa63bd7c4e09c78525427533a2b2df909b14741d7ab66b902597085a4867eaf1f805fb955262313f2a9ec8837c34c73595e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b254b239cae6732c69ed4039b8146fd4b9069d6ecfb2d9c6d0183a1e7ab0c4bd0f292c9d4cc4d9de44becb345b74d3f790fb09e87515ade109f4522100f87b4fc570fec859b571239be79ade8fda13cc4b681390dc1a417d847de1519ee380355ef4bc2bef23bf25aff87b592ac7f9a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3ee5641425f0fcd0a5fda0fe247dac75d77984ad93b4f71830fc0beba60a16ebf1628c5a7b56fc281f7391518fa94e395b033aabe0c94670f60ba6d3fc51bb714e97295ef3a1e7bd1b89b3bd2209bdbfdf7ee7e28c624508d404a6cab91e4bf816d963ca97f3d73d1d4762c86302ad65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5992d05547bfc7d0aa99d92a8434bf23ffd1809c1104d66c4e0362b30f60182f895241cb36468550d895f3a7c99a05c1eb9940eb2d7f8f4a175d1975455c73a925f12477a83c81fdc779a40009aa1e5064e024a5cf67a24943ddcd474f480ecffe31f409a1bdc9d29a842bb433883b0ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5550bcae0bec877e6eec037ec5dd052079d17848265fb5e81b2e664588b14c399350ac436d7214e3be93e19eae5ed2777a5bf08003b61a0b96cf847ffc6a335f9f4c30f2f957ae6602d8d32b85f247435a9efe0e245f068e116d66e3a9cfeaaa46aea0d10774081404bf4ca5d8251f02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc868397027db32b48858289894ac225f4e714a449fda250efa91208966590538ba4a977665002bfa4fbf4541231c3728c710e10d4f24713427b573f5ae27d9ef1d08d3a6bed86b3fe532529591c1b8d60d6b0681524b3e27c671bb0603bed0f2c7b82d6dc83756c819f131c270bd2dd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40356b3ed4f24dba01f1393b1ffce81737f30ffee60eb06586e3dd4148b8e9900c6131ac45f3d71436f448325bb5d0247c220475055936c56db3a7ad007234a0215e2e09727b94830f9c1ddd3dc75ceaa93d36a6a5d04a46399f84358285db43fb916a5f1077c51e4ab094a94c8588b9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a19d636db0ff744aff503c2ccd26cada8df673d1e2a0233fb39091ca86efe57a2c76d4a0adf88c43c026f5db03dfdec83946c05472c7f3b56db839ff2312ebd75e32d4c426d8ddeff83fe254ed4b935c4b28df6268d99153370cf81eb594b101dce6385d2f01110d46ccf58b2e2ef20f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69a2ecc252f6c00081c2c4231340e891d3f3931becfc689bcd3372c44212ae48a0b7dae7197d9ff10ff4f90f36e14ed1dcac83ea23cd392b520b84c749e922ec7b7e0260dc3259d433a424fa54414bf69ffe1127d587d60f6584b653bd9d4ac9b4a42cdff9509e0d0c8395f336b5215d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd16df4121bd89605299f7656248b15531f326cfdb61046a7de7af8507be1f04a010b391da89d52b4234676121944cc0b85d4ecd5306472c7332516add67e06d32910104b9714ecc1b9f04ca9610b7667ac0aff05dd86158495afdfea987709dc13db45b844c93fdee82ca0709b8644f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8c8ae68f89f8c8c76d2425131c4bb5616e8c99055138978f515b926fef78b01df935b34921702baeee1ccd0acbbd94a7635d83ffd8c6bdec07bc8aa0bd5e9fb7f10d9638ba1a473b10a5d790426d47ed7267603cfd168c726c2608a245d782cf9e0f8c7a24d48ae41c09e6c99985da00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he02bb720be7c573cef7261c8b1ab044a92b4c1d8e5dee086172f97bcef73785687463d2f67d062ebbb0b4544a45081f366cab7399b6d67c2231be1759b696e41153f1867379635aae7cdd3a37121297cce85677b93e59faec3a8aab9815e86d410e7d13c1012123517c8f03769ae97f51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87547d8ef58ed33dc884d9e7f0a039b352e02dd6fc69f3f439e3ba0064bf41477d7b8cca74cee3e0bb8cb718836b274f4931e2b7f839d4afb146880316277a0fcd50011a158bbf7e49eaf8ea9bd687c3a01ba5be7ba9f89a82cba6de81a0a91480d7201e0bd88ad6634b6ba4ef9f84a1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f03ebb301717935504b57abe868c68ce47d8fc216ccb93165bb05de7f33a3875b46a8afb12cc56ca2567906fd47bf238c7f76aeb114c77536f7dbba4ca5ba05541c3967ec8f811c97c1c1e0827a4d3c774259ba8e448bc3c7ffa9ed9bc39c7c02d46b99128ef02d43ee7040156320741;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h786668c52cdf9f8bc55fe9aff6ce257bf052b9d3a55c1f971ba5559d30825bf03739aa32b48a7c6ab89d43abf3a0f285e1dccaa9d07d9e50224e4642ef846b2aa3c8c9a892b58a95d255fba8dec60fbcc8c836d96b9af5de306ef9af189aa920df7986d07228532ea8cab87a6270c6b34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b5ec2e81734b267bff6f06c79cd27ba0f71f11c239f1832bb69f56acfa32a526eac1f369261dc2705883b32c9fb30e393473a922275b6b00a038a345780edb095288927b6c9a567c5b8668492368da0d93298209dc4b32de846dd13b925d95e53736e997c2e65f5b4fee72237f73ab5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb64b0d680b589605766457e64025f22e26103e26e963d0a34686309c9fcd95271daabaca7fc511566ffeea98faedfa1e15be29234bcf90627756880b9d4f5b1cc2ef1161e5c57fb26ee17356eea7685d29059d91826b2edc98cfc003d241ba1ce01bb2a511af9545de664fb8391d12fbb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h480b0330a33dee633025968febd6dd94fcd4aacdcba73f5fdc6afbd11bbc45111589112cd58eee1b181242a9030abdf062a49ca5d92f029b0e847fbd3e2974619c6eef110ec042c578d3e742c7685820941b3d9ef79118b32ff0a88fde74bf0ad748498c32c5021019b8f741ee31d5baa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a4055a58f25004e0ca51c7cafa4e96fa892c941b0d2266e5db4378792898a8a9c926512a84defaaff5177222a4ec7e6081a5a615977fb11662e520a7800d79844c43449e69546c9c0054cc944806179b60c3e1bff09e6e17cb399d2b6419cef82eb44381c57a19287c7e5784fd976e99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he68da819991c306832d0067dd06f51d786e55389999a2f01532dd38caccaf638c61416b6a1b69a8a4a901f9a505ab330e29ff3a80555dc14cad0f1cfed913539d230b7d638bd8a4fb2ab9c27141d8e3ac13b15657fa57ce08a100b562e79257a538489bca100306f073447e1c3ece6536;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21b51862a8542bd9ae463e99083d6d7fa861cc9a1d80f6a0ace7358fd2e801ecbb46c4d5cf9d613a80f3e204f248856b188bce8c06c2afa1efcb5f43e3d34faba233e493cf87318750957e00447d67af932c2dd6bf475c98ede00b3487f671ef16643633849b821a42bd963649fe512a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbedb240e042018fcd46f6b386639a438982065e4bf395221b15581796ba83b7e9ee0513603496e52f75ab7e108ff05ecc5dba63dc9d41a5112b9109b90ac167adf1d45ecc4938b1d0207cceec49089e2d2c3865b655f252d278aad5aad63982aa6a9d0e02ffe34467741f84a66458580;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9301864d636bfd8c163af52acb1c7cb0af29690ee6e906ec8f3bb9f0e421329b68ded1582417c4259aaedc88ae385ff10d9ba5f9617a9c9c44cc1ca322ed6b4ccd995c9437ac7d35f29b3db642bc59fcc02a1edec6f47eed9657a3c310dc87d637304f22dba861a22d4b34bce234c87f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f039b67c9ab3d6420d6bb58e79993265a46c14c07d63beb59a07f4354ca582b0103cf61cc12c08c6468fe2c584e5ae7424367de2c9c7cc0c887d80bccb1d11280ebb2bdc8ff24993ee26114b39771303f53b44c3de7e7d544a21a0b404d98a1535db6d0e48c78f6083ab58bee68a764d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2dc3804d71fb7937e3c2953da81122b40ba6b01bb324587216af8ee737c4b026223dfeaaba85dfd2f9938d098f07ba8ec897e96ff75f670091b99d6e411507d618bc7cff367197455b4b62a63b7234e470ac728e665d7ec4929cfeb5c56562ffdf898a49eef94c520f3f54bd79fa861c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he515fc720372140bb90dd7b5f8f6851be7d5398cdc462c36f31c8d569138e5f5fb6812aa8579c002f2dc07e845baadcc11bccc4359bab436ff507414b18b745f612ca9b59a8087ee3b2a225db894ab55c066dcbe161ac85b87f679b4c6ce53dc2a012cea843ba5c53df0e023aced2bf46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc21b274f690055a355a0d2548c8f7019de5b68045f36ce94f06e417a8ae8bf7a7fd4b55787aa742356df377451c6bc19e49d32110e09774d97753f91edf67c8b9b048f68fac967773eb7757539bac13584b1791db7026883a60e01d3facac65d6123a3e9c7c0360028208908627206a2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd8cffa1c610905fe0701b376d6490ee7324a600603fce5820fcebcbe5b0a06e01b3a287e47fe8502fc5730b547f7cfdec318e1af6a3e0e76e08bdd2da89006cbed2fb93ee2052acdac7753e4c16c07910c38db23b0ab47c1e25bccef1c6aa9ce3080f8ccb64c0ea6bf26534f82717e06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbeca0f312f1f6b93f238280405e24241bef50c27fb3787de5f0740ac7dc880a49fdc887a5c9bb3fcc5374f2e8d7157550027ae3d63182d3fabf12b0bdc7d0c6be3bf89c3941e35ebde88dcc0423adab9c0dbc571cf990910ac950ad3889795e9d075ed463572b34a727be21765ec9b9dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hced7438775c16d0c4dc8bed2bc814fe2dc9b721128f67e29babad92ca1c209df99d3ccf6290094ff6f0c4e7a065ecce07cc06d64cdee62d0b32e38f9dc597928b17e5d2107afcbccc22021a22b4d043951e2b910d823cfdd8479a9deb1891cfbac0732e2d3415f6cc008c96c5a283d8c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42062ae0f0a9459ac7d144391c6bd06243986b796fa13deea0384ace80f6eaedf59bd073ad742071dbe029c30152cf3ba7f58780b2eaea9d7768be0eb61033f8d45bf2ef234810a985d5ebf608e14150e7cf41207a39c111eb6fd8a7602134bbe453d331aa834aae785ee71fb92f9e7d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe304a3e47a82bbec834daf1180e00a5dcbecac9c8f1cedb9b0df7f8334a1f5d649e324e2bb752911a08e313c83c2831879e2f24578e308a6923e2dc0ff9dc309ee10ec52ae16851f4c1c1c45175349a60eddb3c4d10f2c73af264020f87c3ce1b4b2c945fd6cbb18ec1cdb966819fd5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0d166d6768f19ccffb3ed232185cfe9c10ff4a32ca385363d2197482b05b587321c3e51a777b463c6812dc94d6fd81769684d4a4b50d2ce55aa83a6e9699506e071d2b599d291f4af379f0c0170c27d9f2127a6611c55c59c06fd99aa68cc6a554f0fcd7248230449c5f50fe388eb997;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he84b1ff6529b9d7dd7866fa3cc4f126003c72799a746c4e58edbcdec491ef8dda264dc659524ecb15250905beff69fc5f52e9bd7595fd5ce2e7b74c91ed53400003c51a98ece6547ce05a059bc9bda07ffe3cd5fdb428eeef7c79ff84d5758bea7d9e79a23b96eab099033537ec032c79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h694748952724bc93af4c56762655028c940affb4fd1c8d884cffebc5123a311b8052c76753a3d0e9ee569ef72e21b40f2db21d11380928b8326ec8629e2e6a823d4046a11ffa0f1fe5701a1863029f54b2e1d4046c2b9808f135d226e28af14dd311215bb8f5ca20a379f33816eb15c04;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9efb6e274a93676366415e250cc5f26ef1bd78d1aded5522676aa2411499c059a0b94f56ae4b4d0b4355bd83b5352e5523546bdb02b15bc340f1030d37376bc30b8e8e99c2a323e8bb081ca0c449f16feaaa2177d49b6c8f899a774a602fbe1dc312feb9ff65803ad9e57420a36bb51e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8189820501d85ecb6ba9d34857126abe123a263dca71852d775837f8c67eedbeea5b7b44bd33c56191da6ea823608d269f5e7a0a18f0b69aa02de1d5540b1b47e2b2537c7475842e491a19a50dc75189f40f30c8d9c23e4c58c54d1a1e045ad3ffc372030fd267fceb1b7ec2457fbeae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e58f706d32dbbdf1226d37bf8a7eb337d99dd57dece2f88c4d65accb0772427bc834798b0bb7fe043ac9c8f147a8282a9725aeb77f29d2c4b3d50a8bf4a3466c2d7978ffd4dfa862d9fc9fd9d15a2c872a613b0dfb533ba755374b384ada9703022bccc1528d0c1b797ae37c58750b71;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7899247fba33158a2594cebcfccf8d9726a6d7b76a79bf1d1e7f5caa02426a3dee830d174a35415dd61bf3b2cc9d4643197765911c83dad0d859171aef5ce2049603b75013073d483d4c03faebc6cbf09b1e27e8c0dfd8ef63d4ccd2f0e00a378ad2db8fdffb1b31b1aa0d9c5c59db6be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8aa0b76fdc1dfb41df7472722eb88038c14ce32fa5bd342d5b1b44d3996a50bdf0fac09063fd12d5e9b945fe1d813a577c2a5a25b072ddd4379d6330b0cc086f8cdad5fd576cd52bada3c7f30c11df1e1ffca7f3d8230c7fc7a88e9bcde51eb1d560435c5515711e978028ef73b9ae73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92d766d8a465ee64301f46c28251fcaeaaea9cbf004db9c415e0c83bd94d8f7ff726404a5fc359cf14349d172f0df6ef463f66366542d41e40ec751cb27bf8c9867a4ca63957a96abb6b94fdf665033f589177102310929db7da7678bd13c42e67f184a68cd793a3285df88b0f9592178;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d37acdc3600fac63452a591a998d5848114e6c44144bbfde628a8d9db19c00f8d79d965ac6f98d79383a7db4c601b55c0c9c153522586241651af107475b442e87df7d5c3ea0ff57bb4b6da2c55dc82127496f3b5895a243752954944ff26d87830827741432df94868fee2de96642fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5a87ee41d43d93f2b46f2fd32652819cf05d01fc94f05b26280d3070473379a50b19be67e52d64f2fe8796b553284a2bb3798e498c2d50048ab9c54c45ced232289474f2a2e274bb5ee20bae7af4bc48917b1800e8a38d0947bc372978d9fb07a80899dca5bf32170bf4d8f29ed1563b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba6c789de2f591427f424a2b91088c6d35aa38f77de62dde447456ad10fff72c59157cc9e8305ee6ccfc2d9824e338b119ef85dc486f91422228159866ff61bc5f1bb3a090ce9ea2f3f6022d733b99d33c5bc92ed4049b9d9e8686c982a7b79b737add83bc913d90bbb36687e0efe89a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38393bc3c20a9dedb3a7db0dd0d17aaeef903c0bc48045c2743949f4a3d22788cdee890c853bb8555d721cec16d37b45e71f7c702aa5b706ba49f518bc14c79cb5498a0e48ef3baf86a22e4e80a95bfd12aa997ce35e76aa36d540d60bdaadcc00ef2c30c46b6aed8d43547a0c0d8b3be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5565ca3280e65c34a1291f223505598cc3c9fd0570eb979a95e039378a904445a96c36f6d070eb1d81d1f59044a2818d0f74bef49adff0e6f3a24da0df7c156166926a32949d64e8837327110b83117b2e1915d2e883d0de1ac11afb94a1824aaa8589782181f25728a68a4df9e727016;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he603974996876e3a8b8b69e06e0a440d90a4c75b7f4d41273f7ee75f2ad4dcf06daa6cde9beaa44ac7ee2f5fd4027690c162fa8de7cb4955566c60f9437e5087dee0928e17abb23576e64b88b1424f9ec22f47bd61e84fac4b415606eebd786bb938f2c6ba7a13418b19371a3ebc50587;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e19fa6d6b49c0fd862ff49528d4740e1992ea8a6a0b5ba418ebf560683d7ad05043810ba3bf274a4c36f76f5fe4e59ab022f3c8047b6b2a15616908165dad38275452ab709bdf2c5593a08f99386f54acee6b2f452b4b03cb1d5ffa01a36459f4e49f3736c6a6a0c1379f8b2511eb478;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcee0fe7f267aed513f0137cebf9a1649b08f5c23d20c02600a9f582b4efae60cc610cd97dbfdda95200b1e9ad2c0ed612e1de7da72c49d9bfbd9dd6eb0e18ca0ac886509da5a0741594020733296be7ef8870ec9856ea94aa93403f4322daec763436ec0aba3dda746902f2243b126e4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95ef6d41372af74ac6bd3721e8eece19e3d0a7fe1fa69e35bd6ed95952c1f6ba74c878ea918ed33a6a229d74b8dcb6dbe6f6732c81f2427d916b4da2044f0cddc1bff9e5d4f7b6d752c93a1a053ef9b430bf8112398ba6948b41b88affe4aca75ce7d1a18deea07ce3b6a7bfdd8df599a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h177dbfe5a955017c160ca6195f256b09798135546064b9e766c173d408b469f3ebcb6ffe5735c835934daac86d5cafdeb0c096d83f157d49d06f26ade3c548efc1f990c92fa972fb4d8b233885fbee93cea06efc9bf2cbd180099d8d59382e6d2d5e7cc4f43a14afaec2f54eb62c9d8f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0e85893572134673c0ca5ab212fc478b00952fc1222a8d3a6605823ce5dae746eb1b3a8bd320a166d75a17d8cfdfb0357ce8ed8b4d067d0af84d260cd7bd7923a2c4e03918e858f3f2aa7a408b7c809ce48625cbebd26193f8b605aa902a00c037f63c21d29550cbd58d123d7699a308;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91922603ec683223ac3439483e428a0480c31e968bc419e3995a1773a5ec60d15a707e3509fb5d0576e79d3b1e007e93c2b0cf69651ffbcaef965da9e33ea54534d1c05594d17b06d8a3bdf4c2dcd78a58a4066f45b3f8a5b460640c46e685d589158dd36eea8be43c6aee76623902db9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c8eaa90725fdbd7370872e9efba5263450e49d626a29afd591b054024cddadfdd7e19fa0939193ba55b6c6d16dfb1fc16d6516a0fbc2cffcfde73c9d162a5bf085f760db36c3c04535a89875a3821c0cb5d16947c887768d1d0c8b1b791b8fa4525935f9ce13e05ffc6aa004d738b067;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f7130019649bfd54b5be92d7f5002aabc5c555a1b6419c97bdb1557b08ce6835222659678d52e71df84b084427308c992f3a49b0369bf3d3c36e1734cfab1b320e1e800057c36b2dfa351ec74e7979c9fc185eef5a2d09b1216bf40e09fbb91abd71b9f0a45de4b8651bb296d146a1ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d87a0d8165a98bf774c9be0efaf1eeca5fce41621602b92feab10428e2f371b7dbbdb6ac98f5124b434cd2a640e2b7972f0c8cde74c731964a20898535099373e2c9330abe9e1306b7c0fd71177c36e536ffa50d1a84f25b7dd3f32ee7ea3e8c318595f40d48d78a52df0532e259146e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha96dd5f4570705b3f645ab477190907511c2793ea4b411d582aaa19f57aa141ccc91fd8e5ebe705534c65e956120a17cd65bd93bb4ca10ba31d587455f64aff85127bb5021b760d01afe185ddc48aeebe2ef31ccf1ef6a06d392c247535d0fb85b6775130cb23df4726c3ae31d9827982;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc94da8087fdabfb27434ee522109bf3b80f05180fc7ce574505d94e2efda1cb50ab4c73a7699ff40d0d7ceb65d14ea2a2d7432891af85c9fcf4ad617f50dae822f7643adfdd0d4b40f4b4eeec568005ae0cf7d66537354b3d9ae801da782a2195749a41c68ea9a74a48c36b0700127d4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd136d70973e1c23c4955f0d0e67888c792e9631e307fc23f88750d5b88fbe5cad6ac056e2837f66bcea899c2c015289a5a0a057a256893219767b5941d24281ee675f2cf24759b9b3c9b6c319ed479f6e5c0b0f5b471d816c254003cfd0de59c1bd93bac2b59cf87fd21fade936a4221b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3b2f94dcdeb56e460d04f0b756583cf23b8fd3ff9a003b48ff51ea40c3e0d948ee604590bf022e19bfe2a3861bc6d4a48749ace2bac3d7c882180c33d48ae66f29799ab0fc913beb2df86051b4232621eff032fffd7d175e09880372141a235f25bd6e69633b8a3fb95985c8cb94d9b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec3fa46fe743cb66bd701cb1a61720b5361c4a73077589dd3ce053217d18f469e12379df2d82322f9cb674a7cf7fbe5c77f5eeea70fcdb2371bc694e29992f2408cc188205e55b477cfc8c28d21ab1818ad7a65590f26fae5e97c694fbf7e4fcd0e131992e906ed2d51a00ac7b51e7fd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e53fca008e074c944f56b0972be8da0d3d38ea8e3bdfb9cdaa872687171d0aff6e2530a72592b9929810e6804069918e1507ac9a706c7eb87822eaeb450e5be685517443bdf27d0010e9ae6ece9ed1b2ddb0db777cca98eefb90e15e1dab75d54999b47c9cd797700a70334667177700;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2227048da70b37d37833ca3d2bf26a9fc1d2ee668b25d32f1b9cb327b5dfee3386c2dc6360fdc7e74c8a15c2ff8d7e1d746fdd7a9f586a5da0c8a503e3439583b42777904e4ed7833e3bb29d418150e73ca43a4252c7c2dda70e131cbecdfec29752363069b7c456b2d5f396972b255fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h919382a6dcd29b8ef712f171be579a22b1863a3eec7cf5ab7feead6188679827bdb4870a633d80ccb89bd02b8aa6afeea448d6d1e72ce3593bfa164d164d91863e6a914b8bf4bd7dbfdb147f0ea90ae7ca885e5073b07c19d467ddae48b524c5fd16fc075c909a1bbd2c2e9b845bed432;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he18db58deb18b7ad33f6af75305e9d4057eda12e9d4de0656b5424ef3793ca1c8366438b97d678c769f31d5ea78cd5df70b4ea084b982f69a6e4676e05b8eeff5a3e223645c41ca310e26b679794b7221b7de7d4e645ea78c1f90b20202509e9afbd11025dd3c6d65c2d56bfa3b9c7497;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48306e6db02e120e47a9dc159766f82eef39500a73ddba99b913b23eff9918b72bcea14e70e6e62e920765d71c9f2914dd40e9bd31ed4fecdb00fe2a1324d3980f021b3d373a921aeea0e144795b134ab29f83afd1cd87396a45141c4ad3f4037223364b62f7936527345c1db20040d07;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h336085f0a04ce81df00920e8f0dc089798068a7309fb3b450ebf799e9478f28c39b057cdd69275da83de8964b1549cfd72695b11b16b3945e862b6165919515d16d24c9253f6fb712cb78beee875e51072d00c6797a11dac6d5c00ae693ea3de4fab510e084a4d3c04be189d8104270b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd54c2255436318677f9fb09bd4a9f03df830411da26b882ae16dfed68c416fb4258384aac475fdb3460d319a5fe5e8d3f408d6bd15119356f14d85b94ed898239af6ecaab260c46e8256757f1e709a7298388a21082eca4234b5af6eebaf7c35404975c5572e69ffbc9f31909c22e15f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfbc702459ddb1b5f0767ec237c59b74dd698b251db6f72546ae1b33d0a5a59615c1b8891d32ef55ca578a6e2710863f28483e9664b913d1f508007cfd4f867180968a58c1492360a767b175b3b836b14782724e9d6dee59f1179e9726cc5552f213bb168c40151cd3eb0837a63a72350;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb68cefb579cb071e5868b1c913bf25c60b4c76be50993811dbdb8a69982fe4fe7f13cf68ef452da1f148deb4151fe4089e95e0c2e802b354bd9b96d6bbd7f5b13ea2600aacd3e930a60ab116850ececb9a3e67fb3f3e61f1715512eab9ef02e8a78f3215920646ae069d0d8baab4d8b26;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb504f92f8ecc3128b898236e684ee70f5d4ec5a2573990ba0cf66b4789520b62e1ccdca46072a3a5aecb0ad08bd6adc1d7e1a57a75ca687f239f141dd8b80192629433a1dee4eedf6b2ecfd3ddf38c0cb6cdeccd635f6ba6fc07dd8b9b0fdabddd4044bafd94f0c6d49a0eb2fa774b377;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h792e408fe8ba1a71a71cba17134e6a4bb3485ec231ee78d94bd53388712331ba5d4b22d319bd90efc1fa812e01159ec1723c8c749c55d857d11816c9a31df16fd97e86759834e67667d308d4ae3ce786f2e8722574ff212b6829b0cd427361a4229085117c554f2baeb9ed11aec497df3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba37f1aa1d7c81661af7c8d79735ca1649f5da20365bc32b28865c4ac5e6d5a8a0f29d18778a8925ce284e2e18f6bbb3a540976fddd12c500ab8d6542b7aa9dee8528f2d76cc93aa5f17949f25e584987d42b88ba224ef64e1ebe97b9596d62f0a084416817f196ef7619661a66a7ad47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5157724babf670ea431db1415e654eac45007e6ab95b3fc371907deafb0636313c1e8978e47a730704957863b0c357470219e922f6b8a23e64a971ee32d76a3a894628f84149449e52dbafe06d515d59f4afccddbd56bcc0f77ec9665efca0107d1c1ee2bb96d7c1152e000dbfb3c4537;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7abe5f7d11e9720290a58181b6aafc8cd4c3a540f17c01541c11446f4ca134afbc0bf582f48b6559231d9c3cdd74a42f67320e164248755dc6a8123ddaa7c4c8dfff833654970b1809c5fb33372bbafe810daf09fcc532aadedb7fd267fcf39d5cb3575f377515d2b58619f39f9a0a958;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h329cd0f12a75c06d67cefc008f75a973f436d25125549da727ee754f7eff363b7b6b5fb318acfbc0d9725bb287058d89c7bc5659020771684cf2e21c780741559eb2675dfcddb3042298591ba50fb590b3433b421bf467f491ff7802443a1a8da8186f8ca3d86887fc75c875522543ce9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89f914459820e44a7568ca0e8f97a4379b33004e2a0faf5434b9010e605b55340d45673e6503d6aad3a4474c9d34a04765e3e9c39bc31e7c283fb3ca2f4dbe4f25935ae89940f4a58f56fa555e135c401866eb77b256b799f8dc6e9470211b6eacc34deec20631e1a305ce82891b6c592;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbda21dc36c1ef1fe646560a3c96ca8912e10d9c4245318d11146b762803bab6ba11e43a41a4a985ec33602d7c7b1805519881d57e81c806926034114d159c74a4a8e276d14ac0c3c77e0615347881f49a795c029287371a8f78db825393754da526e63fc5bc5710b2062f9e3d311f4ad2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56d9d01cf7b20dac4f93a80240eebf0f6d04ff1aea0c814914e9a8e7fdb012732e8aec0e330eb79b19c6c678fda15f37bb0d6e4ce1f79eabf67e417bf0fdccc119ae49163b45d469f778f9ec5f80b6b9aab24a92bbc2705227ec6aeb61882dd72f5f50227390cb279f2b10c8b80c79340;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf879bee2514d33d4779726ba5712530aa5f1e948255546c9aedb25d0ced89b6ec3603391b7bb894b3e2dcae555016645da6fea094bd071a1d8d0e12923f6f4ce76b5c062046ba8b4a54af294bcac687077715862628cee23343ec1854b7ff55bcabd0d5375f33951d986d64aa72eca061;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74357c7edb31f63c791ddecc6b128cdf71ec06451bb70f5bcb0d7b1ec7a5fab8a7be0f99a0b3c50da340186c4c56bd75dfed0bf316fa8fbc84507522a153911ba40dbb3f3f574f83ff1be37da69392c7ed2f2296f30a360631c74b430cfbd92b6cee66a835801d601dae94ba8282e94fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcedc177901e50ac58f6ac0666d144d3cbda0520a9a31ac94cb134d7ac3fa41dd4a542033a0b41a912922ba1db6fd7619bcda3051ed159858f3f339cb45a93ac4aa5d9a7380d1d151add9f1a12148a3e48db56f4eba85bd3621a070b21145917028997898d3890a6bd7d3640800bf2626;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab8d03e678a56dba6a492f2e35fce16f0c8bcb762006fb5b5b8ec0d2480d8f80a2f45f81dd0de485a591ff539c5f3914825f3cbeb86ac7f2fe8b4cdc3e3b2f1613d1b3fa97ece24627842149b5ce768b5e6a72aaeb4041878997a837ac4a366fe5c31c48554ad76d4cd6515f3217004;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ec60134f48790366ca5371dea937fd922d8057c55532cbcd55d18337d8f1f0bc9fc76431cd794c496767c440dd50dd3063a474d2a94544877f6458a626e00ac6ad8995c8096c04e72998981fdccec151cb2093ff3f4161285464fd04a181f7419c0cbfd03902cd9f3bd1bf5cb0405adf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h726ea740a2f30fecc0c88960202afa5ba9ca69f4dc67f028db96942b6aa77cbeeeb56bb6d69db1efb513115063707838f23eb5704230e8e8f388755dfedeef0e811b37ce600e1590c7803424791d59e8a742557d16d2dbeec9b7f2be8c6c0d8534a308d53a4e3c04f1066420415e3a760;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31545263d0c5425a5aea2719e0eee78cedba7a1aacd009b17a81b1fc39df9d9d8c8a96bb1cd3c6228df66f8d37ba41a37f7bf7d2e8f04575732327515af517171553b225219fc583c501631b9ffe9405a9cdaeb57dae5821e51f60b24bf68c48c7db4dcc3ca276c08cd3877c638d9df7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a2a4ebf07c9a0580ce98cc0c5cc78afd3788d1248822de31c2350c90ca46002f8975e1685d623e22e984e92cd0627557bbf5e05c0afaafa83a4dd7f3a723c224754ad9da757df76708e130282ce17787bd0f0114535dc4ae8d1d0177728ceef877b3eb6430cbb00a83399f2f1ba29527;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f6235d620b04651d0935395cda912b201d424292bb56db46865273c98c0776bdd203973d401fe7b957b0c8e161231c524fe28b1275aa9b4a5e785239bf13c5c7d5fa987d9b8ec5ec13cb4fcbc489ca3888f70eaa5b6169413c4f0c00f8c226a50df10d25f25a0f6fb239173a6b1299c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45ffe91da6ad49171ce0df932e658d69f513b7212415a97bda0404159852c0880bda7d2e5411eb98f17b9f41c8c495a5d0a17333415b016ff0710720caf039bae2f2c7c948ad23594c119cd15da67c5de1cb0c031b0db9ac64ddb8b8d0841babb3d822b4b31f9a1949eba51b63cd77e9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h107617d1fea47940f273ececabbd24e0b2c2c898dae01dfc227c70e623cbcf1238beedc240303e3b174aa32f053f8fa82b6b0b22020b0272f71fcf54355c2cdb8d0cc2f1d3e0ca17fa5d7e98b76bc170e21c627713a0173f8669e90d963bbe45a6dd698537e7c0b3f0cb0619369dd6ea6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ba56568d12202064d193bac5720183872f8a07f38cd243bc702b9bdbc8f9ea9a45f4856226f09c0a8b79835687503ba4415e9288ad99d5015bd7a7e68948a53365c4bd69f7f2a6d91f047906a6707586e13def57e86dede5023637d4473effd7e3c7f3eaca4df091a584b722a6456623;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e3f2425590b06a2c85ad86dd0ff13424200982503a42dbcd03ae06e5f70a220f3164de4fbc5a69dfd6072bf5607527e4fb4f6c30e00989a270a7eef310f8b58a7b2f5159dce03e9a89b850a4a5110419f08dc70c8bfe656ae14079fb329e6fbd91c1babfe4a1f0c3245b92a02b7d10d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f8da7cc7f1e736574ff83bf1d3d4c38020c867a6a8cbf3dd10d71aeb4aa315e8d32478f0a4ae02a2bba54b6423faf2eba9a5793aada4a8b40233a416e1220c93dfd4a21f18e354fb5df8829cf24871436d58d4bd5d0e57ef19ebb4efead37cd00463c01f919aca8deeab3ac28a594f53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd74a6d659ab5e7b6a8c8db4499896d6795016a7fc99c52c771143bbc25e55d2b448fa5caa0add64ec2d29810a9899cc7d9c3486d20419e86dd56505be070b1a24e80c31cb0acebd9daf070315a7ee7381367ebee65f936e659934f8d47c7f2e8c55d02c9e91a242ba6386390e4285d6e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e26576292688e140e2603feb8812d994bf1417e271fba4d9271cbc47da4c2321b7fe8ceabfb80fceef1a9428bd2af4a94647cf7b6a3e8ed5d0244bff9489700824f712b8f3309a7f51d7543df2bb7fe61ed43a9dd55c6aae4b8a4a872947a5765514465d2710745005f6bab16eaa362e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9944597d38297716a32b68ebc687ad4c31f2073381546b11272e798748e178913bcee4e925b6759863461d4ffeec6b7277e6fbfa842762636c546519c64ba87749dd170e5b2b46b9b27dfebe80c04291b69c9453892f37e6ec37bed69c8f7935acca5020f55d165d67095db976cd5b2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0d779429fa1a4083c9033ea40e6298323bba8cfdb126703945d831827f232211add7d6cfaebdf4ed8df9bdfe676df43526163a448508cc014ae614c8fc78bd3016b891966f302fd48a498cba308e43f685f132b56954dd12346cba30ba9ad204de371f648fc9b68a3c3440ecfa8fc5c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5bf84aac11cd49da7cfa465fa6e704af48fa3b4dc579b6962e2228252f70926563a7faf065df26fc989a5a9c10184c97c63bad5a78fc942d63de7988c8f5cdbab495e6027e1e511afeefeb29d04768dca48bd55c7f85cf17ade03ae577e4c7f6777993146750325536a9c2cf09aaebbb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4513f6d6a1b29bf6bcb4a75302738e991945417e8c0e2ba3be49f4b2451f84a9a85e484cab0eb4adc5a6a7efc6b5a64184db833f5655205ae717918f7a1287068e7d4fe9b5b6209135e54bb3d1e1d2bea98a3548dc37129cb011242a062f95601b2950d126b6face9fe72acbc7d8b3b05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10a2ca4f968c48af10804943da073a97dd7896f41f8ceff3468693b0a0a279f6a4be8234de9c9c54841da2a383c2f82518b3b6fe2443b065985d017044bc42402ae32826e7d5f1ab116de5752bf155a19d206214bb58e9ff5fea28e0bb08cae3b425b2bb4284e20e98c459a00f1f012a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2993054f7542692d4e047a3f4ccd34df14c5f8257ef427c139ff3e10e95672fdd39a5059ffae03f496fb6299c08869a917437eaa3c23122f2130bdf1a00a6ba9d519c5e7e67ee7466dbd970ad30b0ef6b450dca3405425d623f3b20b7e13bbf9ccb4ff301fe10632aa613b4ec2082195e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4567c9139f7361372726bf12cfaee0a6e5971689ad1be4e58ac6014b91de6c8c3b2e0ea5c4f00adaa31d908045f6ed3d42b2a971791440bc745976ac165794235a1939729acfc3e74796f4b2b557b3723fa2d8a8ea1d9faf4cf3bd9cbb7656f35e2f8e26d55cb8aafa8f8abec961c7d64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36e7e2b1096450b372a1d0a042d180c41da1a5353a8ed54ac65daffda9c0de9c127520cd7047172b2824d8d2b7d099fad276dc11c37a18300933a6ccd8218509b8036959b8e273f9d55e712bdc29468c859682b56b4cbbecc3b65440b4e2907f9eed8a85aaf27acef6a5a3c5b75bc8bdc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7a7cab5574d610de62d43ad621c4898716cffe7e40431181bb83b2cd55cf912c0035b23901060c333ee897c0ac3e49ea4090273ebaca6f7db487f9fbc1a33814019f712f1a553a882e5c86ce2a5970fbd16d166b30d2c4418f2352343ec0e28f7e79dae4ee49eca6771affdf92960d72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h380375d675d76f067d59b55a352396b1357c4782a4c9b69fa36f28d7c3ab29f6e0b9ba098f28ced542cf036fadf19e95b416ba04cc7cafb8c53bfeafcf6ba2a06f4487f43a39efecb3f8dc44248558963bd044547df150c82d42b44b150c008828f77340fd60c291cbfccc4a59e93018d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h238b3ea325aef6362a9bb4c876e4beb871e40bfd94f3fb33a8737861da514e39cf89d096588c16a38bd9bcc80e51835f4fcbd32626bd0c0e18c81c8041fa0bbee9caaf1533c7d54a19c2d80dbd7b0224300622ffb5712d2f0049274cf55a1e640ba6330e815ffde7a281b36ce36d5e75d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd22f9ab1a9548a1f1fb3a5e1598dc3efc91b0b96aa0d7352803bb2b2e5790c2c591d766ca593a5864337c634179832c771889b06279e6898d62b86255c7ed0a5073ee0bb81056b63ed079052139c684a0952a3f460226f9c39e9aead961a8940a827f08ee34a8b790db81d741c30002;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha11f91242dc9ee5c4051ff744c769f8f8a9bb9b229c8bd3e2d4d3835b0b6c7efe605b852dcb3b657f082df2fe5abc6e351dc78ce8430b35ba49e5d97232d1d7fcc6c8d8a8b29827611d30dbfdaf7344d04daa9fd762977f177b6773f9f9e104dfd6a83ca837afa908f066d45fc55ddfbf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cae7bcd35808475a7687dfb7b75b7ef6bcd4295bb5880e6742d07a359b2f1a66aa80b822798572e5f75cfdfec0f8cb1196b631e14d924366137b2fb300ad075e24fd63d40a7734d3c7cf0e68a5703c231d0ba5615b84c6808f94c233e4f76fbcb0fb18007623bae64418c654cd66d73a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4addeae1463bfa4129409f1619a90976653bf2f6976ca3c5e63859e91adbca19fcbbb558f1a4fbeef2f8be6665ff09a1175535f26179b755f5da270a4df7d554e6cbb33b1b6f3b6dc75d65b4687fee758cfa35ca77afeacad0e82a8660b359b1d26d8dce1debfbec18b5e5439529f527a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e7f0b826a83f033bbf996ba61d7569d638faf32f10c908a9f5f240b3fe9a6027c4f0e80ff5d1c934c6641048b99d64bccfef225f9acdb8252bef57cec43c84ad75bb9798fba0cb4537354f312dacb52163413d2cdc6f9706c3c7714048b63cbf79a9d2620d1a0c7e817c7f056b2b6365;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c0319bc4838deb6f3878a730dc2396abbd1ccb25187cbd7ae589f2f5135ab2329527c4ae1e3a0a063ad93a09e5e0e44381eb6a36553f54e1503010149190fb6e6d04c4c8b8f094e19128d732593d855da6c613ceb20d28a979fb74ef7227a5b89f0d65dfccfae7efa4eb2e71c5239e7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfa0b21be50e47e5c3292c106e5990852b44830c9c417c5086e9e09973f0fc730a50ba480e0267cee9eb8d16bdb3423a9e1b58d69504e2fcc8fee7a7ab6d5b425cb3b03db4b42a25fa8fae418cc362e251b82d2233f159022f20f8f4b1eab1932fe3d497b347e22de6c719ba95adfc89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h967fed136ad84ec5ec22585d196200264e51fbf1f9197b4703308efb9a3b948f2e3d3cd96866879ac6abf0bb557ff199c61a745f6642139f053c8dffcc1e4b62ec71373ff8d3e2f2fd3de9e2d98ee1a5def65499393a95be5335149a0f6af21ea5a8342fbb394085a17a8f43fdb0f53e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe41da48e23c33f31bba27b9167ef3bd7846923c14e48c3772112692110c8cc4143de6ecb35623e5fba1e49689c7c2903622cc70fc1c37d210c481b418725ccd6c65b10d74981834510872dbd2257320a8a352da49ed7f7153bec2cb7d04414acd6f55ba0b7e667907faa6640ca22869a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ce1a683521fa230111f9f447e97d2d0f610509181e743c6ebfcb05b435a948271fc2524ea89539d7f23b7882a37f3d8e2cc39dffef69b420fdac5d41707c610cf61152960cf4c6777a1d6da8bee4e430e1e94ea7a783686ceecc2661810900d2de31e6f1e43e0ab2cbbc1c14c4bb4aba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf280fbcb78d63676e4ba1b0d6c063fceca5c003cbe90424a99a8d517b02ee3c75022db62dd4a169e83dde52b545e70e5fa451e8643c3c0b67a6843ffb48368e0dcc19b9844b24a83e948e604597441202d067ab1bd1b99edab0f1d3f08699a4af57ef2487c541c69e43dd77e25c0f6c7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h603a94b39bd5f7e212ba1cba2cb40648bc3b33eb257e4349b308d7e9fd2b9125842dde5ef3709e2e31a201fc539fd0d9a18297160eeafa9641897a912a474a72d8e7608a8f7ef7bb6c8401d6ab7346691f77bb7e1223d13813bfa78223815323c8b1d7fad52b513cd2034ba73a6d0a41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8a12eecff5d9b722439f13ca70dcd3a039a8bad32d7fd4421bdf0524c86cce464af2287e43ec55b43ea0887548efa3ea36ea07874678653539f8628e663da6ce5097efff7404cc15c80b4258427a8767761b3fa7279fcdc3a583b22ac10d1b99e293dcc222ff9fb1ea3920bbada6263f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdd6a5b6a23255dcfe6808fca29e623e50d1ee9beef67570dced03e49545ca7a83d3eb70f86ee7f5abf77b806d2378a48b83224a3e97472c6f08f325e34f61859a7d39652bde657f0b91b3adb0157931165db703f76a3acf255a453a924ba05be98aafa5251c98c9359a2ac812823273c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9d80cfa271e204768cb8a06029d62e0f25b453ff642acfdc585a07221949b09dbd93f619e78e237987f71cbc1b0846fb7140a114bceab86fb7191e381e93417bed662a134e66891886ece57b474f6e26729a44a9a6c183bf745ddf8668fc4d77bc5568a25689ac4c07962ef420382156;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd710a65d546a14486d010a9aaf9969b6ebf04306aa2c2902243d2500be4185711c25ca2160a958639696b532f300ec972333577821b467f289b65363308aa9993b46f44e6807d525b2cc3b0130718ac127a3ec6170e435982a457ae004792de43ce056f4a1a6f38129703a552eb1e3c33;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd02d0107c44c67a69a12e8a797f7686f79ed7580c47c14e2340f34f81c7ba3f2ddaef4b78e069cc755e12a7edde4e0c1f059835311cee545892f0fbd4af7519e2f0f2063f586501a13da5dfe37b797a12346ce9c48edfe953f6da274d945198bab8f0dbbc4b4d394c1ca261661fc2f516;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9cf6753a4b7205902979e84d154c4023ad1806ef650d25e843aa900b2a255eb8417b00ba53c358d6e5a7ac81a6e137bb32f20ab6dd0f7a4ff2fa8ea9cfc968458401650dfdb74b4a0978fb82578685b5a1f26017c1c50b2d9082cc2b2081a2c3e7d0781ec70563700ac02d5468da800d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47dffafb0a72f3c0e939479cfd66279c4e796e37d55c68ff0319165d7bdce2e93461367f428d21ddbf47dfe14acb6540a6014995965953d736cf918b1f362b2ddcc62e0ba4cdfd295238b051be1c8393669907c7d537bf5721a43d01ad36b33de11c08a0303fd8f9819da6a06a6539060;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e8628d049dc84bb2b0ca778412dffc4ff2b4e3eb0386c84c93ab229d3ba50155e57c4217f96d864c54fd8f43455fed6b1e54109c34a88f0645d7342de44115b9b629df6918fcd8017aeb1c659099163bf341d4aa77c4d3f12d48d09c019f10efee187856e4822759e99cbe1f7f0fd53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he17db97129c00d380cb9a242a9c840bc42552e0c2f038181188b74005ebb5f193118db1ec8fd2cd47c29148674d601bb7a77f94a1f4b61bb2726dc6367e020b7f0fa2a0941d5a128361b9e349758ef22991c2b7125895e5de55514bcb0b05814cd2345a8ccf7bd2e02292ef898ced0062;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9e76eb8863a2bc77a66b69940b57175f2d8b1ef29dd6d885ccb22ae63a5a5a3d57d3dfce0a15cb3c21beb322eb0175346636195db3450013a266520fcf70d635a2025602c60b2acb3e933062fa7abe050f0406cd2452b6c9f4b84c8c7c4aec9697d6f15081f868eabdb710b32571323b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78ce5d1bab7b9cf719cca399250ca0bbd7bbf3a2494f0cc218c0be2df7c73ae9e46bd2960e93d3f8e9d8f49eaffe210a23eef8dd91031a2058f79824496a293539e1a43575a4fcc069a2665b6ac7480972679655d11f45ad547a49f602da8d52cb6f423893d60cc1b13fdf9b0100985f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c47b7bc295c6faea331c35be8ed2c9f429e6b9c9d1373f6537700fc483bf79fbf9336ca698b094ea848741616cc5cc807438e9d10d8d943ce78f9440ac707640c039c2625051490b59d44d9153d05500a50287ce6f84dd16b6b102f917ba82fd1c2c6bb6c6fe346c6849142157f21404;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72f12ffcd10a49725097cdfedae5543eb6628aa0868edf5c41d3beb9da09cc1a0eec188f0d706db0b4b3986d20c2785c7d990534fc37e11d63787e4106a3ce5238133623fcf0323374df5e44bf4d24e6b8d3f4d04443dff5e317908f95af5b885da4b9fc444fa2f9b444d77dbff3341cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef6922fb6905367e9b27d25507ee5cba802f02e8b3fa12068808846a7e5778bd851c8c01263453b09e766bf8b5de2e28108c4223a185fdcabb8cae2de8549d6052f458c580b9a376353239980a5ad7d08b0976067427ce8323f46e4dff2d1c4d96f0113c83d085c3fca7c6718f734c070;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a8b82668aa29b975b5caff69821d46e747ffb32a441de7db89da87a3a75ce60cb3828cf3930a2a1fe6caa462b0d80292cc0159389f22b6a5a718f9193567c086fa00021a062646c3b1eefcd3547c0415367365fa2145f8cc7008e93e0493da8a65217eb345b8681e563baada360a05d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h999def59f0557b6791acf4150fdd09f574ee381151e4044206ec636f52ab634248bde50c16509099d49566ffa4fe5c3927ed89b31b6821961cc394b2731f7caaddeefb8df74ae4531adccc52e03e27a29e8b89a7ed962eb96b086413ab557ba2bb27da9d393909b1d2ed1b42563ea7431;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3dc3daed5669cb24a9db1ab1e6be013590ae35e2e1de80cea1e01fff1ebe7db3d46317ba23a5a1490d8ca68cbbfecded49f00e3e6ca85efd90d17cc17c55d4b3c0cb4495cc1cf3c33eec59303363a7d6cbd7f13e43e0b62fe89175843f03c437ba9b2e2aa3e9782bf62382d8b2a5a39b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h932bbdd2a7511d1fa331178847a514bb56a40e20c5f68673841f741749940623474bcbe94c38b94ab03ec41b41e218061abefe944e4e0fecb613fbf1046838d7fa8802301c54081b29c53adec63b67ac17947a221f86e2458778a5e0423f94eba9ae0fa7479e3178efe80ab79035fd2bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b08b67fe86fb0d135cac7895e02637e4092f8876783c5b7577e60335d60d5f6b8dfaebb7928bad2152315f1488a43af4d96b56ff4453a0be7cbc7d4563b6754f8a47833c0ae287af3dd4446374e109e5fab111f564cb9cbcf01c163bc5697af5ce4b59012ad61b3bcd9ede4d12507297;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34106eb0ab96c4cccfc778b3550a746084789144bdb7b13810d2d3d33e0ef85f5eef832eefc3c92984c907bbc16f086f0e7ced734d32a8df8976781a69dc7816c20dd4a85dc376c9d1ec14b97a760b02658adf095e638e44d5ceff2fb4b0554609c612eded16913ec208c55c5c1faeee5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42522725a604e669e36825d2ddde1e88fd8e1cb298d43e36658ec074882ab50e9ec1108a922d45a2e23d8f5a2908be521f4960fb82e58acfab2f3bb43333688d5bc4299b2724b86f63ab56c31578a407a80c19efdb63bf7468919ce6b8ef88c1bc3ecf100bd4267f58785c8aeb8a01509;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb34006581e17676167131aebdfcef055a3a3f0b6eb83c1b9e12277c96ca94d07f6ef1b16b219eb2446aaba809d338122848bc321d59ac5dfde9275e4223bf66aafee54457869471b51cddc00d22d7ef98870f0731c3ff577d6c746eedcbb404644fe564a492415c809e3a4a7dd18862cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80073a56d38a40134cdcff632838f0ed095449a73fc47a3ad9e1f65bd967582f9dc3e598c5700cbb3f01f2b2f8200c1aaf0fd414011a39e7b3010a4dd19be7f7ebf0466b40e860cd28da9014fd0aec8e531e0f61047e1f64d670908c0fe8d0d60351fc85da1503353220da464b67bdcb6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f1789e68d15cb9b71afd12fdca8aec5404abaf4d56357f6845f950f1a1f5ec7921bb355571cd2784ab6221a845e3c2c30b7c73999f6aac6882faf63ed7ffc6d9068bdab7d5223b344dcbee00bafc24b857829d5515221018ebe185a2d93b68db400afe64207ac6a75f64073d7e5108ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he910c332aec34d7187f7a8218e9ab3bebc1e4a1cdeb01dcf6b20ec5e2640eb384a4c5709119dfd4231811de6dc8f56b5275be5c018deeb59bd72fbdc20b070bffa69a826aa35664a6a77cd8a05661fe5507833750005e92b40dcc1fa55a50362675e447a16eb32f1c67ad4818e4259d78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha05a394361517b82c56a5462866df82933c822c52ade0e661facdc0526be5ea9746eddf4d02295726f4925e6752161b0d7fa34af02e02792a078167afdf53a4e8fef0c422b6f8c26d08af13249b8605bac6bbabe902d541d1df020b2d342523845d96d7734e83c91820ea47400d9b3b00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha381c7435270d10124cb09d7a2d4fe1c9ee94cbd4503c985608dc4902a52a2625a002547ecb95ceb1a1cff2205b46821ee81306e83b3946e8330f5ca9e536ba709f9354694674922f41e0d688f5f222063055c4cd42401030c7433f9c9dd05a6617dfb0f1f287b92f69a2e3e3e14265db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ee153ca03ea3d94bc905a1cd41b005b9c216b3a630568f7b0f988b9f625016b07ac1d0e1c92dce8d9f62b5e18351a0d4042ef56d67661e2956411188456742dc738c387dc373d95653e9ce0d3a014cd170b3ec87cbd7d14ad93ae59d59426afccbd7774cfb5e70e3e7dcb282cf9e70e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d73e5494a76156fda134b9fb86fe227fe9f7c929ad64af4549528e1fbb35679a2c7f28bf77632f1f5faf5c5637424efe287fb44437279788e5c3afef96999c660ee6f697f2f4ae7e25467eeeb69d15126a4c896db6dbdd2fc6b4fdd5524eecbdd5fd7d09218af66ed5c287319f4a19fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1cc5947ff20aecd962a47598bd2dbaaf7aa5b741dd4858e236f964b223f729d401a139a970e58b24c40f63d77d4529ae51da36a7890f7cdf2ea4aaed147af4043416daf71c398dbe97cf99a660911a3a8b25884fc8b3e6346df1a413c371cc39bc26a2a1ba879aa798e04956f7418a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4678acdf324104de9f3bc24d3933d9ec6f31e5bbf4b3b26db45d5448e0e617562fa2e3ec2b256ef78719585244eadb2e01bd512300300b6b46c3365ac713cbec67fb0fa0804e0cc29cdb92c4ca51f65ab439fcc0112a3aecfddeadb396f0a2bdf413bd04e90067d8fb10699f6a35fc3f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44c9949df26d97a762ea87ff82fff9fbc89029323d7d6cb8afa5fe6eabc24b15710d67eba46fea669d5f0940e9668cacb61cc26a370cb06be1a0a3170e58bfac42fda47dc68788b806a14c09c310b160d5e98e991dca523e2ff5f22391ae0f224d8b823f926150508d71623a253ce9bb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h847f4173224690122f12dc4ef6d108c7530c93dab123903d621c18e91da7fe01e6981b0ff58b81bf6671985131106731b9d60e2e7c32923a529a075db20c531dccfe6058145260aed60fba2f71476711b27cc3b616850dca5e1d465e46d97165b5dd2fd1555f109b734419cc4b1d36eff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3058e3a156f39dff8f8f5926e4451e73b1e214ce1ddddd1827decefee26823e263d342ecfb61f44efcee1728f92f605e0dcabf1287feb519dfc00553b2028674b4a4acab42e36bdb215de22f41745c7271abfb22da325a6def6d39bc1171b34868a8574e05d94319f5a93249a9aefa8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9dd285a6cc48c5fcc9299af910cd6ebe55684fab8ca1ea97138da2fefd2c6475e04f173345d30f99525489b4a18b9eadf71b3706c303c699ba7afdd3a2eeb3c0552713886c11e9f18825dc8df62fa4064a2042c39ecaadd9239c0f55f2fc409f6f701413f8192e5f2d3dfaaf4cea711c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87267e2b06db44b9e5d516da9da7b894a1618849f92329c72fdb029e1c4083ec142a553e733212ba00a07cdcab37793180bf5922deb6ebb9b79aba358901de9338c54bcfc9bd8f606bde1abb02fe7263cdb5b1f7b0db77a90e64483eae0aa358cd82e8596e97c8a79d13a11882f418b7b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha79316f4a6c53cd798586b254c72698db793ffbfc9f88945ff0bd8ac41a0aee071c2324ae5b70d0765349a7f4181e3d8eb7b3dc5e7a993ca8a26267f9377b1ac756f024563395912c9606906a191a6f6a0f2cbe6f4914d6b36e4d1885357b2a040f16dc51e6940b74fcca719670de5bbb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29754911edddc469cda90589c338d580cd1870b135abf9b86835f6bea5911313f421bbde90cbf43909939b3e34a7b4216a7fd3f898b2bcad4a16d0a76e840e912de5a089be6bcae518b404ab2c0dea43f3084bb24c5b018220ffe6d0aa53b08ea7312e7236c71a24f996ad0a499be05c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6e236f768484717b71fe51c767cad75e7330e000521924f7fb1b031b1b369782ed32a0bb10cf4d6fd7e40bf7920c8a169733831b989d5c13312095496fc76e1d8fa08d2f312f7a7f9176f713e13b255c221b720d1063516ed95a8998ffe2fd1717c9d144cf0167462e742513983080df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc38fbcc4ebe80eb20d60c5945564cfe9ff18681109d1f195c7d3f74853589ae0577f4630bf132a95c468fc41f8fdf7420f652a73702aa1ca7b9e63c55c0819f5c8c9fabaa8a0b6cd0a0c78852236d16a006d522a63961ea47139457ab6d29abc2731310eb2f23039d2c91c902707a5291;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1d7b6227ce163848d69ad74206cac229b10925bf0a52e82c10b55a4ca48a7414fccd315ea17240a56418d9188b2e814a2d47c121b8e6e21cb942d85e79c79e621bcd3e8b72325ada264d5002491fff710696a1a12eec6340394ef9f6b2ddb4af7fbfefe1eca07a6af3ed36a7636a143a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71e9de77f42e19d558e16e4c588a5e38eb65638065c826a7df761098f08f98ac147c48b871a7a79bc787adb943a03354ba49e241e3761e3315534d071b375c5a9ad9470e3c955048047483ac8891448b0e590635401c4ecf461adfd3fa2160b24e9c3117ad202befd5eed4b1974f5da70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc02a5c4fb1cc2990129d7a28f3c73c478557b400fcf99899c30cf68bfa3377b751e881703b0c4d8bf769b1ce38b599f147c5179b7978271ba293c22866083e8f020f6444927f9e4a1b79bf30cc1c7715b0840025a01a6e7fc3df3d19e35308fa54b3af0e887566d2426a0651c37a2d420;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fa652e3d0af3c76ee012d8cc1c003b7b62cf92f3cf27ee9f4b3500bdabcc9c6ff429b92aa74ae14ff210489d32e400bb3a3ad6f02d02a01343bd1d07f68d1fa158322e1eaeeb2a1a565e46794dbb25ecc973b702963cbfc9104048b22d81475b5ed523733dd38f074ffb6a56d3130976;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cdc31760d417d16e32ea2a34e83730ea6d9f182b4c7038a1b2d08aac503296c7a005ef46d308e3b7e892570dacb72d57ba571ef5c581d49665254f959a5513ebe94d9650a81c19d86a35dbbc69cafbd914795ee8b7e42cf513eaffc4246fd0fe3fd7d905798db2b0ef8e9993fe4bb531;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d7638599542b747f53d512659abfc30a553f2a6a4a7f30c08cdfe89a944f5b4aa2a525b45e2553caa466ba6b7a6ed8e8cbf01ce4c94a9392b054c3247b1d3a221f283aa91a8db2b11ce6f09f883d84e58d23f0c11dd292f781ca54fe53204a4d7fadb865ab6cc713adcb81cdb66822a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2acfaa664274b461911058a9626ddaa28a4364512620e9330128432a58c397bbb86168896d89a218d598e64e2f02ffccf12b7e471cf4b4973f1e9b659aac0ac9c98e5be7d48b05bdd8aa38d4c3c1c7b2302f9396f607c8e1bd72825e891ca10d8132d2a12f7313d058d82a50a90a47a61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb930f5bf46957e28efa189df7373f3a4bc1e0235d6fc61a2cc78fe9854bce3dc9a6ae0e53dbbf2c41fd2f7eaefe8d7241add8d9ac33d98174ee249f36d7619397a39ad595203cceb1d421b28dce3fbc197651b0189eb7785cb6d3a4757503b0859760e44b38c78b0799b9dcee4df2635;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc07c2f1eef545d558da6eba3b293f27c537c23ef6dbcb283e57af287e39eb5df9529c67309f71394e3c411f91ff62c3a338b9b2c781c740e0f39bf8530d79f96679e1860dde867d7d940c704990e77e3226aa6b43e0b043f8a3cdf48a39d24501d5d5c4c510b6c2a79f7e317b82c4f3f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf85b3d7a93479f0537e0672bc1ceb3488a6c3c65fc78a66e2b22d384302218e582ee5866121452b5b4bfc76a18e42090bc8adce421e7b89fc4bc6cc0d5637b5abef8021447d9b0e312f7b196aa24c3f38d9f00dbed75008b23d958ea6329e228d9d31574914d448d782c0e07010f0ad1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fc8156a9739762ff26aa987445441b6160e34060beb039cf0304ba0e5f01a7e46393a461177639398ad8d9fe6e28a8306f167a9ce9808037ec3eb68fbc3cf2362f99fb87c697b9312b10aaa3b70e47ac8d58d870d6a6773601fae4b1b16b6f866c6a031a971490a2a9a2f72d8069ed5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1d5a95f65ba5ad76f79bde3b78804acfed8f3fc966733c199ec65fa8825524f09a21945531d0720f45029039b0e217149d60a4f608d0e9e15b318eed1380747ccd89c71fae286b687b761bdfe14e43f5310eeb90b51cbf056b49d14b93a07b2b0284bf31fa1090301b4c1e755fcefbb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1d724ebaf87104de3257b1bef7500daae937d3f677685964cf71b3da97ad07b2263bcccc28a50b80f031996b35a9bdcc8dc4937daf54b5b9afb62952dd1b3e5b50682ab2813c5af174d770ad19a9e2381bb710179027546b2a0a72a2933d15ade61bbeaa3e3f740dc2d9ed8404e748b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf982ce169e045648ad993359a60ffc21c90ad2e378d8cca059993aef90081a789b139756cb4352e4ac840f035730957698f12211d65945dc137bb5ef6cb34bda019634f5fb3707e601670d6ba4709c307c594658925568cb7a9c55a9991fade43d445c2855d37f632d025c799d3e1ab73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ffaf5116f44a8a87c3a8137612cabedef04d1aa5c42565dc90609fee8de4842df8e836b2657b183243dc7e07dc19b7f1c5769a2316c8a5d31a7d96d4bf05c5ace553155891ad76920e8b10e6a8663cd922f29e6bc4746e9748a44302129df47b51e10906c2a5c9ca43d24a07702b9219;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4feff46678e31c98fd99926943722ac94f093d208d9e0ca503a6ef7620e7969a9195589222f0985b5ce68bdfc1cdb83d6219d0d9f4c565391c3032f261b2c711b13aa89d7b6ca93a83d5258331f0041094abd76c74f4774ea23885895e2123d96a76d09ba5e45d4e92b75e3b73186a920;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5146db9a818c7f538806ef0033582dec4608e2e012ed0af0eb1bd139fe33b112a165205f5819b7c6fb707be07dd6ea0bda7c646905cdc1fe4396382d48c3a273bca14144ac2d215956302a4518473f6833ce86845befe842f1ec703418ae38530de93b2f8c12cedb4991750a6117fd889;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c080ad60efbea00b29416f6f39bdc55e5013bf96c770c286d7330d12b64efdf31fa3fb17d4b823e2ed615d0b1a4b8dfd33ebd7d8e50a160f46131a16d8435ff5f1b61c573a07e559c153c98318b6854de3fc2207faa6f71ee6b110b46866e8b1a8d8e0816dbc12254093e32ee3b40d7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f77f4c3243c119227dcf52e4eef74ef7cd645152c168fae659f33bc5c995a612a8beae1852c94192ffc69be5a1157894d681933922134b8c17025e915fe4b8e958c4cbb15ac5b87fff2e2944c364630aa22a08e538603f0ec93953e49b3bda3aa41dda9668368c8f216ed4ba02246c5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d70b4e333633692a37e4b27ce6cd0b9de8abb21f1d37f76d9f56532fce4eaf9d9ed671f4988a6657cb8ac2bb7579bca7abf01fb3af1db00022334311ad1b3d34d65d6921652c23ad26dc78626e0a63d7a6c5e44657f6c69ca2959f7f56e774122006dbb81eed8e2d87da8170e80b55fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e498ec77c706a59f1e1dce5ff3f8b160a177bb1d4ac483064669be6dc4ef708b500669de750b623e20c7f76b835fee335d34d8cfca638c4dc748c303198673f52a6b9b65f91ac4c8af34bb1460f7e93c2b46af9be420e06fb67d62c79fcbb41062e3059cdaf397384bf0e7c18a97ca3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1df4b1aa4ccc48bf201285ad678a945040b044a2a47a4e11e3a9a205d2e211fbe6b45ce175151dc37b834df79fdec68983cd76bd804a3e3bae28465e0572b9013bf9711f080966e9a14b74f3defe5d884f6737434f49a79483d6470852ff3173836fbac5643741d1648b7c32f32a9fca5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2febe645ab6fb7e964f8b1affd8c93fa1a794c0efd4be0f23278f024ae1ef61de1a7cdc99a6efe2c499d88b92cb639a1be6ca0f8235e76001f02d4c40a2bfaa756ad5393e33f6c1255b3349208a8ad19c79e7d21f406257d1e1a40ff869d7a6b147ef36088cb29034eadac6f5ce7806f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9105cc4fdf6ff75df6786d1e06795f921dcc9cf9063205c9d91b5c464c0022fb4e5ee9ad7fab6a4e985463057374168a8c85f51572b586ff40145af53833a6c66bb6e894b9481d186417a0e88be9e609e05e2486ef5935273313cfa92494a9ffc9b7641c5d0b49c397c47f9d61a05c9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h890e4c1b9c897532f81c2f84bc302f31f9442b1dc523ce3c3695a8bf64cb7dc9dc148b641b5ae899a5e89b3778be69223d83be3d6d927835442c54691e0c062a1f70d57bb94a155f1f414ca0766c5fbdb668c098ddf40a3e8b3f6469496db9d22a9b8a06ab56900d58750d1d29f562ae9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f0a9b63e0f426d2def85735e54c681034090739b194d4416b4a49a342c90fe6bff0833944b27aa97178557768484abe43e56ef3556c291bfadaeb0cd193b8b8036649716b91475a2fbaeb8d9d384b7d955748375570f5e6f350cf055313200788c63c0f45b3c4935cd46344df126158c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffb8307748d75f3cb33bad2b330e7b98ce6ca426f078696744c9fe1af9c05e3b5fe00e6f69887ce18247f59e3e42d8c582972d64afb94e1f2cbfb8473d7e25a5f04daa169243dd3336bdb841c824c56a59bd88ba1e2929416d51db7c6c2ce7e8f7af1ee202f297679ed9ca156f8caeaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e87833c5887450c45097c525fc9ee1fb38e7aa23af7e999fe902e1ac26a864648890adb7919f82c78fb9dd9cca9c431abb4d50916e6aef0b4a02e8f62455d5f436d5383f4ba668c54af54d111b99fd8492072bc526dd5101db3675f4423260d3ee320e4741f07a2a326310b7fc48fe92;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10ebaca8b3c7ab1194d513d6df5e1e8e433c82f348aab7692043ec52c41d236bf9ce8f2b14a0fc58fd281a62f78c709b7e91b5f729f69180a3b25be8e0bcfdaf45e278a1c66ac296aaef39ab1c89604180b6b40279bb9bfd7f4e4501662b7609b638c13ad382008dbce15a3a43ab5ec16;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f880a548190b1b1ad8be9bfa5fc2fe7ebf4667fe2b7a180a549eacb624fe54f366ee7e2561a5caa759b793ba71441a8ee24dda02b5c5f16bdd272a2cfffca44216d732e5d26a0c8ac0f4b36abbdefe0f26de286834f3c3db720f123adb7593e556e7704a00480219ab7fc58f4f40fcc8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77542b09aa896225ba1b320ff3c7ce4a862572d8aec67b87ebbdb7a6254a7af7be60cd17f6cb1e6baca95cf284819ab0b2e6bc3d0a5423c494028cc0ff0b02282512c9cb1249f940a8885b1d67933e1cd81cedadb743601334398259d05de0affb8a9eebe2c283ef2bd920a94a781ee89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea441150134948da7a586ce0c8b29ac772ade4ab4569f8c33fa039a4b2b2c0c8c369daa8ac74d0229598fed7e30be207a76e042f33f41257e488f317c66d37bd9db52cc5e3f6e1afbb6ba8801e06e83528b4236843241fd1393c09654f36a4207f3bb6e63db3026ab10f88aa31e2d680c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecf0b99933e36bb3222e9c884d57f5364bff96e6ff99eef009915be3ecb61793d197ef6e02acb68f103a21ffbc8b55b1f9b66dbd4dc200ebe661bbdcf2d4b578f2da9bb66eb6ae2d700bc0c1c2c4dfe95f62944d52d4c0382c951fe664cfeb82349c1946f8a86534726f03407b8cc9a10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha382b1cb9d0fccb3733dfa00d1c47d9bc3c4309fc4d44ace4fbd67759c1f15404600ec55635778ecaa73f938d3d343746fa36222f380578e9a39f03218e54336b3c96ec0930406cec12f656d0afb35a43519048aa3c00501e0d29bf6f8357f802c7bed434b4b7f3b2926e1594638a003;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6333a795ceff4d77fb388e3181b112297d76ece66e1708efe7cb4d8aac2570472a55a93aed367158ad9bb57a8d538f30d5b9d11ef192e09f15fd489f2095bfba33b02fef1643989ee1ca27b0c9375b9479c4fd98cff81ac6cffb3f7b6131476aefa885f623fb3c05e8719dd256014af3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86dd4c981c4d16106600dfd72418c21438ee4757e41b8e403061e264a47907f7243830e12bbf1a8dfb7ebdf4aa27a0671247c5afc41b5fb1d7ceed52e32d1a9adcd32f4500951e88572e26ea40c04e6684eeb6e2c1b5f51cec3064cecea25c843503dc26c37779fc3ed8110252378e07d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9073924a97ef1e72ada55362e628f4533b9fcdf400743377f101557881bfbd72a406247cd97b50d3b467fcb0356f7ae55d715105d9ed2ffd892426076444710471e782de3eb9d659e7a91fe2a6e8038c568f49ead7b1fcf3cc87ba66cc381d37bdf46dbd9c87ff7b820c44f834a226734;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdde847232c9fd4aaa9f6897be2e7a1ddaf983c3312a6c9e2c990a5befb911045d4ba2b540e04de62eb164df540b4d2534f2a69d29b0af4115319a00e0afd6f638fde6a3033fc9128976c4ef6b9abc810c407e49c3d26f65d1f2725bbd315483fe66134890a7f83e801a01233621b9d904;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cf9bd86c6a8be5eb3a63b1587de23d71214a95c15cd7b49f67bafa0f1061990e941e3c09ddbd7f2a4aa080872a9e0744f469b7ec483b575b5b5b1d44de5f4312c626ddf493b75f33de36abe7d2e1d6a08af44b2ab7fa3648ff8f712d50feaef9899ea31b92f076a8db572432fb18aecc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9e0855fba87f8c7fc4f3254b76f4d708b17b1a9953a0fdf0202121486048ea45c53b36c600a3c403c974e19def6a743cb0b381483361268b371a6a8bfe0ebf4f6ae8b75de23fb3c0f1d94ce3b95ffdd856834b1f8fb232fcbf8c1e76d257c8cb82d8adcc49d0f4b7010c37db1ea68070;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h574f4eb3d906ba9c6ff6cf8aad337f8ad2f81d97c29f5a8f15fce442ad9938787a6048034c0a7be4881419e18e5b93e08b4e531314baf0cd914c1ecdfe733e74d8146069d85c1cf40c56a3d37944d5b6facdf83c2b3553a56fa734513e0a11fa87bd41395ee4f12679b1a020a82ab8bb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69fdc078ab450dcf7fab71953c05a278daf9d3951fdffa5add95fb36810c5b7c0b59b1a3cdb128c041dc80059dbd6dae18e15f60181cf3061989130e69f4f36911ad0a5c984b2aa5466a8c809dfd08bb550ccb811b97ffb735b033bef313a014ebb73f7dedea6c4af397211e63d27612f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c1d90c301aafa72952eeb8fb900318c33120b3ade51ab3920fc46ff2dd144e7a3705b7269e793b77efc47aeffb77f3272c3bbb579ec10372265e918369903a880c79800e8d1bdbe2d708278a3eec97b9f7cc054c65a03bc5f21dab28c5d0089fa2406054624d2ce34385bc37a643eca0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd1bbebc71b5c0a42005f78baf0e4595cb397fdfcb4bb9610bd0b17cea4371edb6184e563b4452f29ce624f85836a31df69dbfb9a7685582a6a7279ef5ff74c0f7fe1935b717e550f505c9e888d917b5552e29ea7e73f80a0eddcad9790f70a86697f1dec52e24ad413ec758e6fe68416;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96f0392e48710fe2483102b585a1b8393ce3f4519c5ec7cd530aa89a300165e99524877671da9a53a5390caed7a512b7e34cad4b928335fd7501b6e1da981222ffbd2d63d74a802ea27f3b748cac44154b76218a7608172bc82fa9e71572910879ff5e36f213513f2e6b901045571009c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h756a26f1d3bb6469dee86c57fbe94a0028119994a4523b87b6a0446093404cacbf5aba23ebb4617ba960632d6f121cd3d89118871f6a2092807e842dbefef2ab9f3697f0c61d457365cbc67b1d2335f0e534d0e262e9c7c0df0de4962e5946a0dec505309eb32ea59e334a9d31c6b58b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5346c0c66e0c1ad725700cce78dc1f4dc88491cc5f06354608cce6ce63fc3616b2bc800315c27e0da34cb502e142cf68ba2df95b9759468dec735829b608335c0b2e72be48013129d1e99f105c11b16ae75b4005bc8d3f059c1ce45d8c2ecba9eed3eb128eeffdd5b3cc4a3bec5236cd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbca03e3b1f2e093c1a050503932fc7c31d74f92d83e756d8fe83a50d31104c8d172a27a3d3d036b5416aac890d67a7348053979c1d1a74bfcd24a7dcb51e7ac8900e95b8ddce9913f7471540ed27fad6a5976218e90e49e7372837f4aa14c2ef268e45aaa4686a802379b16a604ad24be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h110c3e76149453648c3a45afe8c5c11e3317110f7eaef2430015584ee6f2ab4e743553142bfaee952c24a0c071b7b9553e7b533044667172e9073cdfc39885a159351ddf3b8caeae839d3bd6766a59613c877b424439bdec8474554613dbc6f00fdbd67e905d11434a74f84f08ee18077;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32944fcca5f1cfbc90c8e169a770d1fdd536fa49777d0b495fc1d91ecc7858f6f6a37197f1c04c83dab8e7af3c3584c1c1ecb1cd4eea410d927c11f3f5baeaeebc898aee693c06900dd10adf4597ce6acc36daa46a77b63c86636b701472541e0415274a605f92cc77ed96a507ca6446f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e9cf1527cae1bbda4251f160cdde6ee7399438fa8b005c08315d04908a8c5a301228adbe1148966f489915aafd62ab616649444ddbcf0170f9a0d413f90697e76b002215e2413556735364091f114ceb83e38091280c022d8c464ced567a0c6e14bd2708c77ec1c8b7814b72e9400b80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa551e8fce673787ef85f5d411453313a98f4d8c083abfef7004051a9f1875406d55333b2ed9ec7795e7af1ed90f40dc17b790d3148caf20e3479dac73c33909218af266d0b00496cd5040ff90861d7f4242bb57495b2c135815a5f0dd8af799a923f7b7746188d380dd67f57cfa340b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebc116b96cce92017dfe118d5c2a8dc6bc1647c9042dbb84b960f4918854c3303fe4d71cf0154c48e72e669f2e6c2d96e4f35716f70f68ac51147395b336474f9891b27752f7a7c1bc3f3b004ec536a3499839168ff1e1343e070748d68915744603592f22dbe4fae46060c8abca315a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0279d84c0477d317e37f1cdaed73501635728f5e68b0f1dbbf7da3b095af67c3d71bf01050fa82ff5326e3f6d7d941c4231d0359e3b6e4d0bc662fa55fb9655be0c67e0a7ddc8600e9ef288a567e2f9e84296e52ca335100b8e66e30b748c002af3782175f11b131135c6b6d2f6d0507;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h421ecb2093315b947c25249bfe176641d7c5a0f9dbaaab924235b00afd7b0291443a49faced3c9286baffcc7eb6f1ff7a39ee94c902e517d01bcc1c3b3d15ff60b8b4965a63e797abd23609e499ede6428d36a0400885f5d3774f8c7a41715f21b871b74a3897006237f40e2d20d31125;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde27683775fe55209daf2340a2a2644b96ef341ca41350b214a9e23933e2ed0097ef039354904e4ab1dcf086916de31555b3587433ef30762ab37c06cb26efde178a914d5affecd0c8a2b3b0e3860ec82e6c4a5c63d29aaf0f18d5d78c54379527d7ae802f43e6a5830efd13c8ede730e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he463a70b61e2684304103aae3b61f18c9fdb98ed13343bcd0d50e98e2588ddf889daf13599b7dc37d47900aa1cf711e3066fd8ac6869a51ea326fbe37222457ded7e0b63111fe396e2ae047b82bc5ab08500427b900d53a6467e51e71d6d5f49b55e19b7ffc01d02d305ce64c22f94b47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce9c81f835ce25f3d74b28478f6c8ae627230d19f33bb36416aeb9fc5f429ca51622053154ab6e77f38b7da23b4f98bd7d265714e38738b8eb69892a501fcf44c24af7fad981476ce8c777a3fcc09ec1a989ecc1328ec0e9588d57098e3e3ac9e31e9973d82475e02efbcecc4be7ae691;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf034d1c20686d216dc6ffd2741096ef762d45b1a283c9699af3bf7485bc6f46bb0d4d74255a6b4ac1f529277d5a6b5bad19774c1ce868284656ec25f3f30db602e34e038979f610b0945f7bfcbf25a5dea71ef34e5e162314b8c304ca33610b8859b183443cdbabe013b2abe9946afa14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37856b0f00a28976faabbb7b38b7f248bc1f996d767e808d507925b3a4df35189b7f0bf64085ace2344170b4825240ed9c67a467edb0aece9e3467e8013c5b7a145283d391f525d7943f21e52ce9b9a2b17e4951c368940b2a963e742e5d2321719f9714dca0a4edb7f55fecc4737e8aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4177361e8fd569338802cf72e0b407ab6424fefafe32f650f9c2acd5ff03c9099eef9f656ed6a326783d1b90ac817d4aaa4e6aab4e029a532c103c473b76836e7f0810a46a045056716aff4a786d0dab541d68e0b11f02788106690b405a27b6e26ccbe51fb172c182b7680de4b355995;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e4e2b6a540b52c82cd51749f24fe4e0e1b6ae33eac8fb61d5a133e6e03f51ef9238cdfdaa327fcdff51f5f572416b33c0373a25365c06b5ce40c0ddf364568d7a21c545af5475d859d0a182815a121a9368b374ed8fa37df6aee4379fa5f54213f319e58927a6d116d517cc2582f5a39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b5d019bff8998bd9c01a5058f4e0a2558aaa4e294ece41ac0b8e72716ae01da670544e79a27790c9c5b2e88a8a0fcca246a185042c652ac8ad38943122af7def35099a05daf0de4c643001edab1bf3d98692af43bd32c8d73910109f51fb6c658b8f868a118b9671876c191bc2e6634c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he926d3ebaa834536c03e0b5bcb079681bafa3dd944c26b1206928786fc430998cb4ebbe21db93d157ed9b08fdf0a64713c173c9a32094a1abd241dd4eb3f6cc054e2da89e1a9c1ac413beb0b1221ad5b6668b626d4c902dd33a1656931901487022490897b9b0c77bd1e111fa052dc7e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4ce73f45dc2cac73f511d0c52a90a2ee0be932cf6dd87ce204201b42fb7e7c9bb80d6976cf570190c8ca0f61a196ceb5cba2a2f8039ab0f880cbcbe5d7e40469b17b76b16c0f9213bd11ee011984049991a78811de722c85167aad2b2f33868831c88b57ed304bc538564a1b78830b7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f65345e0e95429066d6cdef00e764e3b2927921f6b22ec0dd908bffa76d710f4ad88377cd8bd28da2a8f907744cbdd4051818ba569907c194446eac8cc7c38520018830a1b9db5b89879c30b5f53e110c3bee1fa409a010929d4aee58738710f8c5b41cf457f43f1866cbd172c8bf2a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c4a40cac1353f9d563ebf75be8cea387ab2849617e3e78b424f3e8a30b8e43b8763925072118bd88ff92dcca7e0f52574efabc0f4d524f45820b996e502fc0c5093bc917bad8294d22cbed7d514fbf411c98ce654a1411cd02324623f4dbd4b07204365e93cedd16afa19ad0dee8765d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha47f6a99964aa3f7a59771dd93ef922412a51f34f22f539e9abb5fa21e5904e35eb78bc589a6dd587644d21d403e28c985e3921f5eb07b0a11140b6d0d4700971b36428fd0dc590396e033e89e331f4e1e3afc4e39fb52094e1161eaf4eaacba123794e5716cd4aa642342bebb3d42622;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h928a2fca7c40151e671767eb3aeca892a58b66a243bb3bf22cf02dcf313b91255bc8f0be7361cf7cb127286d19265587a9874bff0f4125c0b5b01a3d6cbcd292ff5114f4b0ac429225140cc16949f4a2dcf5b6e5b5c3babf1a5b83d449edcb1507f5bc6f476e5ea9f212cff210893756e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46560e577783640a217d426f85b8a9637ee9b7ac539d4f0709f9a3b9c3a6fdc7a07514b5e430fc630f752a5a5801e7e26748779111b1a6ec7a4708dd1189327ef1d7318e71d83b7aafdf21474eb465070206ebd0062f3a5908e5eb9c0b7cb8d4c7be5bb8fecce5d0d7812e3d402c1565d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h636e5714dae31131c087812caa8f1c6bbc1613b92f27bb092333a2e34cf1effc20db47f374cee9074f3837aeaab99be73d9bd149f957fb03567b74d9a4342a301160ef72adf4217633481c54ece9977d7bd790be3af86f54b330ba46c7199a34870d2c4a61df723ebdb4dd7d4458d7fbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdf12f62a7abea94628cec31ea52cb7cf621ffc2ac2a4d748294888876969c62bcbf05c7571de5d20cfceec288ed7bfa82bf76978dcaf3b93e4f66306ae5971a451e522e124ad529bda39e64c3d4ad9f9211a94304cdc367f403c036c2449383da744cc907ed646b56acbe79bb43fca59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2511237159c549f37d2c5904e787b82f10dcbb4bc1a56fa5f13880f046985f483e46f52b340edac3f2d588bd3078cc67a34a3e1c20314fb67e2e977b4f9dca20d4735cefcdd30fcf553fadfe7745d5d3a59d14322ec53172331bda445b39dfd88fffe983080ffce78ec13e0f23ab81f62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf20c1222ff622994ca6f97cf71eb191929c9162f8286ba143bdfe9b0e98b128e9536ed93a3ee8a558b9a4f50fbf85295c05cdbd49ffb92c2c6fe74cf04fc50db15efc478e3981472a0c0fa86199cfde13a7c4abed474ceafc89bead0c370b17c19c9695e151e581001df8fd41a3e4b00a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0ae97bb3f42bb6e467625a0520a52aa284cfa2f0de1cd89e2247c7fc8b4dc5f3f8b02812c49c0ebcce025a04ed6b87afb8c0138387465cfc97439f73559fb0ac1c113b9933e577e7eb17845da59f68b75a0d5911de9db559a031d38f9c19c7ae754390e4aac90b3b5a3954d43ee82c59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdac50a7ce8b7ce54edb3fcb99d7ed1a306f3a5817518a288fa8ec925ecc75e5ed3534d99dd31a70ef56bdd404bf5440316f0bb776f9cf737e5f9bd7b8e58630122bcab2e4b179d67adbafc60842e810f6850c6c5543d4aa164675df65ccd4e0c060addf432677eb30f5e313a6c0cd6811;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85887f6eacf352f1f1cc315248eec2048dc2801d105391239d26c182a9d4479efee4b6032d55abdaad7e63c2bed823f44ac2201746ea59d576665e4b84fec2ab0cde010300cfe9853d455c70e0693a98b2f9b400f07e1369f64e58a5a13eef13565a834b8efbe769e0f60444d6702c87c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8153ac861719db5e59deda97cf1a1912ba88eef53c2f05298710f28fd9b04dbd096bc7e413a906f504df6141b76cc1fc4e6685d9c488bf9a3e1f978446d284e5a964bf206a390f4f172c8e4995812352a9515f563c2de6669a331f258c390a96ba6000105e12a9c2b1f74f17fc8cf3ac8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habf4b3f120e839dc40cfd8f886dd15eaaa9b7aa80d85a4d5a6cb719f58bbf2983984fca432804bfa9d0ecc9c67847d282e97de985fb8d296743f272abbb2ee40716453d3fc5e83b96c38f1961b7f377dede1c5362ca1b3134ceced2369aa8752b5126520014c985843b0cf114b747e83e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38c82e27ed45618895092c3c27df53ebae74c07dd0177b9560093593eded4ac673aa280d403102c8a8bfec2aaadb1a5ed1f08ab663800620fb9ab320e9a4240cd28769d23a61b17feb55fa38123ca9b18a690d884472400bbfded97b3ed415f40ebcc7f2d6856d5164b376918589d6995;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h377fbe90a2e75d82b6a1d8686b8b54123fbfde83ea37d59b04458a28f0db2a2c2612e0fd8c09c51cb4540347661fa68202a8679b4217a9c594511b244b7378de6418388983290fa85f1936ba826983303f8012d9c69fcb65cfc0ec670492e247217f2d2214f0bebeb32ab285c64cd1da6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d1a58a1155e1176c6c9904f55768a1419bd49ba018eacfde44befcd423c703669ff2e5506fc530ef917d0f42467d49d05035bf4b03e87016897a58329ac879137f0c332740dc6bd57f83feab76c8a0f6a7a0f5ed9fe4a4586a206b34c2fa11599632a6466c8178da34b407bf193fea8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc9fc1c9ab79defeaa90079ce3a297b981792535614f84140d5cac57dae8aab8abb997ebafe28c8a27aca76696e7c3c81c26c8119a443f6523a2fbb4be34fe30b7ad9d157091b20d4847ac7380f949b73ee093d8301b22945ed2de7a73bdb64f3d1ac2fbc9d2de0f9ac1f35dc35835272;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2a1e557def117d145dbc3aa70e2f5741fd344f94678fe5cbd18352ef4528e3289e7f37479455110dfdfd86943151f8cafa8f3c87c01a63eb50d2598b0a044383e921dea18d9d1d0240c4a1b0f2393efb155cbc93021ebeb21759a7899e8afcb951eeccb2d9277d052a43ed16a5a8154c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8b8b4fdcdd61e95ecacf3a8d3b7a2dd5cd2d594c5f2dce3d6ecc64384e7dca3385ae1d931d411d2fc8e49c04126360d05c5c85c466f818744c0ea6a0cc297ce9a23a908edce2a87a21a74508365fa7303f8283038841c285163b26e3e77ffb4a77be28c8ddef64631d7f6cd09634264;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83fe9a95479ccbf4642bfb3a055bd5e7e68bb0ff8181f45a8d0091eeb9b30db6c5c6212f2e2ea8e88db409d5d8de7947a28d5b261f1692e6189282199b394a05ccc40999ef5cae8560f7cb416d7533a14de39ba5047de8d28f9e292e2528a7ec874527f4d6ca66f39c8f22a2646329b6a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91893642759adbf5195bfb57eb164380188f891b9c4f1942722fda3dbafe6dc9e35a91a1d38e5ceae0f84de1c765e011239a4bba45687904503ec82382d99adf7cde9a8c948e7c2a8f48af3791386e23591bce1bfe927ac7205b57c91779972e8804ae1ed5947f653e442c547f27e5df5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8eb2aa85c77ae2816996338b20771e54063c7448542b7b8500617658916a5dabcd5456b2bf1f3c5fee0490c67fd5ab727a93d1251a57c514b9975033aae82b318524d6acfebef610cd97b7e71e80932942ba3d0aff51bb18df5e004d085551bca4b4ccc5083598776ceb47861dab3858;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb06cf0fd7eef3ca5476d9452bbda2fed516915f8a1cf368568baa7fb0cd5ca9cc6cb8df6032fa071b23bf4e8cb9fc17f83f1616580828c51a969e5ed9c5491675e1b4493bdaf1e3deb0a8da64f30fabe7cfce42c75401f9fea1966be618d39a0d0430847b3694121097d640eec93c2e69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6adfa90ec171dddc2185de0c0dbf62e2c109e07cf9a098a72c8823dd3a2acaeca73a07ed5bb8446d486a892c982cc266df15f0edc79620d80b5f038ff69c3bcc8052a756eebb26600ff2f5c4927d72c6711f17b1d12eea22a8ac6714b17a3cefc7fb00add3de524642c5f6fc9728abd4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5a39d2b1865ac8a0816f2caf406e7b6f0953b3b461ecede3a144509b8e7001f5031fbe0641e0ab0194980059d16d0b439f3be0da282e40c5f3f8fe26607f9c7f4b26df318607b19f33783dc495124f0c7a691963e1af751378da4f9f0271cc658e453a247eececd803f38b027bbd0c22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bee662aaeb0ff9f19df63dbe3817dc4a9c9c602078313ce06897370f5cd6f567330fd5f52bcaae0ecc12f04cf83b00dd8cf037958071e032d49b02c1b2e949cc7c2e2e186acc592e90c37ead46aa30f9e83b836dbdda6caa444b52ebae57fe488889f89e11afc31d025b2cbdda4bfa09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47e7510a491da85cb7e6aba4d70ca6e0504b8e32b320841d6f2fc1ad0d6b9973c16181b6a126c703b921e9f2353cf18a0b2936e762dc5af536807ce6f8ce9b4a90024ace260307798614f6a1199cfcdc55e8a6167246a391d4c9e6cf1b988ba749e5736fb1d5965e03a3de62261207566;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd8555009ce528c52438d24ad595b641b4262b41ffe6fedc298968829b61eb784e66bf63d3c674dfaf62f1c19dfc7621211d2ccf1e62065f5e26ced63e590e0c80e2fe8a71af8f5b898563713952ea8e4812ce5a8b34964286e3fe424ec3222625cfb998668f27abca30dc1448cc847d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb62a4069137d911f6aac77d135164042a5a4b535d3a799e59670340188d75c9b5eb7983630f8b493d089bd9e0ad35b91a79099cee41f451c31be7cedf045175c621d329092457e8b0f66b71ec04220589fc94964682a8e3594e2fd3275a1915cd1366d9153fa33aad443fb2ef4bc54c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7931417fb7faa440406e0e141074d0d4b94f34253fdb810ec5ca218a8d38a27c0753c9bc626eccd00742c5e95ec4d6d68246401904beb5f7de3384781f99773cd46fd94d50663a4f96a061db76c7265ab2acf5ccaa75c1d38afe627603a3d72353e2b69cad58cafb158c857cc1f1d1ca1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9f23648642c328c41b2c02bd19e5729e19e7dc5aecb1095c0d14c34edaa20bbe1655aa94f3db5d972f518196b65871e147ff150c91efea375aaaa7e25b1d0389d1487f099879490c0c6dbb3bc0b55a5a33453a4f344da870232ebe1119a361cd05c99ceacdd15c3f9477d41771081322;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2375173f4548e1712de6d44febd1d92bbc95852802f92d2e069113761642fbe8bc7afaadc7b02b15cfa57bd1d93b2e29260ea39caeda49a980ec952fee09571d4278848547d7cba2ef6d531b90d1f89980917dab2093b160c33cd97f12481344fab160323309aa9dc4e0529428600315;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86cd21164a23a9f06e0bf50b1c3b06d4ea3deb706ec439d0b5c555eb371042b6727c675e921c7fa544a89d4d25558668d5dcc15d860885c99dedcd99161d3d1fc93d954f3efc1979ad63dccb419f7e0b955e613ba7eae2f1338d35aa1abef0de8964d397ca8f6467006f1c9b11874a9c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fcce44b2d7556514e798e699dd3ce98ad4ece8f4aa6a0d7d0f9be9f49c15b919b0451e5b6f21b3499d6a55eb67930c8d909a0c9fc33bb9053e05e1644e12fca9731357bdcafa05187dc76da6e3c59ca14305a336122737c17306c3ddb0d9511447fb52af2b87119e15fbbfe2e05a8f39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7a0fd49702728156ab8c5e5ac4b2b61cbb4edcf99b62cf735225f61317825897905692b7fa64e157e1aaa66b59e3212d90805db7f0b7e12a670b7ee2d449e3189fc2bf634f5510c4d39673646160dc92c6aab20043ec2b84223f9b5582403bf728079a3ef6112eb3d406d146d3874196;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h203cb6840b82cad391f4cfa0c477f5b05760d1284176ddd28f7df244ea2f0f4f31e6714a844c00439027090c2ff893982240a93ff20aa70300b7d22039a40c32121e8b00a148330383f4e8bb6bd9d56885fac85f9d60575a499faa1382a280c0fb1bde741d8b4b47ec74b5c7a4ec91bf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f0997975dbeca5fe96cb7077e58eb9edd2810b34fd13eb286bd32fabf47695812b10ac4b2c3083ef34ed5d7aaa1a04adb451b38b91e369e4316418153849db855ad7c8da873b5847eef9874d6bde1b3bd48a355c3ecb0d139e6f93360e208736d68ee99713cefecc5bcbc949d7e58c8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6be6dbf5c531645a661efc56ffd7107038b1488d6f4267fbfeb26bc5755b48dbd344c13215c5c41ba289c0a0cf74fd8d6d7532f1d99eece24acc4c1d99f8825e073f35a6995b2bc908e299d9e36ce4a26006cf5766eeaed02eebaa1773a6f454ae25ca99c7b3ba5a421a1c9b87a2ae929;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f4474c3a27205a61384cd5f98da632b7b62209ab3bcc1eb9ebbc8114d2d90dbba2e0cdd41f0375944d1ec4f9fafccc65d6c0088df8d5776fffe10338806be8877f104c522b0e1d0da47152686084ef74ab75ea54375b4fc5c429dc5fe739536c6d2eb485a6e87ebfd99ea8d8c492ddf0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26bc383b2cde58866a4fc12b8713de748c44c98b82edd7c856b8a5d182010177fff3562111c8a6288a785f753554218cb9b1ef07e6d31066757fa4a9ddbc3c0a4eef0625a8968b82f685b7cfea02b6c8bb088b20b2908d8454a4c3d95442a6b4fa89a31e6717262c674f3a40ea549fcd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf306a8953c7d57d7262ca3a66ff489d6399c129973299bf5ff3da8a8751ffd11d8bc32614f77f9ca9be3f2c3e40656d5aa907d18174e8c910bd56e07663091ab4e9cd780be3ae5177c21c5953806e3cc15c4741549c6035f703ebbbd69dcf586754ed1e94baacfb65fef59066e842ecde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28e3bf2d39c1c218fdc7330e1a1100a25a7927dbd231f5a62ce92a42ffc9303258f3a61d2273f54957063c919844975a3ac70a3c3db782b409d2543e66b4a93f707b47c3219ee6d9e7f61da12c770c39072de764c2b9bcb08be363f5ed610bbe66e233e6dbc1c906a171ec8899f2e181f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b9372e11bfff1f10a9b121196893e207edca1ef3d24db02845cbf822141c88a2bf7e3bfb9a90c3d4ce380432c7110bfc6a9ffc56acb79507b3166572a4f9efa8a8e6366eaf70872efc6f301042883fdaedb6043d1dc64cfd3acd4b6e7a045ff939c62976d0050bb0d01cce7010383587;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd45fc8105f262639a38cf60157130d87f0a683170954829ac0b1027e40e27540052b46977efd67b8a5dd90dd34a74f88999df30d38328b6371272fd1c6158bb645f47772314b5c1ebb52b9b0a44df717314886c0c4e546eb37cda9a04d8ae0c2fb02669c1981e587f0dcef6c92238eadd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f614c996071c838b9b580f05cda6256004fc4f48e00f3b0acb1cff5096f50e4535fd4b77340120851303e7fca459a7e902ad0b44cb05dc8ca3dd721965739020cbf0982bb4a7a865471d71c6c6d87991c476d2bb6d5a974e56d99a2ab5711fb9f86854eac1aed19454b85258b2c37b21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cbe3992716e21500373efcba4a45fa54a0360ffd7bda31011bdb8456a2dd4abd31244e36eb1eadc68cba8a60ea5d7186830cbde072e9f18d718592f71d0f83dc8bccf4d8e890b0c4060292d4ac8d1bd3060980c033ca8b90b1352b7da59042e417b5fe113d957f04af7fd9999aa91c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ebf973332e901db00c5eb6d9401abd1d97cb7ed5c3b7d0c328b0c6138434c83427ca6675c2515514dc365d0cff0055f307e12c2a241e16840d724204f03b0e0c73ec1ff10343d388a9c90510a8b363499fc263876f9b7a52368bb7b2b28e9a3072da91a36e671e160b8fac2519aab177;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14f5d25e8fc196d8200467a1430116f4b5b9598789aa2c73497e267459995141a8a11e0e826ba80d25027aea4718fbcd5931cd05375a71583508cd979f94d69667106fb4c252634c243eec2a2cf2f2c08b6b87e25010ea02d35314324c98461f991a72ee9f64adc5a7998f870cccf3376;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1355d6020648bc49108272c123e5a5f6752eccd77a4adc95563425075f08cb609af02cd8bb37c4be230e1945957f8a2d97422b145d3e24b50df75cbd6a2a27a031a88d8baf2109c51762755c158366446122d307acbd552272c1fbce648fadbe168efe754c16d78db4de38bad363845fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c2aec210124aa91d92a643e5e3f83fa64dbcfd3262515f44250b88f875a963e55eea8dd6217db7806559321a6efc865412b66ef4e2384d97a738beb68946d613bcf258b16e96fb02226f104703d4589cc002ec3860abd1dfa2f26785b5a76c5718f30235c09ca859a49fb809bf67d0ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h457893ebe027a9948e2987fa63b5763d74938cc729fa664826dcb142093e6fd102f35ef85a55ecbc527b8cf14b3111f2b14dd98231550c67db234195fe863a4210a5e1ff6c88b022c9af7d07f40cef8e39b98ac23c185aa18bdbf21ce6c2751a3dcc6215718341b503bb1a2e519a2bdec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3182bb3e7050e3c5dfdf430c24a540a0d47a33868b4cf4d3c0f9edacf65840bfc0eae94ee5a8dec7b4668fa33c1d06a0f1aa4f3c1e99390d712806aeef9f676381a03704312fb3c26d048deb46633ff8f2bd51a71fb1fee0cb7a41a13048eb73bff3e6c77759ff5ddfeb22af6d07f4d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40c7a0c33fdac0187ff03113c3ab61c8321681a430a138e39ab10709b7d096ddf7fc13f7f399d707a3a42e58fcb754073ebb264d58e712cf71d7d8f2074cd49524fa0d5745de4369466034e1aeb8845048d5fe9a08db4e1d4461e65938c195cd3fe58b59980bffc7d831c1960955a3e3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h852f9a11141cabb819e9b42dfde1c589f99b575bb8b3276d61d7fe0698fcff8d58e9988a9da3666e32a0fda187db0c160c0f4b803b43a92f07173e5c0b34bf18f56778c62f61c6679787bf90c8e94463fc06202d117c52ac5209732ae3758c97c6734c3f02adecc9e532beb24ec78645a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d8259bf862bdfd6967830b8f21eedf4d7c1651d31cb848fa3cdb8b04943d0e7de50722b0d349507763e994985c3eb043fb42a23123c2f8764d3e300f4a10c6cf4fd404e099afbf8eefcddadbad57cf80dd8d05710e1af08134f8f1ae0ac38c46f8988f6dbb9271cf6900ed3274fec8b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he076b241c9afdb4e70ab8d487da9d4d295d799502375a91740e2e4f656eb268f0fb45433fcab443e06c38db7e969d03cca7a714285ec5cfdcb039b706a2781f0a5b9c4bbe0c6d88b7b332c6b697fab8d33a6249c802fbb77af5bd583ddfa577183f170f1d9203ea1f48a8af733da1932f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10be83a9d69bfa749fd2d51b5394559dcc0c0a4f86c2a74b29496f57dcbaf567d7d3768b5eda63f1f842d6f4a0121fc94c2cab09fe8fe86736f60c02e88a78fe4b9d3436448bcc6a8de4999624b6750dc6871028af59a60c358578c40a8d7e398bd386ffcd959a216785fe723724b1ee5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb681191e9a4fe29dc1ef9034087232dac427ce3573cc5c145a5ce8250196fdfdf663bb9ec3b15018ee14fa8751dcd999e69e71c63f6bc6c907f3da99122b0622964d70025e1b1dd1fd06fe13f2d2a71c7b15a5d058fc10f340b5676d4195fc6058a35729540c64c475de45a4dec5e6b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc221bfa770de3193a9a6e904aa6ee08925c52c8dbdc71322c1d146656399e6a5fb52302b0b9c5973a7b455e0e0a6aa60e399d77dda1e9878ac725f9e6752a0b81d4abcdd75733741a088861e48a8e7921e19a780eeec5b9c96c706e7bc9dc2024895c0eeb3436a6c29b37d8c1e0f39bd7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81a99fe58f0d2df24a2c24037eb11beba6d746ce60b0661a6382df8764c46237dc5374e5f64156bba2ad14bd43ca6353a09c0b6d7e87bf9075cc2f99d0d217afe71872feb68bae149594627b76dedad8622b775b765d900160cd0b86235574fefdcfc02603cebe05aaf327c9476fe5ebf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c7310d0538c94c53c5b12b3c7ef7fd647cc34f0f9a288b3c90375b88daedb826c434a78bdc06cc8bcefa9675abf193849bf5b31dac94d7ca63bd5500d333acb27c2c1a55c2be12a6f2d4d9e76a4a8f709297e5edbf9f0bf493cc07cf656aac60aeaf4a4b4f3d73f5882d03397ead91a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cadba1662d64fab3d892677ab23de6a74c037bc97c28d6b724c2728ca2fc1ef6f0a47a3516122a31819452c03fd1186705b2c7a796cba398df4e14235fbf301be828d2fff4ee1c3fce54cfa4cdffa85d6046d63ac93ed1af6659123b288d72843824aaf44add34a9a99d6da5b9b5188;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99697827384f273a606e23f03e1adb15088b6ddf39c472289803d06f45df5f18a3c09bed9840022630f72dddab981b83614cb2a56f15e444b1d6512a2ab332d4637c4234f06e38a7041b72bedb4d3e759ba16c0256705d8a29bbe721bd3c880acbbab2714711cf44081f3cbf9639caccd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd82e46a3400ad50799033c29af5c0a95a92f763f80fa4e7227585267f4babf8fd5ccac30f986283ff01213dce1c9d8676a4d9948af96d515ae0c301727fdee7694593b0b376f5549bfb2097aa2b32c67d90ec49719900b20778b4bb1c847077da080a8cf0e37e2116281f7f3064430946;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff7e406f9c9f2265bc06061db1c69dd6239fc93d8c0f6c5be166776c220bac492031aae95ae2939a92e25e92a09e2783c753861c1852b115fc809e259686ac52abcd0958ae953c1f8826508fba911398e9600ca97345775969da8b5e185f876800169c52c80c0ba1cc97106c3fa1f2ea1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0e058dfee4f3e049ee10cf651b72dc5bf8903814686d7dcbe5bba247b1926bc952046ff1a9ab7870d54cf7993c1115f96c7c8963c66122a27260c74a52c621f32984b9f2445f0a0b178628f4f4dcb7767a2edfa8cb65b3309f032dd8bd5618a5f97feff2213d8c81f6f9a9f332ad78a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2cdc7dcef1cb6c63c4d3524f69dfc1e6074b47fa559e6fdd24b9b3f4c37747914665cc4aa36f470709e01e4074094d671f9709223453cea78f9901d033dea71326cf9b63da79d08a6163d57a083468ae2d3a2d7915895f3c690fbbd7fb1eea2f318fa3170070bc89ef6d07929dcc6864;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fbc0b7014d55c7de4d8db6c3ac766b4484072dd91155cddc59ab9a5523d634f980f6fcdbdc1b3a962f11af51a042585a44f57d5d47edbb6489a5f3212af49784cbc29ff8ddc775aeaf24e9319189bb84db56eee85348a84ca9633700c6d0a46316e6ff9822640eff5a5f17349abe9be8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he78608e15a5ca22102006f286fe6e0b6b1812f20fc84d3b70e870b3b2851bbd8f638c4d9acbd580e0275d0178bf6c1bd5a246c31488a487397cefea2b528fb05ecec940cf77667ae329a49cb99321fdb1bc27deb4a70df82f08475daeab5ab6f31cd3254985db22ece223fb4428b5d139;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f726ca70fb71fc83b9a548cc847617957d23545a8ad185b9756b50c38010f9626aa53847f98104741182128bb940d94babd400517aca2150dbc5a06dfd15968b366d0843fa91d119a286312278b6a1dd1a3c95d545457c72f57dd5b6186f18f8d3e6c90a15efa0651976a2ffd56da7c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19ee51c3318e5b1a5254bac73a83d73cc6745ff4b2a34f8ddf326b25c96fdbeb47c03775c92f3e62f0bd5324d972a158ab072439450bbddb626f25306386b6bdfca81606ebab4b7ef0c8bf9931cc284af0b30acbee577cb02c4b55cc0e8b80c12e0c55bfb8a93be2fb3aa4117f55d76bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ec296761682cc8ca9a87c9616b03c5a726681d6877ac876d5b47ed1e006371081b714eae4a489397497eb4b9266c2a148ddb60d6668e718cbe0745f07e885e0f3979e3b530d1fa352c0ad9491957e93a4a57947d049b2d2e9b9c5a24810b09464086f6eb461ea95c5ee0dc6cd8c3fb35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91571b4703162bef09ffed3da2c74f28630620cd4b04a0a7dbea43e98d483cdd07bde87478ff4ae5ea2afd888fbf1892c7e1449212fa17dfffb7292d592dec399edd54d27547ff70e97cb00e0053705de0584a7014ca67435c08a05ee46204e6a4345c4ad4b97a221784436eef27a8902;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f02985957514a8214d6dce80123c1c21e8f246b2fd9f5c1e48a942fd58120f2b9b6550a07d83260eb11bf5fd6d112e9cdb311de4c023275fadf8f076737662a1166949c75807cd6f5d042f3bd3014353bc3ad64de2256c4c2c3744024e891c516df5f67963606297fca7a6f6244eb585;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20ecc4b544c7c5a6024bfdcb8ade4bda69ff112f76d133df86d8eeb957f84a6670df5dbdbdf672db7e36ac555990ec68f94b1c706a32c02ee9e7492b13c5280cee9a0a4e7019e1875586da20d89e66e22c03d66715e3f366e928fea81a5d9939918d38adcfdcf254da449f909170fb0c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b20a621c81397b57e502ceb22dd35e0b491afaf284ddcf99f92a83520fbb09bc33127dfc59e10dec3ac8050968975054c81159a8e943dbf064d80a35f5db10a7b3ca5ce36fce8ed5220daedda1e9b29e02a1403038b2aa6a2f3d956de30e35ec3956b1a3dfa0e3351ed4f7cfe13806d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf1505edb5c8e7c6e00f47c3ae080efa9e4605892e3d8b7a6d3925028f3772d91428afe4a4477269ec676400f5428bc36db105c0cbaeb2594aa71049f7d687a3a675e4a58d0d61f45756b06a0793d2e74298c99ef58a173318daf244bd7c14e1b807bebff71e9d3b5fe527e91a8f74452;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcdb2e0280a33a295e78f367ec9a144bd71b19841aa0308b64e4b3abc1f5db5eb6f2644f40a54f7cbb75c19cceb579147053fc901c3d83a8beed74f14882bba3891245d1948dd8b448687cb19d9542ac58536e3863d6bfdc218437e3167f36e388cf1dd08eec5c4e00072041b373c3c71;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd305f8461e5d714833cec5e48c3609baa7175a547fb447a81e44e8769191f62d05feefc36739a230f4f178cd9c7c19978a04339929b9609e3a007df021f4b8cf9ac89085ee143b47911de9c79216b351c37d67f1bf3264124d328225884691544f9e1683f65dfc94ed1a493197ebabe2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33f7b10ab65fae05a2aec0610a1588f515a9e06c6653186947f58da3fd35c0fcad6255a09304bf2b884d70efed43e93dbce4687348a095b07b8433c8d5c488f3b69602f711925c622f98768501ec38d864fee9ae1cf00cd90971e160b2cf4e23b8fc41efbac5408e8dbfe8556b7801f8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd1fe9b2a29ed74630972ec95216033c196614779f171386d3be9eb5bcd878f1dc3437868d521bfa0fe016a77c3bbc24b11c8678e8dc564d3650ec8d99ce97ea470470be3b105fc597c183d40839fd929b94e261bf2ddf87b944d766fe36a5747dc0737faa6520e4413bc69d657a39045;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5141fb9c8810772f2ff0a6745969cf20934284ac298c573fccbd1d9dd3b4177c3e6caf1c83fc3dcacbf0b2f83028615a4e61082073d866f9254743c07b599674fd5f04a5cb5c7970f5944bc3783c93b73d9c4627d4863c72b2b67bee9b4fdf0d4bbeb5c0585cb881de5f968f6f547d118;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha97469556265275aa9b099be21b2c2c7a217525e7d259db9208763d54431d82e32988d775ee034a8f1b955bd67efdfdf44af50ebcd53dc2806fda00629081e195066bfe19de83cbb3c448f954b840541200b1d28a41f299f48f801e8fe419af1b0939935c86c769f99e8860047f77ef68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9599c8831d9f187f534ccab9a7b534cf8cae55ef884cba233f7f5fe0f5566efbdf0d263da266fc6a0853a9093052fe8d6e9fa3e73ce38d8018d0fb065051067ab4659c12cadb80830535960d43723ac6b771d96090fcb5e99a5a4dd7818827c3a1adf7abc5d18146f950531b1afdccaef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40560647914455594bf49333447c95fe6f344d6aeb493043823fa1629615f1dd93ea22d938db38834775bba581755078aba5321dc9570a7f2f2f9c85d08b3f5a4e7107f2389970af14ed02a24f2729e6377b30c46f8181be5e6c7b0bb20d51f5c011a0910eefeb10b46bf7eaac30fedab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0f0dfb90998cac83cde16896c1e6169662e93c9f910829e593d312040ae73991d96297ce42dea2c3b03b46933f24c3df5ae93a9b0a73d1c877995678c54396c8062cd8c18eb211ced793f32b7840ea74855b3928a52100643918cd5ebcbd4f8befa1cdca0421bf393b767d714ff6070f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52ba1dd6b7dbb254e9ffa8ed409cb5ab079d7d1157040496bd3c54eb8123ac5a42c8c5fd7b733c367e3ded6ca4a315958df31beac0018d5fcc1e27cbc9e74738e58e3bb431954c8d21960c653c657f2f609d27733d4a633bc941d0ab6b29e17d1846f8ef029c2ddf735679ce54806e374;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7adda69d81e1e655ca3f8d9d937a0b31b5cc7c03412165c7fb9f61115111c75e3a2ff328c1d814e8d5e0ba3786fc85a0c3d8e5d67b7feaceac17ff20f9bdc203d55ca288e03f571cb3ff8e1e35064104a290edbc2a39153980886d811a8092b4d907a431dc568e122338604d6aa9e641;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6680304c6793a34e820976a01adcec776fbe06224d58b05aacb95b80845c8f4fdc447aa51d8e0271ee9a869c8db4b99d5b30fd33607eaa1d9cbeb7964b6f39e9a13aff6cf2dd3732c9aa5fcc4364dde00496a56a325ed938c4bc097190ff7e19449b074f57de058c1f04c34328bc909ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8aeb35d436b46d15022b06e6904b81c574979a4f0482e81effa0e96774ba368306b9d93b03660a8b7effc7651cd87d538c01ad47f202362bf0a81de7cf34b49d51797b9198ca1fe5b6e7aaf7405b9560988f9c62ef444f96b080161b66b21edb8fca07f7a16ba0ca0ebd2b991fa320024;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2acb241abbda0ac85645c87e8dcd72e1bc49dd030baf7d11b180161a5e6c1a331b88c983e5129c2b2f0a67a4047fef2ff8c3ec55469648e492827a5370ff3cf6f4292791504e981c4b0d7b4aa04e0fbc0e3f7893e92324f4b48d507bac80666383f4cacc83afd0085e4b31c575256f51e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf7c21203f0032a9d99d7f1f7980e002105a6a9f7f8f875cfc9eb586b493f100fdeef3d75e602c68768643b86534fe17be250f309d2ef41553dfe41f2682fbcdbfe4c5a4aec8753abecfa66adab7829ed7ff98f5b32fc0a5ea8eb40690720af32eb440cab37ea58b7dabaf52ce5a885bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38057b89fb389dd5adee458381ffbc73804a998c3f151bf068522fa4eb734d5dc9350b100e82cc6c3a809a05a04fad4a52edf6559c1cae508309646397196c025222cea419bf65755054dd42f50040cb64626036fd5115a19ed7cd23ca4b0707f38038387787a5749b072d22ca8a48c86;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76eb0d541a660f0f4cc74b1ce98959d79856813665c5a90bc37e118e7ac4939fdd72e702697b362e46a7f34f9eacaab8624f9f3c8a2a92a2fdfc3cba05ceb6586ec21799dd866b59299d0b5b726bbc2dd0a5eef354319880e85d5142aa9cde88f1c4f62269099e5858d3b194e5b9c8f95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f4e7cb0c7adffc36da411c7ee23185ea308848952a3cd673e7c22ba266508fb4b56711fbed759651d15f3860d52fa1b647d3dba3108384c40c22c64b558d72158db20fac545c9afe4690eee556354cc6db6a199f7596217c027cc92d586ab700b63b207cffb9260f99d3f5d551a21eea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2494d1af4ab4ecab1511c7151b006113b35b5ba6905ddf83db0062fb8fb720be7c092b0f45c8a9e89b41bcda2c2d5596fe5d5c33b992c78584ea76b0fd14d1aa39240e0efd4e329774ca5b7eb478f0b84be3eec9f8e1c3f99e7211335f106c4989ad5ce5630cb34d89664369bbb065486;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b65484d3aa6ac1c54f6637f2864a84c216f09bfeaa74fc568cbf7e5e30faa4dca7eef34102f3cb3d73390ade02671c1a715741731afffd4a52d091c2f5059863ba96c4ba92ddeb8503fd6d54f40485f23e845ea95f459434912bbcf9062e49f10ff697a3840e7116ac812c403c0a646a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccaaff773ee90ae533b315df7622a60c836620dd3a25976012fc82845f53e9cea1d34f3adc74cc1496ec7100c8d7d6a5948b6a1b7e4f33dba000f797152b6823f590d14d5755dc63433793887e8e2c877b866ba4283cda154617e34b256eb220ab6354c080374a84fd9d097df13f9ce13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2107a5733520a603ce2ce4b6819f0158dfd502bc1d84a39e97599c2542f751641bb883eb648e85ad73fb31f95fec3c5e362617da4034821127f2682076ed1160ddcaa9faa34c036e2a5602ff95815f66945621028ac0f4b7a1ae5d3e8e65968cb9261f102f5e9fde1ff77b6e0a6357253;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc15476b75902db5dbf5fdd569c53e8eb15b1bd59c92a0192fcc1b79899a9367d5ae54cb566b958d0aa204f0cef75610c7dee05a6626b5214768065c977857e6d8981fa4e60142b7d7f376fc1b203813a699f6f2241083b387765a91f2cf7a4645fb01407493adcaf740c73ad93674bff5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4c95c82d1021b6945ae9bc0bf12baadd8b8fcf1261f5abc7af86ca2d6522786befefa012f254035c5d2e3495b2be7a5e691c47116ec554c9a9ce571ad6e1bb54082504bc171048e357f93d8cdda5daf8f005c1ee3b0804583bab03706a62b8bc5af749fe3cda6db8eea51dea591015e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde6718b5b55d9199fc91b87192550354a765b6ee4c815ed7dbff518945a5c44693301e2cb9c2cf62a5312471a2371e4ba44f8f8e7455a075de080568719e98c8020b49105cfa929104af07d544c0d3781d2af96f6c241bffabcf62788c10f7fea062bfe3eaf23f332ef8c4cdd08eab4fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ea752a53714092b4939a504ba5ae10112ec287d1fd957e245104be712c8990f9328ad8cf34efe49a82b491789cc95248eafee866b657fd296c346d0d13a936db832a28595ffed3e575c7c81486c6193eaae5fc4b92f0df60b2e1af93d2c43f021dfebb545ad3868a48fb68dd9965510a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86b6d6735bf535edabef66ef1fe632a3b0945de8adccd305ef4903c1369bc8a92fccc74b4a0c10485c51e7884d1efd44e23cc1d0916ccbb9ba646957a5b716b6e1ef657adff0b3261c4ee5080f6155b7b9576e8453435bd2effadf635551b5fb65d3d0fb301df43ff3966523d1cd26413;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fe2a6d7f7741098cd036f2cb481d9621a6a60ad1a1e929d2229ba84daae1c3225909d2e9db2fb1f1940d0de98cb7cb577ad7a529c1e587afed11a3f33380baa8e890bef0580e9bfb2ae4cb829837fef2010b503282b08520f3fc3bb168241888615a6e80268456cd9570d11d68aa0a2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha089071966e90ba3f2b259f025c6a90bde50d42270c900430c2cb8e5e4ef7e2094f0fbd2de60d645346e263d984c0e68a60a85da7bed6ab263487679d238c4f4377d803263470509a18dd126411916dcc8098ae677acfeb45265bb063df6479bf0bd5e4fe0c0da43233c0283704ec770a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he162739b688ba6e03c9caa4e1405f5391f883d764295986024a1aa07a70a043280ea9215a815e31b68131b45baa088c818f543bbb21c0caa9e18d32561600a88a05fad6e6405d29babcaa68ae3b91cd5bb9ee297c528a06d7ca5de9dc99828187c9a93ce75cc23095297a22bf1b62f554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b22f3ad8f132cb7628decb26722df626438daa899e0b9c884b974c47290332cdc017fc40e25ed2600eee5092e6bdba6ae0f79d7e1da3ccb5a56bd54aeb6789ab510a6c68e2532a68ec505e6d9aaab22981fd7db2ff7e0154bc5bf13b82c2c05f5dc49d7c4fddc62c8b56f27a8f4e3532;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec2f856d5ba35a7bfb43ccd29169230b683e639c73426ee3e14ccd30c02f6e7259411cd9c248d6afd6f380ae19c5aad9d70995cb06489f550d0aff3b703a8c9d4f2e2f98b72674189c4ab332727add117506e64f44db177dbc3b9e7d879a40df46e2e81e775ce350314fcf70f3420c0cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74f95ca895b4b7b7fc20760068165ea48651aed550419bac553eb8957ae2ab4796c4b01dcfa87c0379d95a880f7acacc49a72b391677c051bec165f57a341439f41b2ef2d2e9ca02f5fbd59d1ebf892acb5d331b72b8607671b1092ae5be940f821dd8c45d3cfac1d665d591891eccb31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4eafba440d5732729263b3c962b78b87859d9417aa7a36a201daedab0786e100681475a6759440674f5ce0b14359d814cf402ef564d03e33039e4aae8d4a952e0c9f56d94e6284762bab522df13eb3c6575027c0399724769c1bcff861adbf599ffc70403386e004f5d0e2f41b75d1d31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58b8162e99a00297f618f32dfe760b9fcce6292da5e37c14100173334d1342bd856c4dbaed095c27ea90b4af550da51597a73bb0ab8467963a5be689a6ed6f76f819aaf626d2eda3dcb903eb6b84b5bd64cae0b7c4c27103e769ba913e0d7ea052191847f1d1bb167c26915d73a137bad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ef824a56cdf337b8df1314298b8a5edc975aa6aef1c64daaa64fef8e379c53c328f1e98bfc27bfbef09115f412c08aefa29866343a7d5cb36cdb3e2f593c12e8350c0f7fa4eb7af5a57ff2dc91d2a4dd6b433b24e226ab689ee901a60d6f62da56ecb627e2b91ff57a6173d192562904;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h136406c8f37f751fbf5bc24541465b9afa36539370e80f25b984c2f736d7f817e1d9f61519f19aac7369fd28903fcfe51e18a4f79968b87cf250547cae0de34f23e9c1b184d7629ed2a66fd6431c9fb9e220ba7499900008707244826c541e498e40434646a9de36e9f7aacda95d3d2ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bb600c7e76a02b7a8849a888b7b434917e76c76ddd58aa6797238e14293c4c899fb0447aa7fac21b53cb4815cea85d2689ff8f054d3f98f6ec40019439b05dd98e07de960924c5a27e26e920f747c20ae744986aadf61edd4974ad934f4a2bb2e119a29c11c32ebcb0da2de642142a81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b9f1056c35cb2d6252abc78d94a747fbdd51e25d50a2a9e3f8811546fd16a105e6cf04bf468c3efe470a33fc8fe140094e695f51d2e545d7a146f5bcc137db591bc6b238bec7df00b3ec450552da17819112c0557a19c28c5cdf688387ba3c86feb2475d397f0d61b03a373d694f3e3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7136412ff06deb28f1cdc2df5b7e2811c910a2bee80bceb16c18f599f49f890bb920439efa424e89dff3d19117da17447890aa88bb2d04db089892a1695a5df455d14bcab0b2c8b0f513f9113fae367eed237c9236e5b4560f96f961292a18e5fc936a7a734e5e75f9f8520b5b77372f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e8cb9dcd763ab4cef14a4f05b43ae94298bc0f8ec6a570cb5bfbd492f232150c5da2c3ac26126ce7b392b454d94dc0514c396252861ead3e25099234f8db609036a0e2f97774811443e9716daeeeeb01c53ce48a1da9ed4214d16f436af4214ec6478b93958ca48420c6f5572c0691c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9749988bb37069b5f6e8ed8e96a40de92fc0fbdbeda120b87103598f1cbc64b89b4aeeb82915b3c40788461b825206ba2c65282bf8e5f0e1bc1b0dd6f086e512dab0925e679749b7e84bbba6c845f377fdc4bf33d3c40a7e0005593e6a2fe3e792361321289c7b1036bf5d755304878e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf025362f761c48eb7a76b71ba3131cf483a23e79df5f91b0d1a3e7c7df9a957fb651d31d558686c0ff3949de89accf8c4124df59c579b3703f7639f77d1157840f575c286251d18b06792309ddd5f0ba0820b993143e2af1c8f9248b9d06b72770feb64196f3878e69f768eec34bf418;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fa54af529c9dbaf84f53f7795ef8c086a8b45aa11367c7660f82649aa4a1a519a4cc7d478417c006af08692ca82aeb7b4427452281a94f09bb76ce9d5704075c977980d7e95164a09254608531549b739f3575b2111b8081b65c11b242605e607d0c14aebef0fc32b1f8a87bff24a8ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc24d919640b808dd5018ac35eed7362657111c4d70b7869122f8a1084e087c293ba80a756eadf21f89cfe1a3f36763ea92528ded4bdb332142ff884973de262009d472bd659c90a35886bbf5f4b9e05fe8587522e20d9f97bca68ee17903081148232970b71a6e09db45d778ccf793316;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h416c6d53d6e3d891c4d6fb7ddd82c079f4b8a5ee893a207d0d32a2d6f3b73684643dd8e138a81e3a52a3730a953cdff373b966eda359c6b40ff90ce91069b50d55d7a617461b41e8027f7d5905ae2cb999d01c2ec84befadb4d3a997da8a63b33b75c9f1dfd7d29ab3583fab7b3593c20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4185350ad7ab0b3aa45e0227587079c217d632e37c2218461c08d0632353d438fbd860829d2d9131d3ed4c56b7ecd11e017cab63cde62e8db0ee11c66ec711e251d6c2e068c2d394dc4b9593afe01b56ffbd4d6f7277af9eca940aeaccf1ce7280e0661d1abccec752c8176a4825a98bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49cbdaed7f44838307b94c883558c050ee8e04c6b30d6e2fd3430c766f2c87811bff724b8a80a68a1d0b76b7f657345c1eaf7e1d597c4c182f031ce34abc6d539f49d25842a05a20128ddb93b1602045c2b58f2e5f518665894120020356f7661c0ec9588354d7d317228273605854ec2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89e9404129ca04acca31d9324ec2a6b7a4eaf4093ee50fb59238595ec0d50a2ac1857369a8207754f3aae4820b557ab0e5ab16084c6d37b7e37d0b1e9298cce4b6acc743ab92eaa29ef0dd60fe1de9be356c01b631beb34283953a2025035d86a58c039dab17d0e171470777a8a4f245a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfba9d399b2356628f4e0513a22e6289c19543c05d6e88726967f32ef0c0d12540e94f022e60b8e10401ceb4d020d8f4bab403851fecd3d7404305522c8cfd796da1c62201979675dd39bfa9c0be030dbc25973436d266fc0ab232e885c963d123a34c5d8ca1e9182516060c8e044ebb72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he40a6137867548ddeb93b37486478f419756dfe5e001d918190f158cd10768e3660ea2efac9bd9728b4925d7a34e6c1142e31010fbdea6bc23f76f65e7a746f6f4140930bd29dcc8971c5f7add780154420414426ba5400ee9ce5d604a6b18fd87148a29b228736a2872ddc114ec4f3d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7348e81e994d5f3eaf61e9a2e813c86724753e0524564cdf84b12cfd341b72f857cdcdddb3b8d19367c87353ac03479b26af5b9fd037f46eecf2cff2c8bd17ab273a973b0478fe9ff1932ccd91496ad65772fb2443634ef4d99681952f6a96b9a74582598a04e91062dd3d96b9c3305f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95f5011f38aab0cc03a29cf450ce1c0a44cd778c213dc51c075ace5c8672bfa158719fb58e6cfacee56baa1ae0cf696059f1fb48090f15660b9166ea7b3b8c036a895c6d86db48db33a74207fd44c60e586fa01cfaec389f866c2162715bce2533d48ac53d22c39d5d311da46af0d6abe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab9791151c78c9ddce7b7f090b0992944c6ffd86ed3fae0f5cc14e6b86b77d0785bd219e8f6ec108b3d2f1732fcc84b841eb3eec5fa590ac4db38f0dcd8fb646db3934d91b5a0a080fba969e03ffb12dd83418210b71bb82caeb353efe6cb51a74abc25b53e7a203aa3dc4b7d2509cbf1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he634fb2321accc9f918c9550a7681d0fa7da8a8483be58ce3b6a8bd1a54c603cffd5a50adacb93bbf7f2f524a7fdb379894b46a742de7611f0795f9470835668b73eed3c120527c864cf0963d260a7ae7a454567d1a81f68975d53adc65bf91260cd895fc9f8093c9cadddb3ec192003c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdb019ed55f68dd444e7783797dda7949a61743f2ae1d094c7f28f2362e06c391ef4403ed58d369c6faa78b0d46de9e56a4eadad5ea4db06b1fff256196197b7d5b4cb2b1c3cea7ef47ce354d72d7817e0b399e31d1f8e0df92d505b47f46e6df5a9cc51b78dafe38e19dc1f4ab737aa2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a6420b2a747f59332b3c29ee9cc86222aed7a871ae879f69f5479513fa7cd9d40445335e67595d5c0dd4f55e63b46622fe58d42669729814bd5f255d8ac0bae7cbc0c842d573d1d41200d24008e4a117a1e39162a021b2dd474bca0afa9774c72bd344783e6db4972c00a552da6b3998;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4aac3635bc6cab71be129ba85aee54be9092ce8de146741170a1f6382fc9c5177998dd5827162b81552bb7941e4b16b114ad650c80b46721c524e6deb47e462c314abab66be27a1fea2c0d724f8ff8f67b9b8c1f9adab80c723349d22dc69679382665c0ebe8934852300566ec22be044;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56408cad6f4e298f34ab714eee2777710551119299c0e5b025ce117c0d68740849b94c7ce206768396f0ec64dfc71c7ad6ca9b384baf0a988eeac17a8fb893503ad3127e287db026726571cb406afc5ee73e2032dce62ee8cf550c78fe7b246eb0940b7664ea87a63de6edf56f108230d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4418dbd6530ab0bbb41b37ca77ed690a764e9ae9956013c81f0b936d8aa6b951b044966d19b5422871d5364ca62e7f83eca6017f1f97c54e02e8c3a463c0ed617631df8d2a4235761df24dd2416227aeda5b3b2980b7bb4d5c4286432bf4c8363b5b82b489a2819f7edd947dc35c150b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h328f01aded627cff1bb6c2d152a173a59c696894941e202bb71a5057777652a70556ce1f3f22060dc592d55f5f3314c746344dbd74ff842d0bbbe025520c01360be2f7db286978b745fd1e8199342896f3e78bd16eb5f312488edc31425953127ab1c6d3601d3333057ecdab6680d0bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h630a0de97ec19cf26c9b5c21355ca34c9285ab7c5b87354ef07726615bfebca09ee7ed72e4959bcc05b750dde860eeb1d171a3ad3c9552c2daceb9f3a98904a88f3efa745530457fce477b6c1b89509ad4711c62d71a5fc9fc724d5b153549f75cb5421bc6657eeb482669547f0741399;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bf4234ab5ff30b4bfabcf482b3755c3fb640c62610cf049254f7b013bf0aefc585d886f2f33bc9adf47c18257889f5a3178f6041a3784c14ee291610b57edbdf10c8875ca6dd18e70af45fb8fd4db3f8579c54c3e926117960fbd7bd7d3148e343d78e28a4eb8693ec6bf1d58ca35507;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44e47ccc558f99756ebf5666aeb4f3b7e8a223b7a5830cb44449631283f12784114aa09145e51c05ebc545d4122dac67c7c1592bb24ddb046da525a0de9c7c17c636741881fe10e09402f14ff5b7a20e2e3b639bca09f289874cbb38767a3ce34fce762128842821bdaa5ad70538c8f13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9d12569d47a95bdcd4ddba9095fbd6832b92d4dc49f20b86f8c61e54673640544093199c7f7d41e3d7a16b8ef007eb7ecd5ecc6de6108e721b073806d5e6bf8ce3e26030420ab13373ce3a3beb16a8c1773b004b60afffced4555285eb53c11099b5b1bac10320a98bf766f2ed919a77;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdb353dc99f06bbc832773c5cb55200ea74b12f8fbb6e7c8cdc8205054e1434ccfe4e6e8e60323665f1141e6394951789e23d57531a268d922d01074d6fa27ad36af9001e6c4cb767a5508bb5f484d83cb6ed8e35197c4f20fd4cc5c01bf4beb3e9c0218632a6daeec37bfde89e882cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2566336359ec9f6f87ac2f65054597dd21d3fbd413f3840faa084f91f35d9e9856a8b19f78f46a9a55be5a092f63e8f6fac8dcc9e18ded85d12262baa09ebc37a9f32f0da1b2af784b3ff9315e0445f516efcb923a8f26b3805287d54b6b22ad7791350a7c3363dc4cf2abc5d5c28e6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66c86191147da31c99ced3f308c6bd074dae85db00acb10b8b0e6355cdc7566e94cfb5e36532465c3a3eda6bc628ba42950e3f55dca5df9a839f275b49c7fb2bd9734ae2b33592de3266a97ab758ba278046960552836b210a4cb8ad1b3c73d01fd6fce36554530fb13eb4c405027cd6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf89d2b0765e793e6dcbebfc22653584b51eec956585d3d41848a1a92f064bb79ce8d28336f2a902bea40faae1ec4c3a605aa20dc8d4236ff99cdcaa73cf09da941f60554393de4adf57142a35d2449263d4c3800d79e7ba3d1b5e1c6c717affd5b5678ac97d053f38c14b317a593b1e18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72e093095aab27f6d901f715d7e993e742d8b8371135e8fd9342350ac6cd5211fbf4fb25f72b76d061bd60b56b5c90490ebe7dd2370e1715f1a31193cca32fb91d891880eb96284fb2632870c5e5ee2b4cb825fc06559372f3cfcc5a62783b4101dc4355d4fc01be6a8fe3af43a7c598d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h309d74703e837e479339c0aec459f0811006a433c9ff072a52e4be3b17ee1f28668e184f62d05ed3e672db32f1d7cb04c50a61e19daffed46246066d8e68a0fd52cf2e8a2b1455e45dec517bcab5d380261efb686b1e72f2e9c9c7684abb00937125bf0d3b80d92677b463a03d3c16bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7718372bef325538884aee29327ce33dd1b829c01fa68c0d8dc346ab30d053b74f6c142462f47409697431b4bed58f6af4575e8e732fbf3d7c2c2ed10a32346ed3eb56c40aa89062eac6914f60dfdbce09350476bda4ea495f8516537ae010dfd6577100b245ba77889b38da67aa5c53b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9165df4dd8ec007ba61bf69aae9b0bbe776b370b8161f5d47f2d6d7ef5131df8828914cce97038587c550cdad988c3facd5ef147eefba9e68b342595931e97edbf9c46ac31f9740a8b6dd08897771b59792933c92178e4ea4a5ed60ffbb6471519b105f11b9d11a4ff9c68c06be0fa84c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d13532522638b8b6ef0ce11fd9b5746863e69dd16a784444301bce559439d9dcf3f79356252151e3104540b0cc670a4b7600283c8c10816312f825dd7c1b27955f34f669aa849012735555d897769a00749c33a3c44ca3c9a320a129ae0ad0f4e8520588c558a17bf2a7c329739ec78e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1b19e22f7af8668bc47a2508b9c83e25e1bec4c26bf8d9ec48f77ffcde38008bb5e0ed6bc33ceab642dc94d2cd254f9c9408abb982c5873db50124fd403484678e37c0d8cf212adf5c45a9b16ba268d7f7fa059af43478078772d49d3b56437225332cfc81825e0cf0d9165ee43ffbce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb17b05d19165a1b082cbe14a9f006c7815e02ecc24cbe5ac309634bd9f6b4c9dfd485eaf9f09e8a76f17440637f91df54786fcec783cee689681a6676782fe0d087964733b6427f1199ec1d6a95e470be89fbeb05024d682efd223afd1b88412a743a7d873ba02b036b71a9632595f533;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he486935fb9834a0ad0bd0f74cc0c3ee8a8b838cec420e14428018ab1ff7c03ac37129464a724f95b1077940e05354f9de7f0d2454e5a61e4fca9dc9ffbbdb6e30650d48f9067a3af98e9eade8d3630b4513c3a319f287d8a14d012eb23502d5f1f70e4c021025c2da845526d595fea8aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2f2a1325ec29fe0f42b215963d51e1f4f9e74c6f93604e49b461f9d5bec8c7067fcab749e801a8c95d5a824ce3b473da12b4fce45d512d93f428148ed1938aaf637a2da3d7e6e54200630539a8588b642e646e29309b33ae0d2bb7c65e9605341530220279250f5d74ab791f6fd04635;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d4366c4f689694b3a122c095430989e4a44b71ae7b596aeec7427f9dcde46c154f526a1eba79b545bab174f2a6075690655901ff35867b818fca85ef4cc04d3fd29672d6b9931061dbab213377d3ac2f0ccc27b383cad80976e9ab794d5c78b8733f011420c0c7b38147762b7e584d94;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e972df4786421200fc3ec819e543337fd9f2a21442b161205d2efbc1a5520c22343fb8b73358e79c9c66c8f6a1f6160ab58ecd9bbb871ff53584527678da0c47608164a24ba61f15d7911a38f83e980ec9163c2a917904026d5441a3f3b710f15ded2a5b63c1ab75c7e0974db5446d02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7da790b5dff95e28fd62ae0fc4b2152de7fe8cae8a06597bb8eac56cd5d022d083ecc47749002a156e7d43449d645b92a46db1ee3766f98bbd9c23a1bc49f0d7905f4bf4c7de224cdbc78de930b9ce6155cd4e5109223fd17ac43806261d6c5128d8127f30e8581557b52f9d2d834e36f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4077673693cc757a0b2249b3a1e0eb3a75221a58376786c9af24e42293bf2692f1812daadc4c2ff21edf736dccfe27cbf58a17ba6a259e784b57cd19b513a439751d5c4d71b3eb5b1996d49776276131aa06e227144046fe1a36ca605ca24f0cb8682420c6e02a76a724670fcda24fdb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9194bc8102ad25b65b82490c5b52fc80fde1b4ed3429b9246266b65c944eb89ca9ea4d911d56d3c7adb1c8d7d36af17d1cec37c61e6d61847caa985add3532825580cbc070f1011bd31bf46ea31c7796c46f1409d7cc58ac4d2fffdad7102b5de1771be5dc69c0cc02fdcb387e95eae4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8416382b5df92e038286eaa777c9958da5a906a58c16358b6588fcc671026b8b719438ffd344ccf22e979f28544f6e9ada6fa12292e9ce04a90cb3e334497c994ab9792143b15cef9fda25d1f65163f21708e2d8d9fe322d47506921ead3b2ba53624bd78cb8b8def0b70c09b9182d7b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c6fd70c68929dc73d75b63126cdfd974db814799365c22a6e931fed2c142f76dd286ba887fdffccbbd05b0ae72f3f6636cf5b64dd78a7f9d1a6d1a3cc9a7a0ea4541e8ebe4e83060fa170f948fdd5a237f7f91ce7e1c42288a3dbb91b6264ce9c9d9a0dd7da0733b96c39da23832a538;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1aa55f965dde847ddd1d8409dd8cd26fe6d3f6d07bb0fe414221517a0d2bf49621e5dd47f3890bf148b84e618fc77b85c77016ee21834774ef9b2868cc7278838aae22fd694981e3778316bb881feb28999a4329403d416786add8e8f974af0920a9933553d8fef16aa78ef67bbe4accf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19390ec378248a762ff7d1dfe7f54f4eb54e286b99276a4726157e35e1d1133858dceebd0b0d9325ce6ee3d1bc3fc071ea92c60422b0975cb50b6a394d7fbdc745e361e00fbba8041884902bf2f887971de43995d4509e2ec588b209c6788417b3016bf014ec04d4f24cf09da0578b390;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb168204005fd5077778c9babe65b311a987b49354c3e86411477d637918aee8a2edfc38254f2d4a82f55ef0ed8bba7663df452cc9bdf9a2ae012a418b2b0ee21bf49f3d47c5b2e48898d15dc2dd34dfa61efa2f15d722f6f1448cc8685f5020f05218c654e3415120760c8c2cf5bf2bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h610c9438fa3331337e468365328be365b15a138b32f2d0eaff35d31d909390dde4dc242656dc238b8635afb3d22bfa936b97299812cbb7fa47015eded32434c2ebfb24733d652aa40e6c59289f7cd4b37f22ffdfd21bb7d84cc4b2352b435386e3245ecb69a9e5baf414c7bdf33a9b3b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf3377247c3852be15112d759b0313c77921bd24c23657d2072b852feb2f60831ce97e6dae5f409726bf306bb876b733483d5d66b0fbbc4ef6af96d12a1d245e55ee3f232df90f0a1a44c080a41a7fc9e0d08d9e67b5fd8969f796a79d7edd963728c1778223c7194e859f7535a5b06ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he02fb99d4e0965c5b33be930e99f8ee3b8ae0caa8785bf2c96a70d9c1b9bdd7dac0a8b0cf2030653a546bf65553fcbb9adc4ec4156aecce79450855ed30b171cf0e85276821d6d7aa715f868c4fdee202ffaafb59adc27353eeb9b6637986090d4cb35ed3bf7ed3bd5ac94ba4a0966980;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8a6535bc65778f8b1104b9abd3062f7c39135ecef3f112bf3fc31b5b1613e95f409f87e9efba5578d27634d493a2af404ed250f77535f4469f4c74b27d9e3ad193e859ba2f8da168220da2ebf7805367dbb268aaf2d3392378d17743891bba9fd1a0f51d79129887057db1d3b16c9430;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8d0de0567941ee3f1424de02635e5e2e8dbb55791234a98953de9c1f220afe8bbf5402f27cfd532b67df3baa5c3e64cd96688266a2f910ba64cebce7e8e592fddfd5f9b4b4a065bfd34f6d8c261c359c811bd9e85696b0dfb82a256c308479f496f628ad154bc2db828d8924c3f6afd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32e772165941e0262e37272d3dd74f86aac624c0db3b119325bccf323b2dff60496beb43b09ba75111950b08982f5f95c93fdd5d594a00eb68e60468bf8fdefa8fe6b2814c3088d4c83441a26ef6f4e4cbb0e5779a0d5a3c0415331a3e88772be3ed71f4b271b017c4dd300e32d1e7f56;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h355ec66a9387642571183dc5453e4e9cbe635e346a5cb64fd1f12982166870837b9ca2069dedc92d9a3336990fa2b8d4244e04e4b61d6654b97119b6c60050c4bb1f52405f67be425c19de74fe89f0225b50141c793de1b88c7268b2ca291d0c017fe4aa222fff8948db51273109ce7cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacc4b5218f4562e440e39ba6c9e04b2c2f476c398f69d046482116ff1c31a1f0447ae7a395fa59b82efb2bc31dd533aa2fa7f9e6b2e63e24e6a02cb7a991119f78b465ee8eb4a53b6d76330fb21535d4eef1ee8b5c3c706bee4d2e8359faed264201b902466f49e70026cb8176ced1c4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9787d91b5254d456208965ff31814dd6f4e975a6635d46d4c6e901e1de2ea2cb02a9dcc8b1e0a4844699e041a839d7ed626829dc60be10690c3f388b329ec13345a4d3e6277ba622aaaffb8b06034be580eb5363712e39c068fe702ccc8e5d75dbb35035757734c779cd4ae5ce337f96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc92708c55e0fb625e37e69cd123e5867a059e2053ea4d79de7d97c96bf016ebca77e6b093d10e5fb5505d425f8ec189290d000135ec1954d22036f0807d902dd07dccf31864db590454148c9037afdb9b38bfbcb47024f1300b242b15982aef14e80e47c030fe55ab45c5ea8ccae596d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90c06ba11f95ccd42b6c56eefddbb56b144b29a89e2b41d37192d68a895194e9a4ff469dad10c49d781b2ccb85e6b92dd6869820a9a1ac1e0ba8c2e5093bb06d3f2630e965cd10e9038bedfe6586c1b28e4748a50ae901f9173e2ffbc055668e7e375fa721dd1fe567b86be57a346fc94;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a1f6487e9183161db65e15314aff004001e4539365caa79d43e4ec7a52867730caaa4f26f831d8db6e72aca0ac73b48c3aa48ec26637e04ef5ca058275c8e1802740ee40539cac2488b6fb87e10f80d54c0589b4556c2020f526324c1741af96ae6f67a58e459f25d5bf407589fa2897;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1b91cdb9fc6f80c08b6a7cec69612f509a3ea859d155c9224d9c55fe7fba02c6932af803770abbaf1429408ab0d65917e3e973068808fdcb8d7f4805c7e5cc44cd4ae94031906ef1a38428f49090654db948ebe7230f68d8c4be3f44b4254f06cc5ad2c5fe84c9d64fd6d4de3dfd6b4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h539263d2dbdbb8b2b1a7ca6ef7612be3d740ff4d0fc6deb8462dc488915d73815f889fdb3e39b122235253e87e415f5c84fac580de1754196fc9887a0e9d08858e8af86b59fe84ac5540ac086e0afb557a30eba26e293500aee03c7d77ce791faa83f495f9b4c06c4f4d4753123de14e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51f9a3a5c8f3fd08082678bf1cf40af8c49b8a6e7c914f04dd7dbb167d6868b1c8f468d74388641b819e2dc1f28b1623a3fb6d806029a889b3cb02f65875febe735d1e4e314d996dd0ef9dd8b4c1e37e7cc012526cb41375892d16880eccba7d8d15a1fd77e0190a55cf5a63a2f55ba21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2d7dd71440bac6cfe73ec8546592490d481fe6654ea86209bd67d8f57cb54158a3031a91019d0df7238dfc1ce5a139cad5f49daade6c9c6e779c4350c90a7473fd6ebd76e6f4776f8a181f35c41fa794dfbb992d01a5b68b06834fca3124a56b5fafe63fbd858dc77d02401704d1e5fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb5c1173797058af79802065f5cf0d4fb4353fb17c103e906929a6eea466552c9358e4db9c4cdf64514c615b68390362571aea451122df7e1c890460a6e924ef51c7a0e08891ac49867891b34ec4d2c93ef23db4c19c1dc58881bd2d6bd1c2fecd4a2661dbe5f78d92058ad7ef9fb91a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4923aa2d1580873f35a44db5c7865c613dbaf0f82d5e3265148039ecae16395844bcf8c1e34ac8dab2a6f84d3ed06f99cf9d2556464323b1329220d22fbe09681946ac44fee7821d5cf8182ed75583330fb8aee815520947a14e17d789a06d0ed00eb3cca4f830821bc8f8daeec95c185;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb799d75b380b3acb34ce0640baa42d4bb71199df9505e97cad71a53843d6a423956f2fd1979c5fa7e5b4971c0da872e8f50833fb6a023a1b44d545b8559ae16f60cd56d3f88d05cb4c92bbc918de616033fcd5400efc1442f9507c107179304cd0ccc1e245a83689d657cad383049238e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a1269fd38f38adfb51123928a02a73795499708c532b5e8ba5e24b584a33b290f02c3686cccf141ff4543605469f45f9ee1541567d36a9c00b54cf832746ef6e15ba5b0943d49ddb33b31f5a934557a32e6635a0fdaa71c761ae2ea5d3d84746db6e2d47ab7f14046004b152190f27b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec2c0ec65c443249059093f7964b608c4bb52ac9a3f3c756354dfd3b898db31707f9d2d25cae3eb1020825b183d4b8fb9bf48cfbd2e5014b8708b9ba23af646ecd9f49461538c3ba6a0e4f288b5bc4ebd3e45741e8b62f7e3ff19e92dea68ba1cef39d5c96a37bd8fdf923126542b4d7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h496a3c7dad6a9d790ece4588a4a09db7af54ca460e626df93cff2e6adddaa377b253aebdf4148f35c7d07445ee1275cd5c991ac30fb0273b3a45740b644708612395050e7da5fd52f4516ab617a6f163e634135e7bd44053d2cf0a0d5fc5d17a66d86e1ff2205eb093d537671a170e258;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hede69f67de0a42cf84f829887c36ec9a5a95c3856ba784ff908a91866d036ed589f98e92601674bd6a34bba75ebfea8943e2d6b354e2cf983c4fd606867ac2c20402f7b22c1e82c31ccc02f72683010205b215af1e075ebf15f65966660b85b91c8e5db4ca37fdef52000fc1a36b11006;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94e9e01fc303906bda0f28b83e4376bfbbade8cc9fad34aae075cf51418804a7e447a2618eb47f2ec2593eeda6bdeaf020b99de5adda304ec7f7dbfe3f4116f6559e56069f214373daa3018af18093c147b90550491a4597541756bad6807fe359f7a7f184a771e4cf476437d3c7b482d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a73e7caa0a46dd626f0ed520b351357e16659afc3a10f29dcdc56ad788eb40107faf0a0eb92fca89edd6d6a5f605b4248abdfa5686ad53705d2a9a2896d24437a51b23220eb3ad2f3a3546dd58faa4a08a8f97dc8534bfd171ea5e0b6750165c8f9eced53b8e8044331ac2c18dbc7ecf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e5bb17f333b251f478ecaa17561a010622e5ba697da434816cc158e9536d6bb2e20ca770589e846ffd4ed23eca3075a865b036bbff7c4296762fb3404f21ffafca2771151320fe355bf15b0de95f59b661c97bca359a75c82d25db13099cd00034973305c6775fb43c3575c9bd77225e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bf7cc6cb0125d54fac1c5bab79c820705574528cf0819494d5bd930b48f7787f804a6a18b8659140297e5b4771b900300a42aa6a4ad00eb6bf212be3bf388fa94e9151b62d50a6b8bb66789d7b3960837406eed55f773096ab39a7e9cf3041f5fbb8649d0ca529a9c71889ec3c32f96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42bb8f6fd94b92ff35e61ed17f3261c0c61691f235a01186f94b166314de9d4a163522d33f08a332d03eea1f0fdc44f72c4178715b586ee4992bfba20121f165ed75841ae175cae477bdc9404beb34e3f28a1fa342ccebee6c4ceca981559525d5cea823c5a7df0ea30652d507e96a6ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34ecfe67fdfa0a8d53867b7cd47753cec57b279c114072810732d653337288da40e1a3408e807bf303bebd42b6d5b4c9fce85c04fef59381dd65fdf17617e8732dba6a0c374679acbe8016977069b1fd94be86dc882894a93531b0e57ae858156689a1e3ac32d5a3bfb0028720040c075;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6cf71722e76304e1d241931e5f497e78e3eb321ac741ae36a41fd967572ef7f0cfb25eef8612c674d6bdb0d511e46308d98b7169ab0e779689e5bc8cb8a8d9559e1de34564d22512caae40d943efe1b2043715db66451100b4e35308a3c645142244d42c899baa51189c05ba2cc0dd7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9938067039121cf3e97b5a4e6e653ba81338233dec2512b068048afd390ac771f91b7f62c64dc51f39b9b3f57dd365b20769a5a8e8608cae51452a8bc9a395bb0eff439758ed7d9d7b78250f648e2edb126803e1103e12d902d73360241adf356dc593ab7982484ff0a183b42c4a67eef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fa645a13d5d3bac479ce00fa1c705c065916392a2c93da8015fbdaf57c7c49f7da658903a0cdb95fbaab50c2b0fac135c266f6b3d2bb0ea784af0247805c8dc8eccb4a3d0135b6ebf9f95eab1669de319dd5f1d4418ba3282d41371d03a9e8930b29c54933bd5279f01466c46690958d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb19cc64a7d2e308dc1e6b4e85ed1544adc0286d564e340e95f2925f1c91dce9c5d498f03ac930bf69b9cd5c5b765ffa6b77c11d3f6b64401d2dd17b11b1a4bb257efacf553235abb65b2a6424962677cf0b41e5d281170325ec86aea886963ad316d11095c8c5d0b6206f0aadddb0848b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2b369c29c7a82ece887f8725011603d9f1817c04bcae38f8d5363b9b56b30a37cf380a2a6b87150dfc4aa06e19d06a07167a1db8be609854df6c55ec22a5a20e970126f3d95cbc4ae4583f03e148446c9b334404716afaf43701342ad05ec6c50a4381cbbd3a38edf6f9f5f32c7bb11e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h557c34ad9d07ce3dad590263c51b93ca70bf7fe72706196f054b8a622316ace4a1e9a21351584a24b925edf4088f541356e6d4e8b4d4adf136e81f9f1c34e5778c0d5e1a44fecd9f3591590fbd8826450e7cab6c1e027d1e053dc1302510b8ee1f80e2852409fefb083d34a9eb76cb609;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfec8aafe5a405235c3a81d9aa19a285d6df805888c06756a17c307108bff87c05dc0ff991857c70efdaa9a5b900e3eb9e56e7f624c096202c21cc534ac5944812a36b11ab1ab4c2e59411ca4ad81a3872ba17503ce37d581018def742866da4dab5428626c57d9949ba9730ba80644b00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d99ccf078723dfd8d82360efe41e6cb96ea89f48edfbe302d707628d92ba4bd65d1380145b3db01c4a6b4827c6f9534c71cfcb4a3057b40ff81a3e07271168e530a3e5b48096203309b5d4ecdd3f7680d4c9dd2c5289c4a3865c0f9b1e65e4c5b3b4d856d7aafd12043491f38f522d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fe08d6b2270b340babb10bc38e130dbf8fb6e8cb43f0f964e3b3994eb46f3fa4280a5cac2916bd32139f8d8c12669f9ff1c96a010fe6d861eba1013e46d414f7f4633ad3c4b40f5a1c406dadbe70891e94e19cb1aeea6d7b4b0eab0fa9d8360bbd05a5777e08acbf2c79b5a83384795b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7135d7770321b57a5a46a12fb5555d2bc908231967ba5655be3ebaf7004c35dfb07e77d522a024d3c2647bf9f0ee14319bc747e7e012e7b5b49a5d87f20ecabfd69e34db3d8a1b3a45a37ed6078f1acdb19cc1ce0565878696d60a5f0847a0106debf9b66d977550476c8add82f2feeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6a46b9b01de2eb57a5e65d270c5801d30a09ad6b6a17086e069e8b925acaab2db9ba1216e6413a0518a84468ff2d1eef4fcbf6d22663e0523c70488f7fac8846258b7442e65f50f48d0ace3c6f37d0dcbe330154b215b47b1f50d4361ddbd6a8adca9d05ce39a967cb28aad63838436d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea6dbb985a07c39d8c5d2390058f1381a00f3115bcf22dbc03b2876a16d04a605abdbb4307685c04483c9a91a8ba3d736b596385d7cf3977e1be467b109a579deb10e9b35d1cc1eb847f7404610d1c6fb8fb6315e0f0a855bb2340e23b0724c18968937c1fb840b4e4d88a15edd1d056c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf35d4e10ff8e8a49726feaf064c18a4a11312c99ff219efe977bae3d39dac27d2f4af18ddb3d205002281d77e7b5e29be01121ed1b1273e340e6e746c162f069b839299f2c2de573ce0485a8ff21fc33c77574d8b7f1c25447f33031170ed9ee12813d9b0b7be64cf72b6e9764ab2f939;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb0e739658a9be929008f87bf33ffe65bdfe50904b57a2b3c35a0f793d890959ff743d7468a2aff5a3e2bad07120a50ab2d269c32be5a1089f6b13af0fa59ef91b38fade6ea9e691ffe8875f3fcf92c86098d00e9228c256d5d3dd806b50ae71e10b1cce1eb2c826b6be258f1314e7219;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85b0e873b29ab247bfc5e72d46ea38a93132af39c8ec666b213b26255f3293daf34f8d2e0e3dcace832ae01221f6bded119c261c234f9a47306beb354fc5eca07b42e5d630a100a1d733e858c56fd3f5aacc6d7ed5fc4c73256c2eedd6528b321470313c69957f4f9fce0924cce3cc92b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8273c312f2f2576213f6d9e36cedaaa9f2cc5867d200fb76203c08c9e5278dd9423b128540b5b8f5735849fc944d82edf6c1202aa7c9d585df42fbe561925d5eb7a82c0c180aa8adee3d4e24f6401dd2a4f285d76b7a13ba4a5837573f39fc02024e6c9fcafeea2379b4078d020a96eee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e2d9da731c0c8a89aa57f206d71d5cf987eabc8f2bde02bb1876b683eef515c5d2356905bf36fab2b3062f6b4f74697a8850efe44747ed9b11dc49f9770d47c5f202f6aab95298f0aebce813329dfd362d32eb2eeede192f95ec0aefd8719ceca9ef2dfeef7f21175b25d222a04fcafe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb23714a4f86a516cc174e4c209230c6ca84d5bc9fc3890b989186419b228ea4abe87caa8209f50d7402436911cf0c6e55d3bc7e86563d1fd6a404c879cfad850b81bfc4d75efba0415a28436d9343f3c79c106fd34b95a685a20b4d799e421834dcb0b0cca8cbe2de6fcf0de17ae3149;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94015cc1b1a68868c8a03449027afda28239a1b4527f5ab9a9f055dfd5922015cc551441ae8c9808df41bcd687fc73a593ce10e72bb6f2c053adaf931ab6d2338279957df0caf709fe759576fe22a249640dd7ae25a54ee684a2fc5022c4fb5de515e116000af98aa566e4ba69ad49936;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b2143b218cb797b9f4cc8019048b86cb85840cb291e129a011a987925673fd8cb28e3e79691d87d3ed036e0073cfffdf554b71ed68ced6ab0fbcf513c31905557a90b296ec5e69edb034daf056f62fd27c9693ae8aeece31e5828dd0b37393942a79304289a27e6ac498f8da7d7546dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1efdefd378b0bd4ef26fbfeea3bd557b20a68b70ae0c6f840987a05c4023594482ee64f46401b50e147a962f3f38ddd386337e7d572f5f16fac981b1268880a00ef5538e3d9d5193b5f255c0eccf32535ed1d649da09dc1b845e3acb96be82913f65216bba72c553f8b0baa58400e3c2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5b0ec5d5abe94c4b451ae33b8fa604b12d17bfbd924c21376b27bdd627c22ce93c3e1623e73d5d2b1411740ae54740f3bd7f985fa798781af5446b72c7a9d25425aaf67d4da1b94e37a5d3da4454ce89fa072db2420eb2a4334fb4d5c3784f43ebbc239067b3c40b68a4eb9f5b7d57c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21ff3732896652f574558fbd2ab320fda9678e0eaa1d5c3af2cdf10de1c1f619703bf9eb75605f1d182e007f88fb53ad01fec2bddd0b3cac0561e4b5972d706c84ad0fc769d1afecd35306df28dade77ccf07eda91ce0dac4096e235d28a1b6e0410e57ca47bf52429abb0bc1e6457db4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd593b08ff329d9faef5540351f7bbd3e29a32fd99cc075ac6ab8ed7802ee3c4f169f7f8197d50c3b6f324dffb3ec544904e0dc195dd8e77ffced7497df0a7354a2fbccf330b4421afe20d69fb921e98733a187b4b167c423fb026e5a0fd47bedd3000961956332c6532702e9fba28f9bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbe8c256fe8101018455a85142c3c4ca3c5803d1e5e8edae3512b7f81786b7bec35a96495be01cd63028962a33541ed364eff08a87750e7383826cb55cc7f92e85e63c77a0b12901e2b0bd8b8c2007748e9b318dd5b39b191dd23560525c9ac1e5e7afd8c0ccdfdb74b1412e419ab845a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h567e1b3f509281a257a1d23737e7df8c45b8d04cdc59891f286e2bf737f88207ea27c3fbf7a4a5eef28d59bd709a0986bdbb28c041eb7a69175e88318043896ceb44540a01851e03641c663309030e54be9348b2260831fe333ebf95ffd8c5f0ea13d5cbdbe7c19f87a16ad3c7da4e434;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdc35ccb3c57e5cae929351d7e9ea853594aa496e0df656c439dbf3b79713574c2763d07f815155b89072f3cde8c4fd9549ae404caaec09a68e6c4feb074cb4db2868f43142f26e93913f1bc7e39188168fbc5c8ca7c6e2008ee33ed93e896e8363fcff01755991550f4e673cfe2cc829;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h244b46ac5052164f9a8ec625e95f6f21502dfb93e891342b3077341f39b56671e6474a186f3647cff042071d711eb30f8b8fa93514d34a791d1a169b49f6b70b0cc1df5240f0af05cdd16e1ffbcfb0cd1461ba5571e8daa8e6d6e02bd613304f21de982847c5f81ba20f89bf2da9a985a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e0e62e671c5853dd7f21b1785aad11c0b7518d772ba350e8f25e347852a2dd3076a531ba38e199ea5bf5fb5c2c87ce0b5faea6f6cd966b1391637f7673068379763649acc1c02ea11908094357aadede62a87b8059b311d3f49a1060a621d2194ddecb1997021ece99b844058fc3e809;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb418ede74f9400e6bb22c83c47cff6776a8e26e45b728ee7e9ff0216ed13a0e9bfc73f6e537bab8af08005c074487fddb22ffe7058888e5dcf5b088cc977ab6b8cc66c79747f256547e87f9befd65fe0d517738121e5deb71dd61da7a1c96d59700a331f4d77c12368abe5d1ba5448c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14d7dba1cd1bd2bb61c8b88e65817af062752115bdc023d001068fa27b6b1db537b2002963fb9ec0ee4621186d44733181b586da0d164f477c9b1d1995b90fff30f0a54a49633c0a394e3bf04ad49063307c75c0a826abbe6cee6031c2e590a701bba6683a640b744369d3c82134c1cde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d79ff893e10e03dc65c06249d66a3844afd33967315ddcfb9cc199ecef6a17f9d0856de96e9436d1b67ee47694c266658a0d8385f76e4e1d7c1ad9f7e02bef099db645924c11206a8b1aae62a6bd7e329261dde00f4a309751360cad4e4597004f2e62ae329d50c44ec8be1c0c8c0017;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d670c1adeda9ea4c3ce713f4c9d0b84b90e62ee3b3d481e8febf822361d64b132c05557517d55d9318ff2de443e6b9e2d24ace562ff6cd6c739faee8de0336ffa1103426aa9bd38ba553229b0e883371a16759cb6f8f3e6fe8f6781257dce1f52b9cbec0301bc27d37d6423c666f6603;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e80db2de54e44900309841c4dc79ea0b5b09c5408c89c3abf2b8f2d0225ebbf61d90c5df1ddb5a45924504ac6ba9cd34f5f50dc9a3c4bb3fd3078b160c3bbd5ed5e26a0bf8d0a5998dd62a66ee8a3e3d27d712544f620e20a0c96db8363ea66cb140fda710f0ecc3da33d36ee7c8d0f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99ac803844474941b623d4185feef52e090e9c16bdd793e00cf7afc7f2969a2420b9969e3bb8be04e5a38959210ae9804a8e513865b7047fa938e7f7af837080509ae046db237429ba09bdb2fa4a524a5dd95f9844954e05b26e35651d41647dfa8c5604195993919609ac70763309194;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75126fc2d2a59cf8dd7936eab5fdd7667302c300a8cbb4486de8a68cc7be79737dcbe27ba54e607f0aac4ee764d28b376258cbe6054138d0ec1c798c0a27e22ef9c0c7861be1bc5f6250c67761e5c446ff3dc2235418f8df31502b5709809e08748e36aa0f7fb4e4fd85d6a9a6690b923;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5763bd97cbc049ae007f8a3c94b8acac0a453a308f73e65dd835a05a579a30938da48aefcd3d340c306faf79adfea57b88178f9dc2cca8df27fb2511ed655b934ad6a1bb1bd6dcc0cc5aaa6715477e1c869365282c174553dbabe038ac67078b58daa7ac372fbdb5e2a2bd3be900067a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h374e6020738e631b7addd9269f30ef86269b518203c1745b8e8a432a7a71177c61755154645d492d92fc93a94d95c3d6b839f8c94f514b5a5dcb2f123c3cda111d89ec9189edfca4ca06892e4e2fe0f97e6f4050db85e1baf4da99dfe263b246e29d3710dfb41921672046ba4707ef022;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b9a739a28ef9e9f0f895f7e64fbea46acddee76c50b4d17d17ed09adc0c02854f451dbd1c434da6bd9999dc9c35a4034f1c8b70703475a2ea9902d52c464dac2466a29a89373ef30585dabe5fc788d11f0e7fa20212e4a8fb307b7a0f8d285ee1aaebc5d7437b83c6bd9ad1bdf3c9ac2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h352cd9c0e252b84871a8a0a28244c2c9a23e36e4239797d591d17065681f2eeafb7639da96d9a19d4aa37172244ec670f033a3828b4de7ac5f5abfa3a445796d526e8eb12f9762091e486258f436a33c4970d94a2a25eecacb16473bad9b8c0aa322fd565bb7683b1ce7ab7f325d37727;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4eb199f1cf04153232fa513696dec874e9ba0555e2aa006e7684f977bae80819805bbc3dd36b43c1fc983cf3a05ba1e62003557e8f11dbb37619f1207d3d5c718cfefcb4002b609672574376331320e5325bb299556f26dd7bb5bc52e45987af9975264e79d792cb6a988dbabbfec2ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccdb1b234b4cb3222567bf49dff48c30730924b709d2be31ed90fb97dff13882dd1a640ee0d9bf8a000dd90e0faa9c7b02a35771af77ebf157e31d73b1a46640e0dd925982aed0ebfcbc1336d2c876eb579b9771a2cee0fb3a266205b64ea02c1b3ad32bb1f274ace76ee1eb9caf27245;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49c4cdc1b4418a658bd377ffb0c44c044e8cabb1e98a45954ebe4ef095424913f37b1f94f03ed90c6f0ae8fbd98575c0796c3a4a26ca9d3fbb155c2a33c24f797c07466ece7a115117773d007513e4ca1023d6d02bf3a5ae54921e96e1eddac62cff55370fa6c987e3c209649ff673314;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h658ca08abe848d7ee4b817fe98121980272cc66a741859161be3d3121b46fff2118f1aec10fb86d4da77c795311f713283246ff0c491e3511d19af61bfeec0cc04df88100d7ea35ba10deef8736607888b621437d4ef2cafe94a6cb83b28e937f0b5da625c9784fc356af562a0b2dbb73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b68aa47cd599c810a346398c7243f654e5a0b72398c236c3e70d507fc343b75cc5e55f2930692e1f958fb4a92527de615c237f31a80365727969e27651b7a61c673261955290116918c08014ff72590e180f57e69a709720d93d459edc5fb4a6584269e689aa162701d862905f56aa71;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4797902c1f4d5eeeb3500a70766c3810c6dcea9bc8b1caec963747ed05259aa967f12afb3113dffbcde59c30fb521d180560fd9803edd0f13cf57237a5a10da4f2bf0c1bc14f24051606f06461668c42cf1fa441d8e519c75acb6c9b2a368ccaee428fa919acf6b012657316a878f78c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc534ffe907bdb187720e2bacd33a0b54bade6b419aeb8e51e0dcda07ba9790b77a2ed35a385dfc86b23d066f1aef6cdc2d64a28d910a2f9b65d8e8f4bbcabd5fdc7cef75f3898ba6385021a252b643dfd266d8506bf2c03d9af4d9e2953410acc2c7179a4dd3bce9ce0ac28ba01e0e66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6de7d0fb1e829dda761e5fae8b6cf32192932fa0ae913ef7ba2e7e6e80edac8a610280eb0578f381c22768e9c41478042bb180cbe369f4fce947c1bdefbee662f77ae882cc79c7f1bee9af319b5744eace14a526070f2556549bf640b11c5662da5d4b7378e6870210f84510e0f5b55f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3740ac7b8858a7221b9062d1afcf0eaf247fb338c885c1833c1ce371d2f8fce5ffb0433964707d600f092eec57ba2b2a2fa6dcd6d998f72f7c7ecbf17c3e6d27860a0b81239787761b4679445cbdd7f511c349454ad247a44b5c15c164d6a17a807eee5e55c4eb3115753640272ddbd75;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3def59f8e175eabd906c650c4e01d3a33dcdbb335ffbf2f1945bb91923abf1888cd5942f939825a4baa903e28a1f5b1d6a9ec9a0b7fe286a1cd544b1229ab6effaabd6ca39be8d19c067bc8ed7445c0464084647379a55ba8c2f2557442b298f79e0d00f6ce05191fd755c3e0c44ebeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf592b820fb6d8ab512454ebc8850d70703fb121daf053110f579f022c7a1762692f01c677d3ccf675cb0d4797eeae23e10fc09863d95486bc6385a7108252a9e1682a323ea586b750a97a22a60ea1a87666810e590d98f7e6c321d5264fc936a2151c2a6f03c64192ebd40367b123e46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41daca49149608c6127c8ba00199f8f156a768400cb02951ad79e72b79b874b6fd26295dc34cbc859289b5f49cf634295d4ee699582841db9bbcf831c3352b0395b8e285bcad37fdfb94de52ef88cc914232de8b1986fb0b7230fb80d0591044306644a27610117a28752c477b056afbf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab744dd9907e4f08be5a4b48af6bd501b3cb3adb9374bee94d787e4a4a9ca4c1ffd37e4c77618dcca3b58c880a6728a8c7f09b7c5c6db801679aa35d204f9e6fcb689736edebbff3a6d2dd2d0999c1ee2d90d30872a8f5b43dfee41583a3fc4d6bf7aa3ce23e503789e41739f6ba97cbb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57683ec4113cf08c74ae3ba1f2d92a3c825d566f0f054c15785c58ce2dce74a0f4f908c1217159b6b59011db6cad8d5376f44033330550bd31e4e74109db537a1cf764468c97fb1ca5ef106c3a386b7ba1dcffbc4b455d38d12c1c85dd3ef4afd868fad2899159002b767cc0c4b3d45d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40806030228a0be9306a19650b1fd3ca712539295c435643fd41fe36592f71be26b2b63ed0e8f4f2d2de6d19d5fe8d41f75a6ab498a4cf4a6e89ce55a79e508f31db25e4014c00ae404fc5a5d2d0542bd7f85386a1a1f9d10189a273e78d4c27a565cf6100f5deb07d4828b9143b0b856;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84e5261819e9b5a08c03c04136a543626099349f93debc24de1a9d959d45ab9d2c4e7f8568c031a372797d86399140db8d65b77568f875da54edd4680a7948fa3aae8fd33d51e5b9257db7415071bc630b5b2ec7a5daedb62f334ea85fe00d8e2ca80e4bbf10ac6a0ac4726b2a029ed22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ccf8229dda8a21290072a282d016add79e20dbf221cb8f03fb45a9878bcfd230a0379a9f8301c0e5acf8332d1fe944310df8a89e123f213cf6c64d2120135ef6364cba14e898a8736d1a2daa79ff115163ab3348ae02dc7ca4335468608429f9e2c8a428b45a597ff69f0ca1b4cbc0b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha781e7b6f662a34df8dbfac404518a4c177962c1f4e2d4493f5f8c554f46b07f5c29da7c47c7b7a2c66a45c28eb6215163ed1cee7bb583545e09265fb69990a5f02905885b3e472bb1a7fe7a36c1a922a7b9a7e94d1be7284385094130fdc87db026806173b9b8c444ece8ba3e2e637f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he167601984afff492e2263d6f000e83697a6b9ba5eb859ea7cf51e456906c206b67f51aff9f376595f9c9d7644235473470675b4c4c48f53ba667322d9b7a3e7d3ef211d826c38926fb3add4c7a8ca73e292e0a6bff7bd7001644dc59f4ebbe10795a63bfb1f79e6074beea566055ccc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcbbd79226fe4a829a342eaa5c9903799c21efe2769cfd87ce75450ebf036f83bb996c1b70cabf9b803e37982bfaf53524704d9eaf9053827e4166e8b07c33bb6bc37b1b409d1be2cb66095bc4121587a880c859124f50f96ab8a1d5b37bf4e8537a0840b8f8d6a29c91db08216e83588;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22cdbb6e97727b5b9f0e42fc6764c99efb8b936dd82cfa5a61abf571165cadf22183dd71946550a6f9819d7f1bc62a811872dc84379f6fb743e580ac897b7cf6cc4a7126d6332e8ba31ee206ca42fe5c0c830d55b10d1e1298384b80e76604cd827b8eac10dc9be8f5661536ff504b6e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb7b33c86d568365ad4b08c301ea18200c478d7b342fa8224dc1028e29904619070440f43d2c85f31debef910b38ab91ef8c9cec1627012c6131b7537944645749df7a1732b50f986ec5c3e0d1bb90a55c483d28c5c27aa47a64f2425bc3e0a42fb700b9e15bccb6ac5302b2e16413709;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5c4e6ca340801966281b07f49e3218dffe7c054106a9743efa0ff1d874940b637cdc7d93bc00e69f4cd4d428ab6fbee5e9ab77fdc372b3eb0d9285495e041e42f0730d00749dd1d62548a12b0eec4cebff7d277a12f45051471a36f752e9ec4697a273569d2bc62394e909c180876a50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3123bf7c9c81e6667627a94fc61afe9c6b06c7a7fa1be4f5af795d5735d54112f50821aa7c2feba223dd50f0620f014daed4093c8334d58c09e6186f559bb6d49d77829ca3c299bff7fcbd12ed20dfde223d75b01e2a013f2740c8c04e6fef69ffa31836ec773947da1c6cc85fa317629;
        #1
        $finish();
    end
endmodule
