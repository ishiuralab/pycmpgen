module testbench();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6656c88104be4c15f8c1a26bf0afdb44cd41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8d96adcc3fe8e0d25051584d8f860a6d22d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb91252e00724f93b40dc826909e57b5f8771;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf873bffed78c88d27868b1631a1a9ab6ac4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h365a9b4b800d75462f79fb826f20242100c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha88e4ba2d7821bd0a1c86a8946dbacb0da25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33a78142768db8511476e31712c95190ef95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8647e59d2a10eb5659e1492d6fee70e7733a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bbcd2b5fb3d7b23875e5c61fdd641dde2b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf587e3e0c89bfb5f5515c2f8d2c7100ee11d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20a686c1e4bca021e3315df2379e39f2235f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fd8b18044445ffe3546525e4937d98ddf02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2781128cd1394caecf4099efebd82597a08e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28fabe87d520c08868a0ea23708b46b587ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a8af2a4657faa0c7e809ebd1a95872bed26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45ec1d535a635029a01f57661bbd48dc40fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3295b61b99b9610a0a180e7954c7ccd4f96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fe870a35058343f88d9cf44d51edc203142;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7ed55b76e0cd4096cacd7b2b42a03ac1b88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39fbd01eec7f63b5a8b1cc0c069081c86000;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33162938f234b5e9f20d57e24f2ed94bf802;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7896dd510d539805537732b58a7c0b9ac78f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf13c910ededad7b5b87d26f60b737c393b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf898d8ec58a698b9eb4faa631f103aee821a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb54a1fbcafa134352f700de8340e7eb54019;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha81cfa78071ac02dc57bd6a90d1aa8ea044f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b43bf10c83d1918338406a3e896f96757ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74269ac185464942a331874fd7b419accc88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58121476e8e9b7c6591d808057602b09fefa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d871a9d2b7539eccb14b34258f5cbcf5ee8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84eebee32b2e65df4f2197341e3b9187b3a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2a7ed061b02a026a300b26590e718c99bea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4efa1a095a839c6270d1ba12d7ff9420d48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc8b9ea211fc3ad9ce87b88d4cb3e7fedd94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h400c6aedc72cc86bbe595f5a5df138360724;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3589ce749230b7461d57e083da3a93dce982;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcefafdece84417384164b8f5ca31e87e8a42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h140d07c4608b2e64c159f8420a60633a2d3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1644851392ad16f4ced734df64dd5a54b121;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha02241e04e291b1997d022f3ee86569644bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cb566abf55967fe6596d943ae95732bc6e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h564b8a561b987a57ea52bfd97b4fbc72a431;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf38206247cd9ddce2ca67a437613284d74a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42eaff73f37abe5fa0bcddbcc0fcf0cbe535;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h830594f079c2de5f99837dffe2adb110856a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40a0df4e37ca4ecc3d2cc5dabb005e56d170;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f88ff30b177a722204cd4c7a1a672e835fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a15779c1b18169a9df9bf44220b3a389bb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62fae5aa67456a208bb1c1c146300f570737;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h275802f9c70ba04e530db12e7b3e21efcb2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha52bdada51584bdb336450faf620a830f7ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h159307c1fc1d0e43d602436814f88e39f2db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd726b120ff79fa77344377917b18168f2df5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cd30e0f58c54aa27de1e7693511946e4f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4942a40a00bf9927f6ea12a2e3432cd7595d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6062d8fcee74ffd52065ff23bb5e036b81c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbef5af667b5d51fe712a541b3abb0ccab397;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2421bb86fdd03e49a5286f123cbc12061860;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h764e66359cb6ccc7073c2a97f3d4bb25dff9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5708ed3115afd66ece595626867b4c4ac5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28ec40beb93e6cfef37cd966a16c7073d5fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfea67651f03771331252840afd2122ece9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb77bf28fc407a8279c5b6ead3f2cac91cec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53e8946d4f903bf0c8fe66e4c180cdc0e7b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81642d2bb65623ff74f818cd49962085dca2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa1d00ca1fcb6a72c4647ca8b5de25d1969b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31c466f7575583e57e9ec1032047a8e424d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d66e29e24de6afdd7a36d04d8ad3cc0aff6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9412a4aa21acbeb1bb86391e7d91ffc222e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fcb4b6f7bb91c658681bde674fb1570169b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h983b116cb6607af1445cc22be260e400b730;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78c3fb9f642b1331b005219048c104ee87c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf82e29e8e2bf0d78baed5bdd7a97eaa192b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbb30a89890588a80596e053f56000fe5587;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a1bc32ed8ab3c19d8233977c73326fa4ff0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6120bab48dd9a5ffccbfae21ce7b4667e5b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf6434803b22c824101f527bdba02f257331;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc58c5489b3bce8dd2028c364a15c4147dc62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42e52599710ce6ef4d933a26150e2f4809e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h637a89bbc4755a74224a718382fb02237aae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f8aa3064dd51a46b5b1d2e7c2cc3a81eefb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacaef2190b9206f94ed9180c570449be9ead;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f086d0fab88829f11dda92fcc4ab0af5769;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf454dfb6fa4335d4ac1a1f7e1b416c1cfff1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffc1d0bde36cb673901e0b349bf04472a43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h995db8a481a37ec5136578287f5752f5d758;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1627df87e2c4b9a53fabfff1f85656ced59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7c6421cfcb7f7295b4d5ecc60a83ec0e6fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bbc6080b81b9d5aa421fb1c6b67b16ca355;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2473e072329b5478fa9d148f7bc415aa32a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a3d54d3064e841f079c2f08449cd476e2da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc4d1cdf8672d33e2628852831664c3c6a5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd578ce27928726e62375253a6da6d17fc2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb184b567572f7e3eef4fccdac45a28bbf662;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c4605fcc1b521f84edfcc9e52aec3668013;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56e7d896f8d75e59337181003dc889ad03dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed5eb8a0518a304f21ba158c034bb081f396;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6ece07af75267be4ac3379ba0bef5f0516b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a93747f8209735f161c749561cae0856388;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7a0af37acdc3d4adbf7db53288717d67049;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a11fb7e6bb902a2048dbbdeab7b47d9ef27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habb569043fca7a6397c93cb7054dce029982;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84cfff2346a583818d13bba8fed54f024c90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ccea24ff44ed52cce1dee53890482fae449;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fd839d8235cc5718a35e2d121cf9d1f3de2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h426bdd00b1ec70013ae044e3143e6d03deb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25cae59a16eef03ed4fb91a31778e5082ecc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b2c4e69f322031b5f4dbaaea547100ad82c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68ca24619bef12b8c34c15a70825ff1ecbc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcd32d0f9641317746b7f3ae11fa15cd84de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc79e3f09a6b27823824244cb4ec19a72720;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfcd5e07afdba5058186a7337afd12cb7353;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h917f57ac743eabbfcdaf5a0cc0fac25825c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ad57afdd24b8e0a201059b2f231736c0aea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a88a7e89fbd00b2be755c9b5e4d4493d06a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fc3ad0db3860bdcbbe3d007d5e2884cac59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20eb16bd4f3bf922fed0c20392d5c4a16807;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3fc09f99754f255fb5565ae30963aaa5ddf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d0ae578c3b7ed47dc84ba66737545c50821;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5493ac6ca14cddb44c3659165417c8580013;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6b7a0a1de4d30196aca03c0e5653ffa7a07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbcff8b79319071b84420ca83a219df97516;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8566d1fd92c8419710801336df131746976;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1ea4ebc4aa8e643e6a1e64e4f3d62993399;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h335b1b848de928dfe7fa0d86d5405678d920;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7b1903d02f809ab0b6c04a09516e0fcad4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7099c3446355ea8a8d24e15396cb860ef9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4af959bc57fa7c14d871bd6b21e2d187622a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2c3e3ab7095d7bd7efe33520fae71efb477;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1b90cb5d420b4ad3bb4ea3f144d20d6e780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a985476e9fa1a1715bc3def2330cdfcb575;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27ef54146167a6a082b266483d83113b763f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4918fce1dad4157ee78435beae9719d74879;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69588f964f4a6450aa57d729be6d1c3ea5e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74030cdb0a71fa444c3d88bc4a39b4201c71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h907853a7b749ff48eb7a0252ec67ea01d005;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77fb13bd4cc794563bfd668b03af3629111c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b1ac8b28900657f8ae5c75f8af496133b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3577cbb4968b3721655afd728a358e06ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0e65770997a0259a4099bd63d98eb252b8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec411d76e90480099ff015e98de4ca922204;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb740c43fddf80611526b5d81387c688e0de9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd493c59e5ccc415a4ac1af165d2a4c01ed60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66476144f8dd817f830f197cdf7b22d4b920;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dc9c5108cfe767ad2a2888dc661e21bb671;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0d3b49c759842905d8359dea79885030cb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6c744a94c9997ff699a7bc6d0daf8f446c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ba0f3b8b3418ea09580902bafbf4622e706;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a87535cb732e9a38b700ebcfe467eaaa949;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c300fbcaee1564ff447320e3a9deaa6ae5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd150315895b7e231cfb70f2e506ce6920e51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he87a7c4854963a77ba6bf9ac6b8d6ef415de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28fead9495c643ba677893039b3371f524a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95dd6d87280b3f7176b21befa7ffbc8f7236;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a8b58ec06fba20f56e69f09e14f43117fa0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f581a11ef973cf67c3a84fb390698db19ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he74638c4efc4d3203746deda08a1f388bfd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h507443aadba32f138dba27e0a5267d0b4bcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e1a7386096a567f62a87b946639e493a6bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66ac9931554e58690b8d7f25219fd1ed8676;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf67e1919afbaeb655fb56c7cc6d6c6c1679c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacc168c99b6cfb3911e9bfdeb40eb09d4f09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h247402287473a03a25459d01966c970f0dd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h499bd59b9b5c8150efdc77f32301352253cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e8df7614d31112e6d67a04fc658a8ee9056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc8f24cd03a237cb7f5f9496149ee1d3fee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc714881483004549fe5824d724364fc8c369;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2d46d685a60318c9f97f333776060ad01da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23badff9235fba0e3b7a619e48079bf2c423;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd91f6ca2ee0e05fe727f246d54ecd65d92be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a03a02bdac871b5034a7345138cd0899e0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddf43f53981f84f6e2a429e4b06096346cb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cb392e2a0eb824ead742b1e4e67c22c30c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48fe22ef0fee4edc70583f0277d765b0839c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23b989bee85fa9b62354b773f31e9a2a6b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3b75150eba19506d1e206594d2acc218eca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e8f58a71a2037a12a43fe270e08cf9c6a71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9001231293f536087fb62905664972ad90dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a78f626d1b508090aa3a709f883c5f01c8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8db2dce5b424e17b00eb94455eb3abf3b999;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42ffbdbbeb012d95744f065960048e805307;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had1ca38068a7896e9ac463d155fee1752190;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5d539f2a64db02d1424b5ac579eb49ca53d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h742cc6c18fca6b8a1bedde258f1300939e8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63503039f513cb8f002a801484feb0c8989f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45fe1e1aaf4fa0afa1020f1da282d6b869e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61e88a8bb120668c738b02c7906cd64de45a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93b1edf5c0d657d67e8d142d47e39ab1e7fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbeb47a17184c5dae6016778e50bf22fffe23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbf8c42a992a57b9a285d1247de471250f4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14feb9440e213a686b5be6f2ee7c01bf4091;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he75acda3fd2fe89064d1c08bfc5c6707efaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1d6a5fa242bb114bf03ebe11aaf9c1fa18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cccde8fbbd84051c5fbf442bfaab21025a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9609328c7e53651551cc8dc555629635dec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf509d313c39ce3040c70c03cbd80aa14dad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c56bd484b60fcadeef94cbd8b7194d3e53d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb7e356eab1f4480b12a2b6046a56ceb4400;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h644b12125a3749bc9a3a2abb1e9425d9ce7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed2d388fb69de3a21a9dc448bf9ef6490f2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha501ef69b1e751a247ba31b5c49bdaf9e7b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aa7741266c1156b6b786e34b4f3b856913d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he450581f7bf8bd944009142d644718f14166;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h764370918baac4b519df413570d19ef10d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbae80d23fb6a8819259ca1bb6608dd05ec9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c7617f86bca07b9ae59f1170b8d34fcf27e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdeb45936d373f0cc640412441a64e906ec37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ea8c16214285f6c689a191b6198cd5cf7a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f322f21d8ae6bcb957b51ba406d8d0736b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha078bef4177421e3423f2cf1bf53ea04b0d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h494de956ce1d070b7c0cdb9a8d65b198dc05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd77b2e5aaac6627d947ba971da4152c153ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc722b8e4be92cdfa19227336c0f8f716d1dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c7ff78fed32f169abafcb6959ede7a755f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb7d1fd1ca7ba6e484f997c78c2defa1d8e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha79eb042952236239222758a20ca400bd84c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7590f26f9836440de62611b2f8352eaa65a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1bcc8dac80fc1cb95dc8091af31997a28a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha27448d6bdfc093cf55706d14ae708a1abc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbde4fbd3e5487438e2168a6cf9991dc6307;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb16f1a161c343164a707036660a49fef759;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2b0563d048c9fd1c3cdecf9b770c818d3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a55660ad1beac39b3e8070a20a88bee5d75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee19a34a3bba5247f4d74261f5908fa9f2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha84f7fc510d11df124ec5573ceb63eb278c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa62e4a53ecc59e5215318d89d2c2f13b36d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91706f8bf6a969eafaa89c56665622aafa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h871876d8de0468ad4569d148be54fbf7770e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8cafe34ec40d6b33a9d8e5ccba6dcd964b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf90f3e81c8a2f44d065d1a3cbcbac6402bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdca62c4b1fb82615c57f173dc79f4943b49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he292130ea507a1180e710d7e194ca4b92814;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h265717544e425f3e4895a6de3d5fd4c0eb6b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73d98374f3332f69fca3d5783e89b65b151e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h645c77028301d38c9477bcb3d01fd35a1e67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7771150255d26c16604e6d1fc7728f2aaca9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44371917602d4001836b2f8ebd37eac1c1d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79fecdc134de7bb1693d0de646687924ddb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3378be18cf2524c884e34bd8d9fdcd6d7b12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc37e2d8141190606dc58db61095d9f8ef77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd54dc8fe0f9fb68bd61c17bf90f7cc6d5abd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b484fcaa656200a7676469bfe0ef146782f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5160afb3688e8429db5ebf52f96adcb6ec7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13eda62e38d4ee46ebbe76472d05f5015a6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha59c6a3f7fba1e7af6b806fbb115e6a86e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24f1a346beb863e960a161f854cdb75ba0fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h289975aeb218a10c1ccdf8e5f99d276baaba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23ed8646f9b6560d6bfb9dc4f8f5ccb3ff9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b00523d062028e502cfda28b8cc11b1d839;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4d93b173d06d1efca9657581447822ba79d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10bfc341766cff273fffcc48fe2f15b96db4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f028c760e674549b18c8e2fb3b9ebdd649d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe4a82814f3f70fcf45fff127f87a09d0776;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9136790be915e1700dd6e5b7e6dc43b75a7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5aefc744419792a3a23df75ff374bd16ded;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c7a510e64966bef0683a38775690f664391;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea68b940985bf27337880cfc37cbef9b4cf9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ce78126383da157dbf3b3b8fb53991d4ea5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h233a555498c5c9fa74ed74561768cc96968c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h768a6f48f9da8e2d19e97116a6f7c8284bb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8345600cb09651877260fd829460620da1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b227913650a8b117c9890b603ea05506e30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd132d0491454e6847ae3a9227d49774b869c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b15c517482958088d32c0a7a135b4f49040;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fa780faabe675aac11e9015d00fb1c14c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha77f6f619668b72e9268084bc30ae85f988b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2fab6090e70c6247e529e328e25ed1d690f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb493aa58e4d21ff7d0b5b92d27249e43f105;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63b7fb7567ec7ef0258cfaf15a802dad5c53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf69ef63612583136cb15739c5e3cd9dfdfc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d38be123d4cc2596ec6cd6cff079de43930;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf813d021840a66e612b2f7612f3132c11c52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba045c2604bd37e329fe545d3fdb629b8f86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2d528571e38cf532a5277a2c2b41497b044;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77cad01c67a6e677c0bca486b56877c31e74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45f47e1827b333d981593f90ac7134f00cfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he78764851ec03647ea8c413d5f74d20373a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddaa9858458dc6f62d30b138565047465fdf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ed84f1c6e9fb9469f7aac75a5c44957f3f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5286a4705dbd9fb6fb75b92fe5febc82375;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9178efbc50d16cbb5c7f98b5928cd74b90e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5896011ce3d3f2c5bc961e24203b2e0c775;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73e3d83b6c77b7355d70b53e52e8281523b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h864c41b27bfdd0e560950bf65f473d279b7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28df8cfd0b26f6ed2f613ee099b334460305;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2825e4fa0b4076a50282a22addb01a4b7b7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4ee40eace0c116ba2316ca8a39152f26184;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30ff40cea1c1a19bf3569b1740bdd8b425c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe5bde51b299cdae0259ce4d99892edcd58e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a6e1f6c35452ecec116b55daf100755a7d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6c9875f228fef278dc7b0de663138860069;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae2e5d4ab51259abce2a0b8bcb3291745a10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8467895c1bec554d72ee2941d8cdf3461748;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6e7f117f5909a1d5c31d7ef2cf1ae947826;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c0b732f1bfacf254728646291523b71d4fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc98c0c27ab0933ea471d809d116db341fabc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5317a62b06789a4b6df2fa212706c5267d96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd833cd85bbae92c9da3cda49d516f421dd70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88f9309f1b20638f44756ef0f6a1ce5df347;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h699ef17d4a1b103aa1df9dac2b08e4a8b392;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5043b0f1e32291f1a48d7b64b2fc7452a527;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd04e3009671f79417e78dfa3c2f440ccd2a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf30e65155713db8048b30a30e93312158498;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec49561d425c84f2b838ffe8fd18f70dba4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9e4528a6c9cd5fa1fb8fb6b0908fd1b33b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35ce38aec6e82057a7d666619f4c29bfd5a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6570635b19f8b8dbb9aae00932c86185bc2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa7fa0d874ae7677281af8c81e2a2dfe99e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h990edc7136fe8215719a093b003922524ca7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61b7c9e23f0a1396e8e3da1ea1a002626daf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h288cc8d66034f83bc1f645dc350382d6a3f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc5821422cded48659e25b55f991d946d5e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fdd7a3d6d9177ebe6b9f23eb0509774fd74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb7a2cd7d58b58d130bcf66db6cb35cda619;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fcca2831ff0b72a4e33117109849823b848;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a114b74a9c1b359c6a24b3ffca3dfd33baa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h973d733b30ad79e8d9c3d8515f990f0a959c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b5b7cb616da5097ea5208f2b52ef33adf5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b8ddf7a125021ef63e058661b6cc84bd315;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea23be29a975918f735874364f073c66557f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72b0e79f9f8a5f69f06133b616eafde6618;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fd54dc46c8d9aa063a63c23a124de67745b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b1dbf700fc858423731708bee17ef575697;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec9769224f7dfd0e57a84bcd11e11135a93a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd475dfc00ebe9cd81198807c4fbe012b1bec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d5fcd5c5562e8df1087ca6a0ba459865761;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca6bba64c712b767514870275ad229d60d56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92e93c25a4fc9e497a730773392c3d34377e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h791a039386075450f1487c005000d8983f39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadd8b85b2a2135b62d6e26afec6716987e12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb95c74bc03ae8709a7622c47f2330fc26b9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3c4091afab745b68eee546909d286f04f5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c2cc0716131a19f75bfbe9260ae21a41e78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefbe8e97904be97bb261757ec4174af3b78d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66517aae48b0ee7b9f3633309cb22384991c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf5585d99f588fcd3a3b80e293889dc287c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a11cc3369a716ec83376f5ff27876987d23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b13ed63533e18033e46644e0b2dba329785;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30d59d4141a223d2e88d7ee31465bd3a3e7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98a80068d30a2e6281cb0a8dd0cb638b895;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h885454e89c25ec89f56e145f1ec57afd3b2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80da4f72abd044cc888d47d5943962d5b22c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dead22b2b6c0d23c91606a77e0c56c212ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h482d16f3d10eb06501506eb7c131491f6d77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd0d5b4258c1076c0ce1730b67edb291ab48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51a68692cb121876026224a403f47db5baef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31604e57f47605cf54e7dc3363af9981750c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde6dfebd95858deca97671e620a0f3dbd65f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c25b342dbb23836d7a38fc5836c6ec29f13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d50244b375ad9d714830afd239d664e2e87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h674ba3009978a86b5320fb375de46a6364f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed5086220b46f12b0dc4e839f846eb135474;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h728280984f1149e120a993572f91e3b7480b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40815ac75f7383f6970f3a8ab0f785c43d0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c411231f824fb78c731f66b633ef3ed5592;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc44570fbcf87ece0b89b2235ccca88fd3914;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22058ddd94b08c7aa8b79854b7373038c2ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h846d947c5e20a16fa1bc9d5158af2725a805;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h214ebbae0bae076c0fc9a50a87f4ac02d3bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h181559b04d0f7d0df959add9e2f1ec4131d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf958fb88a3f556c99efb01d66861ede58cae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ecbb080f4fa93b397ca34eb53472400d802;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82367efd732a7c87975ad8b06be2a668cc81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h628129c37034205fec807b7d603346a8a2ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46fccd7b2d72f0d12685d13fd448502eb4ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc95b908743b1be7f7e17d32ff5a1fa27236;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf4ccd43ccef98d1c86e1c9f4dd9cbfe1313;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79e1e63ed95587d7df47ebd6c6005ec24319;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8334987a1f832c9c5a018c13b8e7510b5f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a142623e54ce20393884e9477726ba3d3d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2e3f81d312aa542bd7ce827a47ed762cf22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d4313f5107b22a81ee482d7f99ac2dd006b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6442b36ccc7617db7008830518df106bb4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a109b18093dfe1585ac0acf6a8e5d07ee69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4db618b63150fc560df21ae8a2e0eb931caa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd17a19411a91cd919629de21cc9ebd574ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cc150636218960fc56b59042ce20c7fcc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8de215f2eb9d148170ad1f7bbd73fb9fc461;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb293563e8b4c617fca495b97865cca318b26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79f62e55917dbede581971c1245dd2ccdfde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14e04954b7fd189b38aa9a6d0a944184390d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h267ce31560016de42b2d20847895bf054f23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33152479bb823697c30bec61fa1c1fd9e140;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9046a6e0a72df67a178632a5e7cf08f8304;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfacf86ceb5bec075e63069e87fac671cd71e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h547d99971f6c579108fb97305558ee876ee9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94d51390d17360e2e30cfe573a107fca5904;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he27aa93101c17d995be20dc33af12c2988b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0545d270544df93c117397fd519d3675908;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b5bcc8a032100d03d1eb73ae6d70f8c7157;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc2bcba256713372740a127ced3a235e2509;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d41c9cd214ed3b49bf2b85e40d6e4e21a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2852cff3f325125b0ab614038b16753ba71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf36e91c8885bd9c7a0adff2cbbe0fbf0aa3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc7256d4e22932492abd21921d7c511e2573;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h732f5f01216748bdeaa2048e9b8629df2a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21f18dba370f2e154cb6f2cdfedc9b85e56f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4556b9d8fbf541dfb49318f91b0cb5b3480;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2758db1bb39e1e25eb3a3aa762ac91d1714f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c394c88e11bd80bc96edbc711b13640648b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d57994b6c5b1e5cb1657e11bb650c97514;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21345e0837f063f6ed609a0d8ec33abede85;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f968775d4679c35761f2e447d8479bf2cd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bf22d22c4c41953ead5b4d622a45f2302a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha901e60a27f9795863dc80f5014bb81e1e73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h536434c019180949031c9d19e7f2a65a995f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3154f40dadccfd9be26b5883df265eb8f5bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67548e4950e7de92d4c68f68db1dbae68dc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c0e0229d2cf26d4510548d41dfcfc7ccc6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb21f520574d1c2532757c5ba4298bb548dec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac6eebfc40a83920b3779aff6c73b80e2aaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75a4eecb877e37cf75489ca9d622217bb0e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc7e2638302e8a039c3f3b4541605c769f5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9dd7f73b6d591107dea5ada346067608652;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12399124408b2138394fe6ac2843cdc91e80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h949521b9cfc406920d8bd683eaf15f25dbfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha71bff9e7753e94d0fcbc607ff4f345c3f91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60685064319850f8f30aaa7b921d78dec037;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1c997b4ee7c3c25530ef397fadea5f31223;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1179d15f9caf1994a57644002a9bdd780b5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h823e79ef8a2f6cb7e8cf20987240775ff774;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5ebda1c965e346682f12f96683ac08f2f1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d189191c6be90979b03260add4e881a7dd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd983b31470dce812f4bca94359f77fe1a088;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfac0e997b172413c9a924da0f0135bc546f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7470118174f9f878b8d6ff2ce289ae37d420;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf97ff1e896635cade9a5d9427cc4d23daec9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74f3553e7107331299081bcb6e91583225d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a999b06afeb38e2a0403c55d7562457d38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89a0ae12a5253d8e547c2c3aef2b7a39fa8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6c18a863b7d54487ee5f13736cb871796a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4bc09100a7cc7ae7d72ea6c2c9bcf93a9e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a9660a325b6faa7d472ee08632869b22439;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60f5179361fb397efd443ec8806807ad3701;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7cdc02abb4dfbe78d3363b51590e7d8e617;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8560d87fa3f0869da28d8c224617fe3229d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16354029a85197313dedc5793eee981ba5fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f2d4ccef4aa7d05cbf3c63be00cd292d996;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha16698ef206e83b9111214c4691af202a9d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d176255db77ec04add7b39ee1bcc9718800;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb243621d7a10c8e609787ee3dd9e08d9134;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea4ea42a760dbf7619ffb5b4fa6f06745906;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a32efe79e91e49961a63a7c3ac69c47ced5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe5ec5ff8df9e4c85261f16ce11979fd346e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43c39bea8fd02a93f10cc79f076509317c29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81d17e9d31d322abee525818433e2fe225da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h490fc7d5e8abc75c7b621367e542ef42962b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cc10b6397bcdf29146d0cf8d74ef84e101d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf998201b4905db8a7d3116b95013793c424;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e81299bfee6ef1ba79c102e7ec3f3e5d716;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd55e4fcb501302e0164c10c21661dd91a09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11a538aa54317fccb7e9db265aa1efacd298;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd7813311e2a898bb140e49002aa173c2844;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7c42c2f012007642145ed05b4af52bae6ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11c35d8489a9e548f200486ed83fd69a3be8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h998ed112cbd1aea079f8d16c24bb9e67e16e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3136e93f27989963c06ce6bd2dd61e8e8d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f198e629520e6b7e7965a9e01123ed6b07d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd799f2e7742dc64ea5b8e7505c8a4dbeb9f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cc39579ce89c29953d9717c1f1611270867;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h722eac3d694fc3327ddb81542889891c788c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb38c1e4cb1d30d111bc6530e256fca097e75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf51967bff54b2037e8e95a3779d3ae6b4ed6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5758b0064915c120b8bf107ae9c828fc3d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadb077910066dbf6f9d8625ec0dfd5e9076e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c4795754483240b9eba00f5385eaaa4efe5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f2c397dd85f38f5a0b36c6d40274b71a73a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcd187d482257dd43eeae577c28b76e87943;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacbf0ced578965a6e27a33d4b5a6595344af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb14707afc89d7ab3a08dfed72e3889b04f91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ed3920bbe5b885f8109979d1588957311c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99246cbf2f99553dcb98bfc9eab1e17f58e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c66151bdd4177a004454e8779777f9f1c05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h555df1d6d47b4f2f940d21947a0fba13daea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cdb72b6acad052eca26d655798f5b0cd58d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c91db199c02d462108bc548601d047d766d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaf85e1ae64e7bd68c6bb9f357b6f4afd49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87d1bee32df9fd60d30e712c6ac947e4a7eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5664ee992e3bba0e2564ccd8bc2b6e8298dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff5290938c73a348d4ecd95eb17960231891;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h849f2cb9d16c51170b59a9f8372b391cf26c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd566394b9a9c3a12469f7938ca8dd468cee1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1af0ae12c8fc06922a5dbce26b1e0fd5e24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfef0584132c4228ee3f9dc7a528c56bb3a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdd206c6593362317fbfbc26c325b1b14fc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8aa419abba9443d1a142f7473d06e39ee06f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cebcf3dd27fb83c02c7ffda153aaca44737;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8abaa1e49f7fe9353df94a749f65c5d11ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70689ae5c0796c1d2403ec99182daf389b1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce955ba3919e0ced614e093f928bd6ff518e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbaf4d8390ae0b7a259729a9447c4db4a175;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ff43bf009af56a12c2ea20a6dbcfc52c8e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d5a03b21d32771f8bd07e03900da3e4283e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26397620de9d166ca7e1e21b991367c09bde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he42deb6dbeae6f2e1a7bb87e5f8bc43c66a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee149e5c728d5736ec9a1b90cbf5e1ab7a64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb565fd252ae6cba8001a5d341c59f196e8d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47085cce5e19184e3063b7390aa8de2d0531;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc332973767added171e793251441d742b1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55eeb58eeff613fb424507488334de4cc05c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4acd96e192d3fdfff4e0d4dd94bd20e406;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb58d3b8076a39826d8888d3873515699adc4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he434ae99fe4f0652bcff472b587c32cdf0cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2399fce89725c1113136857f8c481f7bb694;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f6e4886f27b73545fa31e12ccb323d8d308;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82c66b1a87327908ffdd9a23be97c74fa05f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce5055385f1bcb736d91796ca04a2aab3f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc2e25ad025b0e3e05a2c91033dabe3a228;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d742030acfd39311058ef9f2d8b454bc055;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b0ed9e25daa9a40633c49cd787634f597d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he34af4c57c22bb6a32f29b0d0fb094d5d40d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38d2aded3403c8de5dee75ba7d536b6bf58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47d2f874e58bee9535533ccf3f3c8d64e8a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3a1795a2c683e436f0f4e8a1a145696a8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aef446418932cad9464fc6883effed925fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3969da43ed36020c8e57c35d14b36201999d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bbcf751f1904ebff178a7cd4870e4e67dc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc458c622d76fa10ce2f4efa53808b56dfe2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61b39266c865f137be0afd3a9b49f809c9d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h649627ed05700b195c5285552c4dedc916b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b541b497fe96226515d9d69eb0d5c5d7cd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ef7ddb224a14da19696a3f72c960efe48fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3ca1cc450769a97ad7a7cebeddde58bc503;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17f0d9a940e4b5303b6452d7b4db00096178;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53edf84144ed502e99a4df70297e59dad5cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3e20fe8be5b1f53579b227a4a6480ac9e51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86a7a1ebb36955601d7d5e6ddecdf777521c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd475e2554e0d271f16aed3926506bfe08f4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5ae54bc06ed7ceb1e88da8dba5ea0d873b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ff1721699caea3c23f15656eee37c83cad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5c96ee03f941513ab7dbfcc4ca234cd345a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8643f90fb45ded2cfeb8ef35a2020df6fe2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1fd1a4ae96529f17373c16704ec8c20c6cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21f2f4a4930da9e89467b0f491406e84fb33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c6a1b7a1c5c41409bdfa047be9370f3ba01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74d3e063abca3f919c833c7ca0831c1fd803;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5fc970154b5ad0f3042e63ca9f0829dba153;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0cecc04cd8e499a258be6c2fab480f56e68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0967ad6ec67bfc02ca1519c0d4051b9699f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6885e1d46a9edc0fbce78b0234c23b44e62c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe72a7983c0dc60a86b2bb18acce0cae93d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfd59b018bca1c3b65395b534fdf5704db7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3223ea890f61cc69d9d7afbf81289585d588;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b79b325a93a174aa841bf1202ef8eee9e39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a3907fc4a3911f3f8cfa09f3323de6c7a39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha542f62403bf5e0455b1459fdde8fc566399;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfc76d07621513a5ac230acc90361cdafdc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5ed57d40dad54f14dc6500946107c6b1912;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e470cd6e8e49564d810c094ef1b5e4ba8fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h107326fbddca7567a632fc1814518c0fc69b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc09f5559f8dcac57acc0594472179aab756;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h811a693adc33a91d052e479c9dbb688c768d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74e1b5dcc4407adf920c80b93c6058e9d933;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34dd42ff3104996ed6500d84149f185e9a72;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91ead184750a032001f55902244a09f99368;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21956f49227dd0f8d41f0fa32f929032f0fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29be6ecda5d7f0d9314464369b5febbaa9a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dd2e26f0d92667af0a1f4e38407587d2f84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h596a5780a8810e8567943ba93ca414d8bcc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab0efbf9cd0f38a4c7f5f79c5cf4a0daaeab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76c5df157e00efb21465d965e20324ef5bf0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7ff2f55353adeafd1854b2cca638104d277;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecb3c4e4fda0cb0817c721bb9fe2c9e1fe15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1907644d48bbc869e9323aef53bce6df7a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h353a6c28bf09010e344c4cfcbb9f26edef3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc08fd569b3ddd922c4ce91bc83cb0ff6382;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6be714fb89b7eda029eb19221b15516066d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf252b615a263e57ae9114d6ce5a829dc84ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84e88b82793266e21af6973926e060b7ef56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5685a55a87ed1bc18478ff7f9541902bb60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h406f77864716fc96a5c8120d24d5c7e1dc3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9277f1dbaecd5d8286bfb595c3a9d6bd831;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf51a7c021615d33d0f1100aacd2639094af8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6e18bdd222f1eb6847ee9f0b236b4ab42bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1ffba0eaafe2745b598f1b7db975a7002f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h714229833aab3243a8b3a3b1622b39d291a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb52367fdde6fb1198a326db436861ab501a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h445a024f63882c7cff409410e5279e64b0a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d11e4402542bfdf7bdf912f8f55ec7aaba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e7a00c1e37a9020b3e2b64c82c44cf14141;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdef431bc23f1b763b197c21f0bcd5230263;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h453db074f49bd0655e2df20146cb2eeae9de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca02a1906c5101daf3d199e60b69ec45df71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91292e431548711b507831384f19e26286b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13a3b6a08d93debfd79a12d4ba0123467358;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe3d25741c80766b20323e5e0915681f21d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbeab04156edd3dab9599fa39c2eae61bb902;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48f83f56ffd0433fdaf861ee43c378c9d69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc59bab6a10cc81306a1030102f42f1c57df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc88f84493f7bfe5ac336d983e1b1ab8992ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eac1814ed116ad428290cf143a47d71c999;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbec5cd049445f5f5c25873e7b63d229fcef6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eaf8c929fed181f8fe933d15ecda95598d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c87374af96047068825cbd5a9882169374e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40cc1604100099e41553b3390767b1679a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa7a2a3c0d121a17f8d607e118895e0d89c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfebc914d5f84c1366daac8e4fc1f1f7f34c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dbb9d403b1a8b2c02496e0113fd3a26ddd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h827620fa8f3eebaaf3dd4b03c2b6435b9357;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e82ec3e68f0b2b905fbdc87e5d46c8c5efe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1355d385cf2e6373994f6d6a954a08d43ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdddd4174c5a1976b6a4100996b46e5d25cf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcbd824553e0d00de07223d2eb877a8eef99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e6604a42fd13bfe3847ee28d0d31069c1d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b1adff1b995d398ec742e29b3a9b9a126fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4ebff545547a331ca2ecb15267933d9772a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e66d13b16dfcd6b7bac795bc10fdfcce47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a2e0fa26ad483506b4badb9e4df8a9408c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8e7b820ab624c58ee5510e67a1c0b509e04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfd12af303d0a19574e5505972f5d5bfc2c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd21b33cbfe962075f210338319c74b22729d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h478faea5f55e1b6cace3e26ced403b19994d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha812598c6bcb0138bda3c56b725a7a535da8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57003baedf80ffa38b5ba7e1757656842ac0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h382d02bf2d7cf1d540fec743d52c860e7200;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77a6fc63a880cd9d51ead9092641ffac7f81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h893628b21c561e0ebe380e078bd6d085c9ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6d09e3a1ef1080e7d3fb229ed33e45dfa66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h603cc3392d453ec6676ecd123a8bc2352ce5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcaecef22a7b58ebe9d7e1bc9b0eca5340045;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b93b4c592f8b02eb4593245aef76af93306;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9ada37671a3305be25c75ac6249b5951ca1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdca5e00612903d21739adda5665491a72419;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda52630805a415d6533d906291d142102c1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3de8692f8dc9de6dbc4e3a757ee98609749a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb00367b89e5414080c19f8aaf51707e6f68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80a02d42174c7437ead3aa36322acbfd8303;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8252f654df50834673402a9f664e20ec712c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5d281e172c5926f4b5e09c0db0c7665ddef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34f8705f425026ff89cc711c351ef25257d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cd8d47b31c6f3181fcdb3b7bf1cb443fcde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc60a1b8df04e25352a95a0bcd1a5eb042c1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71d4425eb4b3e13b7ea9f72bff3e5a34672d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h826c20de904110ede0ba289b5cdb4b95a03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae3ac71bbf89840305bf6aa610da02c89aaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd355cc5e5755c7bb564d7a59866bf04c0a8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3798dbbf0f7a372f56bc9ddb91756d1373c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae52a5efe1bc2e624210125efb6b5f614ca3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56d5e00f0fdc121e04cf1eec01a91c1ee4ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4688c87a6b20b105c299c12169720dab2063;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8eff2df838b04692263f155e708801314d82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56262709578b08eb84d303085188f7a260d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h173139f1eca1e7d6e55a54ac09c4737b2512;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc957f7bc2fff51561ce56d9ce89fa9594ff9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac153568e57b2a0334d15709ac8305d347f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4d5d4150b5e608298d523afef1d7941dfff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h202a6a4d6a97510f1b26cab36969f6bb13df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89983f9e9a21cae996110baaeea3285609f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb06c9058c2468e68fa5c6691dafe0038b8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h628754af80f0638cbf4e9cc160c82b8c3ef1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc43498fcc058c5d42fe55d6b5c3768905f1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h355f363662cf6c646e628f1caabe7547715;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aa62c427762948e6a887f449a502a9e596e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf564d73a1889f7c40193ea9f8d189239033e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11bad7152344781f99a462c093802d83ab30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48c96c87b800fa40d42bacf549d94ec3060;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbedab6cd7ef54c24f202a49d2829a11ac872;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf69b679367868d1c7bed0fa0e5a3fb55e5b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h315254df4f26bbd490f38be0dca8f698c1c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2ed6783f61b09d5c23d94690cd2cd77cc9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb87965c697a184e95d671963f2af69b3cc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34b612eae70b2980e04c66055e93c17d6652;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25b5a144a6ea109202bff6ee95ebc826cb94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h340695420fd7a1fb5fa55ecbd71eda8d158b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd205183ff4f8f61b18ab257a6e69c4634307;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ba8fc099cfda3d5cbf4879210dfe948250;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0a02e49ad111d41337873334bcdd062f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h499bd09f7112b440fd7996c9bcdde8374ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb606ee46792ed35588e29d6b10b8269f11be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f50df8fe66dd443563b98752a0b654e80eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35c913a3fcc02f969c1d8be0691c8d4971cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52a4672c0037d826681a1f340ee9f7b245ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8a45e99bfb23c8a5cbd8e11fb306cfd562e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe63a819bb763ae280a6c833f174042cf099;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40875a4aaf27be204087f36da2688b096d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h419f3277b979673e948eec9de4ca4f0712b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f107acdfa3ebaf3b771f010f4e7bcf2d3e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91125df1d4e72d1d71c157d3bf87b800f25b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28b515299ffaf76e36024f2a052159713261;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha12c5c53d8aa7001f919e4bd74a8f1fcff93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3f9edaa308f3dd6399b5622ce37dd52616;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23d946d5a5237feb0d976894040fede74dfd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc77fd4cf90f906f15a4f323f9c73f59b4ab4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd58bd400871d3b5a81dca9da0017a9037d7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67b6943ba41b8b2b01ba859063cee291a76f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e7e4dbef012e744c82351dfa632e1177c22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d20f6757b3e0e1da52df71dbcca848b7c50;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc1f845278e153cafc7a87edca9a466d4e86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b1c5b09a03d7854c08c032c49c4a4da6986;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80ab6b8d627341ac5e44d812ce3e692e8a7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20a34b97c3f24efa995c89c5298ccc40fb2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3232a6f52e97b80528ed7c8c56df3d75f72d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8729910d1a2be4125a95ef79c14f9c37a634;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf033d2591923e68f9d49f6d75a6c12f2d40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69023e8fbccd29be8aba8cb989e831be7097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61dd32e2291aec7159d66903fc0648e46ee5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6985cc365c6013df98131019efe41162fbd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h707b5b2376dc9c8ecc708e8a113222e307d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28bb27433aa2c144df3d06e6455dea204e7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7edb3929a85eabcf66ea390ff4bc6780506d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fb3b6e501c3c59ad45c1b21c2902b1d958d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71892cb32568547fab4c430f8fd5aa93e742;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a7f349e4b2894cc413cf40f03ca48273f16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f116628366fd404bbd791da13508dd87e31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e01f75684c9cecf16d5b8e5630296423a6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3bfe00eef1d4c778ca53b8455d20706e6ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h874cf0f602c9e62a572745ae46b0420648eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75d14cecc233234989fea28e6fa812f95297;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf77f8f8f1ac15d1d284b493feee38be7bbc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6655a4b39ed21b40a17ecbc93cddcb33799b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba125c93c7eba0df9b8ca0b49234c22ef6c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h490e0a14da15d99c2a46400df07d70f18d28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70e204670e1566f62b67c72668c612f02716;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h472bf10d5166f32367347d465afe9cf7b282;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c647ea85357df4faddf85722dbd4559412c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90fc3b5d1447d4012794360fdc9df10c868b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1d7e8fd9dbdd41ce0edbcaf421bc6367c2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b130e7a3e2e4092ada987ca947b4268c777;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h142e948d38fd2c8fd5038bba8df31255c0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2bc69264f161f6e0665a18069ffb931e39f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h345d1dfce2d20984b06a74590c22304a20b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddc0549cfb950bbfad7f6b6903d1b4fa50f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21d321ec480e72bfca0fb89f7411ad586cac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h835fc8d0d902ef54a9b086ee026a1f3c8a08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2995ee1462a8afe5275eadf2e9c3cb0297e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c91a8f24e2cf92b45406f11e17e903113fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9027c17d3997b2eba8b256809afb809b25ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h900abdbbc5cfc3850277ad474177f21085f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefa2fe216d5bb099600a01b5ffdbfb8986e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4b7d05457cec92758d117a0093e644ec215;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h813de1b3464b16aa3c4506a9246e9b2a611c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha62d82822dcb6d96def3c82483055e238d70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91aee8d768784d298965fe0fdec8ba486518;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4582696386b51e7e2941e2113e59c2cc0c12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f549b58cd51933ab853bfc7c1cba305716b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h378f411446494fb2a4bfd016133ec11a71ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58e807aa6faadb0c10b2a90105c0a04df82d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e9db5915560ac8e437b13f4a3a16d44506d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79b1d0cf09d34bd97627d8e71c4e23105f56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf174a62cefaf8f899bbd9906b1d2c54be8bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab077e599485a6b9ea6049cd9fd0df80151;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8e647364a7281dce275896aabb3198554b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8dd3560166af2ba3c98fca19f3493ee527ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7d7d40570894ed6b8cf0ab93d6465ed6a65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e0c04804b09534f4753a904d8fd5d4022d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf47b9a62e57115abcf443a50b8b4b1dcc4ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64aa4d96e61b194e4dedeea33e5afac6698e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82d6a9e91e5bcc4de457b5385d074d8ef2dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd2f4cac338227bb86e68e4ca6d0f2cf230b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa77113550c0ea1ea8becbcf113d96c87ae9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5c15879ec0f917e3b2ea5f966ede113a7ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd4bc46b88166a226d9b566fcee44a96459d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd1e812b24f5b707578d13762639c9539ad5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76b5cbd76269983f753b3b588241d51c81c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60653a25112acb2a429144e3c0a943559f3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dfea9434fa4d4d3cc58d7d88a631119426d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1d7b93b6ed15f0d7f1e8a0b87736ceed3fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h788b817d3e932ac64a34fb01ba6f4312fb0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc725d5ffadce1a4b52e080e8d3c6f4b8aed4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h558517c3539d0a2f65b454bcb3c654cd527;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h630f12c68b4b9a7817ab93b17996efaa9e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbefb34c95c5ec73e4e42302988b06d8ba46c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5e6d38b8411305e80f123c007903789c15f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cf58ce5a790db46106c4ec90830d0e01a1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5b0d1ac669b8f48787f530d4768ccaa79cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'headaf762b0d251d2199739f8b15c07b0f7b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h833f9b21c1edfacaac5861e6960b45a87fdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54b1f21c8b717ed5caa7179c84c82f1345b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82b1f85dc7618240cfff78b5df620c997efe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac30cf16e094f37bed23f2e8a51e04f5b13a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6dd2410ac80dc538c469574a6f8109342d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14afe77848366c09c0f6c09608c022b24553;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5bdc27e7b0ea805020583df80c6de922152;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee81f467071b0cae2a2e6acb6f6f34aec560;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h521ac972c0669f429d0b33bca49c04443d98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h376288e6fa17981aaf9c6b7ed38c58609abf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfeb00544ce379cf596298924f06293f6d43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7478c375b673e261a710e9c30eba8736cfa3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha75c1804a9da4d91bd453922effbc16b5cc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42061d36af5e146b13c45fcd54a8af32a4fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2f69ac34686f736c066dc59266517d4fd1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82f961b4624a6b5d3f7f8fa0bbc2008fa5ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc3037f41180e3870161af81c62088db6874;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ee4e6eb917e2545a1ea6c7e828b7d28d122;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac3c1b64c2dcbd5f01757a7287693a7dbb95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90b6227034f71e858dc21942c3acc1d757ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd1f13e5b54da490f794a68fc3df604e6af0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9573e05a2c15ba9f14d3e714dec19f0b5c5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1091a7178e7d314fae0f338e0655f5a26f16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69167970fd86f1dc1b07c7a304f6db9dab20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h440d280bb0d163cfb9db6dbc3f10dd8b0b51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha016caf8db7e7c6835df6c0388c60efff2bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22dd4d0a2b68f84810368bfe47c496689623;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h198bcc26e206bbfd731fdf05b3e830a52621;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c3424836256435becdca74792919c8fe0a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he621a347bf49b5747fd485753881592b9792;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a29f370c3bca338eb9f3ff790edc4609362;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb8ab526c1dc5ba151586e67f9a583507377;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc236916553c7e8b1ffe1bd2e587b1aafd2d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e44af5659f17839965da0ef7fdd7a44339b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb74e57f7e68f764162996dfcef6595cde616;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10dbb93fb4f90af2ffdf9e46e14db9ad8089;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bd29d9a122682066ef3251bb36475df19c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5fdd5f57eec321152263e7e064a9a24e0d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50cca71f5616d1566ba79667edb4abf6f8b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha06b5ba8d9d4adcecbd3015e8ca7d9fc1329;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a0beddedb784db85aa15ca2acd96d325722;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d0c9985c387f6d0aae51919669658ff45bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc18668f023adffe679984c2ff5afb5d5c1f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h157856d011d5841d990d9c395246a3b61fa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h862f3346ec92da93439b90e9570b60746b99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h378a8eff8edda4f52622adec34984298035c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd513f6caa8546ad39ea5fe98828c68c9a5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbc6fcd343097ccc13ada73b6160f4a1af13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb49f127c4fd75dd8aed8d1d0c7cde61dc5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2107d6c2dce7cce48f90124b4d8150df4a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab1451919cb3e21bcb350b26eea01c7360f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ffcd6f17989bbfb2cc30a90ee00f9dabb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h612957733f4a48a6e9dc376ab20eb8908389;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e66b975fe385633e481676e862d7e024300;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4045358e9d92c8bdc97f89e33235bdbc7d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d91fa0b1822024cbbd25393f87ba1bb76f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h631f8df6ed7f6b6994b9ec6970b1f7ed02fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf785503c7fff16d35646c9ecddd1afb09436;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59f092449fcda4bce73ec9785b122cc23645;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39b637f8aad47aec0f01e5351559027c112;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda14307646edf61967b3254bc09e1175393;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc67b799013591d0ff25cb6a46b9bdae5b1d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3151241f68dbde05dc5b975a28d655e6b54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd14603c9624e115c83d9ece88bae2501308c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8130b8592a9fea95cd1526a2361e6a426f78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e579c74c85ecfe7b0d728f2a894052eaa0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5570ccd543354100442b10a3793f0835f289;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd6525a72de1282168776f27d33f58521169;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35eccf33ab8fab42c35174d2a1a9d5de878b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca976eac4aff15a36c542ecef3a55ead0f53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h453b8a0775a264af6b0718c4e9f6d425ba89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d496accf97c4fbae5c328811a985bfa6420;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99d7f393490e5be141af56762d2bbf144f54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bba245daaedc6c5e46197a8b7adc43c50e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84a1c6a6311e0f7030e56294b45a702a02c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcc07f701b75721b3dbbbc9c743deef05ca8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75f69ca1bb9012de5ec0751f04c22693b978;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cdcd0d1fb6970713a9c012110043f8611b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hada49a8c1fa08a8ebcc99361594c9d8612c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e916ca82f900c923f5d803739ded504a340;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e3be9aca8b1eccc3f485ee570c654f061c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28b3575091f74a932c246538e18f4020d709;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1dd2d777becbcd3614ec1837cadcb28b141;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dc3083a848213fc3b60c5cd49eb1de33063;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f4e93ea306bc91df782cfdaf6ddfe5c0594;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had62601a6b76f0fdc0d5a9ea5bc11292b9ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h815c34801b25f9c2224ab56616ce42a12110;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf32c699e79b8e7ed15c3ebbddbf1d1a1447d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b5d7e0de0e036da7065a39e95eb578ffaed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3249598c21d1d18b93880dd8fc1119e77de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1251787e81626366e19dae068be351b5b202;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf220d429526d3c30d29f4e0390e957fdbcb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f0a5f10b4ec1fc48c2d786d4604c31adc7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d50ff2d31e1af73955ce9ac22e6be10caca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd57a8eaa8e9c3ca6b4225594627537edef09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25896b8079a787eb8957f0d1ef673c807b9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1acbc5530559204f787cc951721903ebd9e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bc681c7d53337fa9c82f14c6822691324f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45e23714a8b4bac3ddbc30256a0b183aec57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h944ad1246f8112d20686d3c0fbe063a0fe3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85a0c3040eb02965a774aff2a6e4064ee0ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h633d63c2eb8baff33d45f6bb90fbdd334cd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7869613441c6ffdc0408a40cc2c317ef2ec4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f8a7addceba32c5993f43f7d0ac5e8f6e46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63041ef4c507125746de14416bce85518346;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he68d90a03d22619bede163aa269f2f7f3b10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5a0e7b630daff5b5f5a594f65ddfb3311d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffe9eefc7fd2b7bbff768d99205f8bc1ff62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h197b80c8c9af14528b9e5462d7253cdbe0f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef32f8686feb02ed42e462b3052cf8d728b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h855470603a5e375b7fdbe084bdd824bf4807;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h488efdce1d8b5138088ff3de3adccfedc6dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h575b02307cd5eb13f0949b8f5b23bba156ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a81bb326c14aa36243d1a978020acf1ad0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc98aaf37bece0b70959f74f3bb9ac50b56b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd90e5c397fbaecfaf57c39bbc0a34f58a80a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c979d4fa38350e12e660755d8b90042151c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h230acd39216d1f92d40be66dacd44005b6bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf03fb564723d5a0217e129728cdc7d9377c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f2edbee142d2196602177a0b17074ed281;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca832dc3129ff85b3aec68825ec4c8496070;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1435a8aac503ca52e8fffab77cf0a1429ecd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cdd1b7e1ba095084f8354583a5c375bee2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbd10f638fde91399244ecccc70d36721dbc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1518150f138e0182630521fe52610f8be6cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1eadb90c0a3ba52bb4da33be718d50277e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4dc489afcb4896e4f2a15eda199387205b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5cea620596b96941b9a6f9307c964c8b9a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcaf087716041948d6485eb0dce1aa0249e3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb572272af4d0806c0db75647e3758ed0ef10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he368f6b8b65f6b078fc7733bbc1887c1d016;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56431b21fcd030a2e3dd57e2539c5796ca1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bf3f04ed86e59f9d77095ca02eb7d2599d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33d90227d9929679b86056543ecf530f8e40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4d8ab2e5dd40f5f48a9178dd0dbbc8d9677;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf29412722971cc875e488a0d11e1ffbd117;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a3f534ae6f37580d0363f94670b7a4fbc42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha03a522a556f1385f8457379d3af38fb9ef9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dacd0ac7e37f14ed4a2f3aa721efe99dae2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ad58f23dbb3a10bf63515954067258c6de5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90fd2ed41fe38c7413e58c7bd62fa04c5a86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f9c105447a25b6cc98c20b4eeff82d5b768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1712e11286f133023175cc7d2b8e19b8dda1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cc343af0d6226c2f72bdedee698acdf222c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bc4002d86ebca11f2aba0616d790ff4f6de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf619686efb7bdb542e77fb5363a36623e264;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aa76c535f3dad8e230112e44ea1d3168a8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb0fb6b2f2a76aca39deeb02d0f46080c94e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95c3df78c02f579a0bcb469728f59af43315;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ff86f0beb7c6b6dae7c4bbfab2a4a71adc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb767a88c6bb33940705beb63597fc9262f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee01b975ed299afb9a370aa38eafb9c724c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70e82725a84288dd05d3de886b052b377054;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83621330d49bb2cd0504e5d1f97199b1d31e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e6d09362c2eb4b9e867125354517b2a45b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h980b39ac03783a84f336057b99bcbebd7ae2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h150f34387b48d3acaf37ba3ccd73968e92e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a5d6571cd4baabcf4e5e101453281ed7900;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16add19c0c1d0a3f0db24ce111e5cd3184b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58367f97a2c34dbedf7ed305b23b148c2441;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h704631de2c9a907e3ad05c9f181428797dfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f24004eb6d2de9acf7d1560f1dda24b671b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce7f032f69dac47b8efa60028ba79d2b6f72;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bc153d12f9c5f47cfe7cc5ebeb0ca86ff14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8d1620c233536b3b3a3339e16e37c0a8296;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d9c71640fe01caa80475aaf0a5118cdb32f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66d2f16ddb7b1cfdacc7f94c8f0d01e79d15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11e354e661ecfdcce726eb3e876442c3009b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dd16630c54f36a5a92f72fe3f4d7476b5e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b45d074821cddb37ca769f0e5a748f7eff1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9898e5728e141d9b2c301c511893c96000d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4038e64840851d4d8f30bd727886601431e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44c2f1b60b96b7b308256a3fd6bb118003bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1af101a1e1f263e235eddd700588e83d3d47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9310248069576ab34f9a1cec8f54f5ba98ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98729eea8335378fe504504418408fa8a5c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7057f973fa20317158589e772792a3f4abb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b390174f8bf7f848afc416019bf4ea6f1a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha73414b90689f1c8dfdd67f1634454037069;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb91fcd8d9b128789e7604708ed9825529bb9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd2736ab7d0573812091dee32999ab88bfb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d0bcecbb8ad545fdb71f6d4deb57f19a2e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70db7086d8e66221f282b98c3ebde0d4c77a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc15d01d69c671a94791631bfd027534a9d2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2aa295e55a4dba7d220b40a5f3f4e60e2ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha720339e5c6ea81f8dccf609f20417b96ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bd7e102b343f8301b63a44c981bff18f01b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87cb49c6a9ca50e95de68fea600bb678e9df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde05eb65a9c9e7413ec5c9c25eb678c0d4a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc327776448401c3b7186ff675dbd6d9fae9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdede98b535e3a671203f4add5daad4e5128c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0e231fade1b8f0fc98fde96783fd35a398f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha70bce5386d5eb02590d5e59209ae3a1a3b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7580998d2aff66fd89c0dc00698166ddb5b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e59d792b87a7f5bfda1f0ca6f274d9f7270;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6afa342510c9bf476a60b566ebef90b68e4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h448278ea03388ddd28a9e14ff9d9eb413bf2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab874c62aa18acf1fa93f41849590242047a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb3c57e95d3d3102851cfe5c0b2ec9c1463f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19ea0ca6eae91c8498aa4a7917abe0d5dd3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1061ac12c474e47ef18ccfb9c5e969681a20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h445b7ba15e4af11957654e34ae94a51d6e39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h176069ac645ee58259111153476420f2eb1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he63b26479e3ea881de17b464f83bb4884ad2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3a59c2d26e0e533e86da1c91e954b527f63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dc2d07581dd65f71c0ed45432747358c2c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ff52af5d6f964de6b148246bff3d6ddcf42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha18237de3809139201d9d1ddaedcac1cc04f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e1c93a428cef0c7c9c22efb7d79f245460a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a4a5d35e065315980c1fa6e489db0b12d32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h525aaba9b1c659a58cff5aa32f84cff76915;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38a60ce2696aef5878351c9990b6728449a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h526c55dc58844b86add841ce301dece8adbc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he76acd2d9360dd7d89bd59d810e9393635c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h739c6432f0af8abfa18e6f418173ca3cbda2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3e8ec1855212f01628bf313e64942fb1bc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f4651597ee65bd92d937f1f38a66b5cdd5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a0b85c8715c2f82e27daa1f452935a13625;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6773504e287436d588a33569e40e815b9526;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5fc5e7e6492cc009405554948b7dce598478;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ba59be39619f4d54fcefc6475b7e0d65caf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f0dc6bb40eeb16c78d12b6705f0d12c600;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h148068260b8a05fd0ac6160806862b360728;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab1767e96680c0ebd7def70819717f164d51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67eab57f6e95844aa7f9fdd36ca2233e9cd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e4943ee90f726dd24f8fbc72f59d6fd9486;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbd8affcef80bad393e0f0a32e2cad4cccf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94808bc46bffb8f96ed030c3ec22e6fc317b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a01c17c257489ed503ef4447335265f03c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e337170ad5656650231c8fb4115adf7cfb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3672d24989c017a48b5bd7014b08b8248bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6b1a56c13257de96ed1d249d1600f703a37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a9039c46b2cb17706d589d39eeeaf380163;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf1e7938f29542dc1f1dea9338083face58f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75e19cd2736b9ddf78aed281ca034d43ed2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf633b87c5d59277efc00d40538f6705f2d7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6e624374e271fcfae1ae270c1972d6959f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b31a1878c0404e46d369bd5aaf648ff26f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha55d99b4a4fb4cc6e5568ab6f3639b4acee2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd81bbb754591607f21f99ddaadb6ac4d71bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac5db9fcdcd20e67ff4c4c5dccb59a6d3026;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h412d0500a6263f8358c4353a05aaa4256a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c30e09666264f358bb02a7b80c99a3c29ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heda543aaffe3640e0efa1eb493a0b692ef70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h165e818986fab41de33412e39906403325fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ea076eaa4625a185b0e49d7928406401721;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccc44a4a5e7393fe39a8a37a07f1038c77b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h874afa8d10e5d4efbf6edc5ed27b9e0be670;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f5500bf7db47b586a99b285f28de85139e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ba49921fd838be21c989112a7c7d5cfbf34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78cfd7a83d2cd52beee1bab56a3ec485dac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87199f225885fc19c169692f3416baa9ff27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h879efb3b839e8ed0de50799704e1781d4bb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc866c04e73ad9dfe0034eca26473900ef9db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4265afb068f19127447c230836a7491688fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha07e04e5e699a0c17b7df0c96855904d4271;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7f9ab517e3b4162fe598caa69baa9aed42c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbd3393800bfcd36e248e79ac6724e225cdf;
        #1
        $finish();
    end
endmodule
