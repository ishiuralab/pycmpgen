// probclass: mul
// size:      15
// stage:     9
// cost:      31
// elapsed:   7209.145937204361
module compressor (
      input wire [0:0] src0,
      input wire [1:0] src1,
      input wire [2:0] src2,
      input wire [3:0] src3,
      input wire [4:0] src4,
      input wire [5:0] src5,
      input wire [6:0] src6,
      input wire [7:0] src7,
      input wire [8:0] src8,
      input wire [9:0] src9,
      input wire [10:0] src10,
      input wire [11:0] src11,
      input wire [12:0] src12,
      input wire [13:0] src13,
      input wire [14:0] src14,
      input wire [13:0] src15,
      input wire [12:0] src16,
      input wire [11:0] src17,
      input wire [10:0] src18,
      input wire [9:0] src19,
      input wire [8:0] src20,
      input wire [7:0] src21,
      input wire [6:0] src22,
      input wire [5:0] src23,
      input wire [4:0] src24,
      input wire [3:0] src25,
      input wire [2:0] src26,
      input wire [1:0] src27,
      input wire [0:0] src28,
      output wire [0:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [0:0] dst5,
      output wire [0:0] dst6,
      output wire [0:0] dst7,
      output wire [0:0] dst8,
      output wire [0:0] dst9,
      output wire [0:0] dst10,
      output wire [0:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16,
      output wire [0:0] dst17,
      output wire [0:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22,
      output wire [0:0] dst23,
      output wire [0:0] dst24,
      output wire [0:0] dst25,
      output wire [0:0] dst26,
      output wire [0:0] dst27,
      output wire [0:0] dst28,
      output wire [0:0] dst29);

   wire [0:0] stage0_0;
   wire [1:0] stage0_1;
   wire [2:0] stage0_2;
   wire [3:0] stage0_3;
   wire [4:0] stage0_4;
   wire [5:0] stage0_5;
   wire [6:0] stage0_6;
   wire [7:0] stage0_7;
   wire [8:0] stage0_8;
   wire [9:0] stage0_9;
   wire [10:0] stage0_10;
   wire [11:0] stage0_11;
   wire [12:0] stage0_12;
   wire [13:0] stage0_13;
   wire [14:0] stage0_14;
   wire [13:0] stage0_15;
   wire [12:0] stage0_16;
   wire [11:0] stage0_17;
   wire [10:0] stage0_18;
   wire [9:0] stage0_19;
   wire [8:0] stage0_20;
   wire [7:0] stage0_21;
   wire [6:0] stage0_22;
   wire [5:0] stage0_23;
   wire [4:0] stage0_24;
   wire [3:0] stage0_25;
   wire [2:0] stage0_26;
   wire [1:0] stage0_27;
   wire [0:0] stage0_28;
   wire [0:0] stage1_0;
   wire [0:0] stage1_1;
   wire [0:0] stage1_2;
   wire [0:0] stage1_3;
   wire [1:0] stage1_4;
   wire [4:0] stage1_5;
   wire [2:0] stage1_6;
   wire [6:0] stage1_7;
   wire [2:0] stage1_8;
   wire [2:0] stage1_9;
   wire [6:0] stage1_10;
   wire [6:0] stage1_11;
   wire [9:0] stage1_12;
   wire [8:0] stage1_13;
   wire [11:0] stage1_14;
   wire [8:0] stage1_15;
   wire [13:0] stage1_16;
   wire [9:0] stage1_17;
   wire [8:0] stage1_18;
   wire [5:0] stage1_19;
   wire [7:0] stage1_20;
   wire [3:0] stage1_21;
   wire [7:0] stage1_22;
   wire [6:0] stage1_23;
   wire [4:0] stage1_24;
   wire [3:0] stage1_25;
   wire [2:0] stage1_26;
   wire [1:0] stage1_27;
   wire [0:0] stage1_28;
   wire [0:0] stage2_0;
   wire [0:0] stage2_1;
   wire [0:0] stage2_2;
   wire [0:0] stage2_3;
   wire [0:0] stage2_4;
   wire [0:0] stage2_5;
   wire [1:0] stage2_6;
   wire [4:0] stage2_7;
   wire [1:0] stage2_8;
   wire [0:0] stage2_9;
   wire [1:0] stage2_10;
   wire [8:0] stage2_11;
   wire [1:0] stage2_12;
   wire [5:0] stage2_13;
   wire [7:0] stage2_14;
   wire [2:0] stage2_15;
   wire [10:0] stage2_16;
   wire [5:0] stage2_17;
   wire [4:0] stage2_18;
   wire [7:0] stage2_19;
   wire [8:0] stage2_20;
   wire [3:0] stage2_21;
   wire [7:0] stage2_22;
   wire [6:0] stage2_23;
   wire [4:0] stage2_24;
   wire [3:0] stage2_25;
   wire [2:0] stage2_26;
   wire [1:0] stage2_27;
   wire [0:0] stage2_28;
   wire [0:0] stage3_0;
   wire [0:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [0:0] stage3_5;
   wire [0:0] stage3_6;
   wire [0:0] stage3_7;
   wire [0:0] stage3_8;
   wire [0:0] stage3_9;
   wire [2:0] stage3_10;
   wire [4:0] stage3_11;
   wire [1:0] stage3_12;
   wire [0:0] stage3_13;
   wire [3:0] stage3_14;
   wire [4:0] stage3_15;
   wire [5:0] stage3_16;
   wire [6:0] stage3_17;
   wire [1:0] stage3_18;
   wire [7:0] stage3_19;
   wire [3:0] stage3_20;
   wire [4:0] stage3_21;
   wire [8:0] stage3_22;
   wire [6:0] stage3_23;
   wire [4:0] stage3_24;
   wire [3:0] stage3_25;
   wire [2:0] stage3_26;
   wire [1:0] stage3_27;
   wire [0:0] stage3_28;
   wire [0:0] stage4_0;
   wire [0:0] stage4_1;
   wire [0:0] stage4_2;
   wire [0:0] stage4_3;
   wire [0:0] stage4_4;
   wire [0:0] stage4_5;
   wire [0:0] stage4_6;
   wire [0:0] stage4_7;
   wire [0:0] stage4_8;
   wire [0:0] stage4_9;
   wire [0:0] stage4_10;
   wire [0:0] stage4_11;
   wire [0:0] stage4_12;
   wire [0:0] stage4_13;
   wire [4:0] stage4_14;
   wire [0:0] stage4_15;
   wire [5:0] stage4_16;
   wire [1:0] stage4_17;
   wire [2:0] stage4_18;
   wire [2:0] stage4_19;
   wire [4:0] stage4_20;
   wire [3:0] stage4_21;
   wire [9:0] stage4_22;
   wire [6:0] stage4_23;
   wire [4:0] stage4_24;
   wire [3:0] stage4_25;
   wire [2:0] stage4_26;
   wire [1:0] stage4_27;
   wire [0:0] stage4_28;
   wire [0:0] stage5_0;
   wire [0:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [0:0] stage5_4;
   wire [0:0] stage5_5;
   wire [0:0] stage5_6;
   wire [0:0] stage5_7;
   wire [0:0] stage5_8;
   wire [0:0] stage5_9;
   wire [0:0] stage5_10;
   wire [0:0] stage5_11;
   wire [0:0] stage5_12;
   wire [0:0] stage5_13;
   wire [0:0] stage5_14;
   wire [0:0] stage5_15;
   wire [0:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [2:0] stage5_19;
   wire [0:0] stage5_20;
   wire [3:0] stage5_21;
   wire [4:0] stage5_22;
   wire [3:0] stage5_23;
   wire [5:0] stage5_24;
   wire [0:0] stage5_25;
   wire [2:0] stage5_26;
   wire [2:0] stage5_27;
   wire [0:0] stage5_28;
   wire [0:0] stage6_0;
   wire [0:0] stage6_1;
   wire [0:0] stage6_2;
   wire [0:0] stage6_3;
   wire [0:0] stage6_4;
   wire [0:0] stage6_5;
   wire [0:0] stage6_6;
   wire [0:0] stage6_7;
   wire [0:0] stage6_8;
   wire [0:0] stage6_9;
   wire [0:0] stage6_10;
   wire [0:0] stage6_11;
   wire [0:0] stage6_12;
   wire [0:0] stage6_13;
   wire [0:0] stage6_14;
   wire [0:0] stage6_15;
   wire [0:0] stage6_16;
   wire [0:0] stage6_17;
   wire [0:0] stage6_18;
   wire [0:0] stage6_19;
   wire [0:0] stage6_20;
   wire [4:0] stage6_21;
   wire [0:0] stage6_22;
   wire [3:0] stage6_23;
   wire [0:0] stage6_24;
   wire [1:0] stage6_25;
   wire [3:0] stage6_26;
   wire [2:0] stage6_27;
   wire [0:0] stage6_28;
   wire [0:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [0:0] stage7_4;
   wire [0:0] stage7_5;
   wire [0:0] stage7_6;
   wire [0:0] stage7_7;
   wire [0:0] stage7_8;
   wire [0:0] stage7_9;
   wire [0:0] stage7_10;
   wire [0:0] stage7_11;
   wire [0:0] stage7_12;
   wire [0:0] stage7_13;
   wire [0:0] stage7_14;
   wire [0:0] stage7_15;
   wire [0:0] stage7_16;
   wire [0:0] stage7_17;
   wire [0:0] stage7_18;
   wire [0:0] stage7_19;
   wire [0:0] stage7_20;
   wire [0:0] stage7_21;
   wire [0:0] stage7_22;
   wire [0:0] stage7_23;
   wire [0:0] stage7_24;
   wire [2:0] stage7_25;
   wire [3:0] stage7_26;
   wire [2:0] stage7_27;
   wire [0:0] stage7_28;
   wire [0:0] stage8_0;
   wire [0:0] stage8_1;
   wire [0:0] stage8_2;
   wire [0:0] stage8_3;
   wire [0:0] stage8_4;
   wire [0:0] stage8_5;
   wire [0:0] stage8_6;
   wire [0:0] stage8_7;
   wire [0:0] stage8_8;
   wire [0:0] stage8_9;
   wire [0:0] stage8_10;
   wire [0:0] stage8_11;
   wire [0:0] stage8_12;
   wire [0:0] stage8_13;
   wire [0:0] stage8_14;
   wire [0:0] stage8_15;
   wire [0:0] stage8_16;
   wire [0:0] stage8_17;
   wire [0:0] stage8_18;
   wire [0:0] stage8_19;
   wire [0:0] stage8_20;
   wire [0:0] stage8_21;
   wire [0:0] stage8_22;
   wire [0:0] stage8_23;
   wire [0:0] stage8_24;
   wire [0:0] stage8_25;
   wire [0:0] stage8_26;
   wire [0:0] stage8_27;
   wire [0:0] stage8_28;
   wire [0:0] stage8_29;
   wire [0:0] stage9_0;
   wire [0:0] stage9_1;
   wire [0:0] stage9_2;
   wire [0:0] stage9_3;
   wire [0:0] stage9_4;
   wire [0:0] stage9_5;
   wire [0:0] stage9_6;
   wire [0:0] stage9_7;
   wire [0:0] stage9_8;
   wire [0:0] stage9_9;
   wire [0:0] stage9_10;
   wire [0:0] stage9_11;
   wire [0:0] stage9_12;
   wire [0:0] stage9_13;
   wire [0:0] stage9_14;
   wire [0:0] stage9_15;
   wire [0:0] stage9_16;
   wire [0:0] stage9_17;
   wire [0:0] stage9_18;
   wire [0:0] stage9_19;
   wire [0:0] stage9_20;
   wire [0:0] stage9_21;
   wire [0:0] stage9_22;
   wire [0:0] stage9_23;
   wire [0:0] stage9_24;
   wire [0:0] stage9_25;
   wire [0:0] stage9_26;
   wire [0:0] stage9_27;
   wire [0:0] stage9_28;
   wire [0:0] stage9_29;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign dst0 = stage9_0;
   assign dst1 = stage9_1;
   assign dst2 = stage9_2;
   assign dst3 = stage9_3;
   assign dst4 = stage9_4;
   assign dst5 = stage9_5;
   assign dst6 = stage9_6;
   assign dst7 = stage9_7;
   assign dst8 = stage9_8;
   assign dst9 = stage9_9;
   assign dst10 = stage9_10;
   assign dst11 = stage9_11;
   assign dst12 = stage9_12;
   assign dst13 = stage9_13;
   assign dst14 = stage9_14;
   assign dst15 = stage9_15;
   assign dst16 = stage9_16;
   assign dst17 = stage9_17;
   assign dst18 = stage9_18;
   assign dst19 = stage9_19;
   assign dst20 = stage9_20;
   assign dst21 = stage9_21;
   assign dst22 = stage9_22;
   assign dst23 = stage9_23;
   assign dst24 = stage9_24;
   assign dst25 = stage9_25;
   assign dst26 = stage9_26;
   assign dst27 = stage9_27;
   assign dst28 = stage9_28;
   assign dst29 = stage9_29;

   gpc433_5 gpc0 (
      {stage0_1[0], stage0_1[1], 1'b0},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage1_5[0],stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[0],stage1_7[0],stage1_6[0],stage1_5[1],stage1_4[1]}
   );
   gpc615_5 gpc2 (
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage0_7[2]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[0],stage1_8[1],stage1_7[1],stage1_6[1]}
   );
   gpc1253_5 gpc3 (
      {stage0_8[6], stage0_8[7], stage0_8[8]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4]},
      {stage0_10[0], stage0_10[1]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[1],stage1_8[2]}
   );
   gpc615_5 gpc4 (
      {stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_10[2]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[2]}
   );
   gpc615_5 gpc5 (
      {stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[7]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[1],stage1_12[2],stage1_11[2],stage1_10[3]}
   );
   gpc606_5 gpc6 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[0],stage1_15[0],stage1_14[1],stage1_13[2]}
   );
   gpc1163_5 gpc7 (
      {stage0_13[6], stage0_13[7], stage0_13[8]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage0_15[6]},
      {stage0_16[0]},
      {stage1_17[1],stage1_16[1],stage1_15[1],stage1_14[2],stage1_13[3]}
   );
   gpc2135_5 gpc8 (
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4]},
      {stage0_18[0], stage0_18[1], stage0_18[2]},
      {stage0_19[0]},
      {stage0_20[0], stage0_20[1]},
      {stage1_21[0],stage1_20[0],stage1_19[0],stage1_18[0],stage1_17[2]}
   );
   gpc615_5 gpc9 (
      {stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage0_20[2]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[1],stage1_20[1],stage1_19[1]}
   );
   gpc1_1 gpc10 (
      {stage0_0[0]},
      {stage1_0[0]}
   );
   gpc1_1 gpc11 (
      {stage0_5[3]},
      {stage1_5[2]}
   );
   gpc1_1 gpc12 (
      {stage0_5[4]},
      {stage1_5[3]}
   );
   gpc1_1 gpc13 (
      {stage0_5[5]},
      {stage1_5[4]}
   );
   gpc1_1 gpc14 (
      {stage0_6[6]},
      {stage1_6[2]}
   );
   gpc1_1 gpc15 (
      {stage0_7[3]},
      {stage1_7[2]}
   );
   gpc1_1 gpc16 (
      {stage0_7[4]},
      {stage1_7[3]}
   );
   gpc1_1 gpc17 (
      {stage0_7[5]},
      {stage1_7[4]}
   );
   gpc1_1 gpc18 (
      {stage0_7[6]},
      {stage1_7[5]}
   );
   gpc1_1 gpc19 (
      {stage0_7[7]},
      {stage1_7[6]}
   );
   gpc1_1 gpc20 (
      {stage0_10[8]},
      {stage1_10[4]}
   );
   gpc1_1 gpc21 (
      {stage0_10[9]},
      {stage1_10[5]}
   );
   gpc1_1 gpc22 (
      {stage0_10[10]},
      {stage1_10[6]}
   );
   gpc1_1 gpc23 (
      {stage0_11[8]},
      {stage1_11[3]}
   );
   gpc1_1 gpc24 (
      {stage0_11[9]},
      {stage1_11[4]}
   );
   gpc1_1 gpc25 (
      {stage0_11[10]},
      {stage1_11[5]}
   );
   gpc1_1 gpc26 (
      {stage0_11[11]},
      {stage1_11[6]}
   );
   gpc1_1 gpc27 (
      {stage0_12[6]},
      {stage1_12[3]}
   );
   gpc1_1 gpc28 (
      {stage0_12[7]},
      {stage1_12[4]}
   );
   gpc1_1 gpc29 (
      {stage0_12[8]},
      {stage1_12[5]}
   );
   gpc1_1 gpc30 (
      {stage0_12[9]},
      {stage1_12[6]}
   );
   gpc1_1 gpc31 (
      {stage0_12[10]},
      {stage1_12[7]}
   );
   gpc1_1 gpc32 (
      {stage0_12[11]},
      {stage1_12[8]}
   );
   gpc1_1 gpc33 (
      {stage0_12[12]},
      {stage1_12[9]}
   );
   gpc1_1 gpc34 (
      {stage0_13[9]},
      {stage1_13[4]}
   );
   gpc1_1 gpc35 (
      {stage0_13[10]},
      {stage1_13[5]}
   );
   gpc1_1 gpc36 (
      {stage0_13[11]},
      {stage1_13[6]}
   );
   gpc1_1 gpc37 (
      {stage0_13[12]},
      {stage1_13[7]}
   );
   gpc1_1 gpc38 (
      {stage0_13[13]},
      {stage1_13[8]}
   );
   gpc1_1 gpc39 (
      {stage0_14[6]},
      {stage1_14[3]}
   );
   gpc1_1 gpc40 (
      {stage0_14[7]},
      {stage1_14[4]}
   );
   gpc1_1 gpc41 (
      {stage0_14[8]},
      {stage1_14[5]}
   );
   gpc1_1 gpc42 (
      {stage0_14[9]},
      {stage1_14[6]}
   );
   gpc1_1 gpc43 (
      {stage0_14[10]},
      {stage1_14[7]}
   );
   gpc1_1 gpc44 (
      {stage0_14[11]},
      {stage1_14[8]}
   );
   gpc1_1 gpc45 (
      {stage0_14[12]},
      {stage1_14[9]}
   );
   gpc1_1 gpc46 (
      {stage0_14[13]},
      {stage1_14[10]}
   );
   gpc1_1 gpc47 (
      {stage0_14[14]},
      {stage1_14[11]}
   );
   gpc1_1 gpc48 (
      {stage0_15[7]},
      {stage1_15[2]}
   );
   gpc1_1 gpc49 (
      {stage0_15[8]},
      {stage1_15[3]}
   );
   gpc1_1 gpc50 (
      {stage0_15[9]},
      {stage1_15[4]}
   );
   gpc1_1 gpc51 (
      {stage0_15[10]},
      {stage1_15[5]}
   );
   gpc1_1 gpc52 (
      {stage0_15[11]},
      {stage1_15[6]}
   );
   gpc1_1 gpc53 (
      {stage0_15[12]},
      {stage1_15[7]}
   );
   gpc1_1 gpc54 (
      {stage0_15[13]},
      {stage1_15[8]}
   );
   gpc1_1 gpc55 (
      {stage0_16[1]},
      {stage1_16[2]}
   );
   gpc1_1 gpc56 (
      {stage0_16[2]},
      {stage1_16[3]}
   );
   gpc1_1 gpc57 (
      {stage0_16[3]},
      {stage1_16[4]}
   );
   gpc1_1 gpc58 (
      {stage0_16[4]},
      {stage1_16[5]}
   );
   gpc1_1 gpc59 (
      {stage0_16[5]},
      {stage1_16[6]}
   );
   gpc1_1 gpc60 (
      {stage0_16[6]},
      {stage1_16[7]}
   );
   gpc1_1 gpc61 (
      {stage0_16[7]},
      {stage1_16[8]}
   );
   gpc1_1 gpc62 (
      {stage0_16[8]},
      {stage1_16[9]}
   );
   gpc1_1 gpc63 (
      {stage0_16[9]},
      {stage1_16[10]}
   );
   gpc1_1 gpc64 (
      {stage0_16[10]},
      {stage1_16[11]}
   );
   gpc1_1 gpc65 (
      {stage0_16[11]},
      {stage1_16[12]}
   );
   gpc1_1 gpc66 (
      {stage0_16[12]},
      {stage1_16[13]}
   );
   gpc1_1 gpc67 (
      {stage0_17[5]},
      {stage1_17[3]}
   );
   gpc1_1 gpc68 (
      {stage0_17[6]},
      {stage1_17[4]}
   );
   gpc1_1 gpc69 (
      {stage0_17[7]},
      {stage1_17[5]}
   );
   gpc1_1 gpc70 (
      {stage0_17[8]},
      {stage1_17[6]}
   );
   gpc1_1 gpc71 (
      {stage0_17[9]},
      {stage1_17[7]}
   );
   gpc1_1 gpc72 (
      {stage0_17[10]},
      {stage1_17[8]}
   );
   gpc1_1 gpc73 (
      {stage0_17[11]},
      {stage1_17[9]}
   );
   gpc1_1 gpc74 (
      {stage0_18[3]},
      {stage1_18[1]}
   );
   gpc1_1 gpc75 (
      {stage0_18[4]},
      {stage1_18[2]}
   );
   gpc1_1 gpc76 (
      {stage0_18[5]},
      {stage1_18[3]}
   );
   gpc1_1 gpc77 (
      {stage0_18[6]},
      {stage1_18[4]}
   );
   gpc1_1 gpc78 (
      {stage0_18[7]},
      {stage1_18[5]}
   );
   gpc1_1 gpc79 (
      {stage0_18[8]},
      {stage1_18[6]}
   );
   gpc1_1 gpc80 (
      {stage0_18[9]},
      {stage1_18[7]}
   );
   gpc1_1 gpc81 (
      {stage0_18[10]},
      {stage1_18[8]}
   );
   gpc1_1 gpc82 (
      {stage0_19[6]},
      {stage1_19[2]}
   );
   gpc1_1 gpc83 (
      {stage0_19[7]},
      {stage1_19[3]}
   );
   gpc1_1 gpc84 (
      {stage0_19[8]},
      {stage1_19[4]}
   );
   gpc1_1 gpc85 (
      {stage0_19[9]},
      {stage1_19[5]}
   );
   gpc1_1 gpc86 (
      {stage0_20[3]},
      {stage1_20[2]}
   );
   gpc1_1 gpc87 (
      {stage0_20[4]},
      {stage1_20[3]}
   );
   gpc1_1 gpc88 (
      {stage0_20[5]},
      {stage1_20[4]}
   );
   gpc1_1 gpc89 (
      {stage0_20[6]},
      {stage1_20[5]}
   );
   gpc1_1 gpc90 (
      {stage0_20[7]},
      {stage1_20[6]}
   );
   gpc1_1 gpc91 (
      {stage0_20[8]},
      {stage1_20[7]}
   );
   gpc1_1 gpc92 (
      {stage0_21[6]},
      {stage1_21[2]}
   );
   gpc1_1 gpc93 (
      {stage0_21[7]},
      {stage1_21[3]}
   );
   gpc1_1 gpc94 (
      {stage0_22[0]},
      {stage1_22[1]}
   );
   gpc1_1 gpc95 (
      {stage0_22[1]},
      {stage1_22[2]}
   );
   gpc1_1 gpc96 (
      {stage0_22[2]},
      {stage1_22[3]}
   );
   gpc1_1 gpc97 (
      {stage0_22[3]},
      {stage1_22[4]}
   );
   gpc1_1 gpc98 (
      {stage0_22[4]},
      {stage1_22[5]}
   );
   gpc1_1 gpc99 (
      {stage0_22[5]},
      {stage1_22[6]}
   );
   gpc1_1 gpc100 (
      {stage0_22[6]},
      {stage1_22[7]}
   );
   gpc1_1 gpc101 (
      {stage0_23[0]},
      {stage1_23[1]}
   );
   gpc1_1 gpc102 (
      {stage0_23[1]},
      {stage1_23[2]}
   );
   gpc1_1 gpc103 (
      {stage0_23[2]},
      {stage1_23[3]}
   );
   gpc1_1 gpc104 (
      {stage0_23[3]},
      {stage1_23[4]}
   );
   gpc1_1 gpc105 (
      {stage0_23[4]},
      {stage1_23[5]}
   );
   gpc1_1 gpc106 (
      {stage0_23[5]},
      {stage1_23[6]}
   );
   gpc1_1 gpc107 (
      {stage0_24[0]},
      {stage1_24[0]}
   );
   gpc1_1 gpc108 (
      {stage0_24[1]},
      {stage1_24[1]}
   );
   gpc1_1 gpc109 (
      {stage0_24[2]},
      {stage1_24[2]}
   );
   gpc1_1 gpc110 (
      {stage0_24[3]},
      {stage1_24[3]}
   );
   gpc1_1 gpc111 (
      {stage0_24[4]},
      {stage1_24[4]}
   );
   gpc1_1 gpc112 (
      {stage0_25[0]},
      {stage1_25[0]}
   );
   gpc1_1 gpc113 (
      {stage0_25[1]},
      {stage1_25[1]}
   );
   gpc1_1 gpc114 (
      {stage0_25[2]},
      {stage1_25[2]}
   );
   gpc1_1 gpc115 (
      {stage0_25[3]},
      {stage1_25[3]}
   );
   gpc1_1 gpc116 (
      {stage0_26[0]},
      {stage1_26[0]}
   );
   gpc1_1 gpc117 (
      {stage0_26[1]},
      {stage1_26[1]}
   );
   gpc1_1 gpc118 (
      {stage0_26[2]},
      {stage1_26[2]}
   );
   gpc1_1 gpc119 (
      {stage0_27[0]},
      {stage1_27[0]}
   );
   gpc1_1 gpc120 (
      {stage0_27[1]},
      {stage1_27[1]}
   );
   gpc1_1 gpc121 (
      {stage0_28[0]},
      {stage1_28[0]}
   );
   gpc1253_5 gpc122 (
      {stage1_4[0], stage1_4[1], 1'b0},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4]},
      {stage1_6[0], stage1_6[1]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[0]}
   );
   gpc1343_5 gpc123 (
      {stage1_7[1], stage1_7[2], stage1_7[3]},
      {stage1_8[0], stage1_8[1], stage1_8[2], 1'b0},
      {stage1_9[0], stage1_9[1], stage1_9[2]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[0],stage2_9[0],stage2_8[1],stage2_7[1]}
   );
   gpc606_5 gpc124 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[0],stage2_11[1],stage2_10[1]}
   );
   gpc615_5 gpc125 (
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], 1'b0},
      {stage1_13[0]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[1]}
   );
   gpc1415_5 gpc126 (
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_14[6]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3]},
      {stage1_16[0]},
      {stage2_17[0],stage2_16[1],stage2_15[1],stage2_14[2],stage2_13[2]}
   );
   gpc615_5 gpc127 (
      {stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], stage1_15[8]},
      {stage1_16[1]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[2],stage2_15[2]}
   );
   gpc615_5 gpc128 (
      {stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[6]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[3]}
   );
   gpc1_1 gpc129 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc130 (
      {stage1_1[0]},
      {stage2_1[0]}
   );
   gpc1_1 gpc131 (
      {stage1_2[0]},
      {stage2_2[0]}
   );
   gpc1_1 gpc132 (
      {stage1_3[0]},
      {stage2_3[0]}
   );
   gpc1_1 gpc133 (
      {stage1_6[2]},
      {stage2_6[1]}
   );
   gpc1_1 gpc134 (
      {stage1_7[4]},
      {stage2_7[2]}
   );
   gpc1_1 gpc135 (
      {stage1_7[5]},
      {stage2_7[3]}
   );
   gpc1_1 gpc136 (
      {stage1_7[6]},
      {stage2_7[4]}
   );
   gpc1_1 gpc137 (
      {stage1_11[0]},
      {stage2_11[2]}
   );
   gpc1_1 gpc138 (
      {stage1_11[1]},
      {stage2_11[3]}
   );
   gpc1_1 gpc139 (
      {stage1_11[2]},
      {stage2_11[4]}
   );
   gpc1_1 gpc140 (
      {stage1_11[3]},
      {stage2_11[5]}
   );
   gpc1_1 gpc141 (
      {stage1_11[4]},
      {stage2_11[6]}
   );
   gpc1_1 gpc142 (
      {stage1_11[5]},
      {stage2_11[7]}
   );
   gpc1_1 gpc143 (
      {stage1_11[6]},
      {stage2_11[8]}
   );
   gpc1_1 gpc144 (
      {stage1_13[6]},
      {stage2_13[3]}
   );
   gpc1_1 gpc145 (
      {stage1_13[7]},
      {stage2_13[4]}
   );
   gpc1_1 gpc146 (
      {stage1_13[8]},
      {stage2_13[5]}
   );
   gpc1_1 gpc147 (
      {stage1_14[7]},
      {stage2_14[3]}
   );
   gpc1_1 gpc148 (
      {stage1_14[8]},
      {stage2_14[4]}
   );
   gpc1_1 gpc149 (
      {stage1_14[9]},
      {stage2_14[5]}
   );
   gpc1_1 gpc150 (
      {stage1_14[10]},
      {stage2_14[6]}
   );
   gpc1_1 gpc151 (
      {stage1_14[11]},
      {stage2_14[7]}
   );
   gpc1_1 gpc152 (
      {stage1_16[7]},
      {stage2_16[4]}
   );
   gpc1_1 gpc153 (
      {stage1_16[8]},
      {stage2_16[5]}
   );
   gpc1_1 gpc154 (
      {stage1_16[9]},
      {stage2_16[6]}
   );
   gpc1_1 gpc155 (
      {stage1_16[10]},
      {stage2_16[7]}
   );
   gpc1_1 gpc156 (
      {stage1_16[11]},
      {stage2_16[8]}
   );
   gpc1_1 gpc157 (
      {stage1_16[12]},
      {stage2_16[9]}
   );
   gpc1_1 gpc158 (
      {stage1_16[13]},
      {stage2_16[10]}
   );
   gpc1_1 gpc159 (
      {stage1_17[7]},
      {stage2_17[3]}
   );
   gpc1_1 gpc160 (
      {stage1_17[8]},
      {stage2_17[4]}
   );
   gpc1_1 gpc161 (
      {stage1_17[9]},
      {stage2_17[5]}
   );
   gpc1_1 gpc162 (
      {stage1_18[6]},
      {stage2_18[2]}
   );
   gpc1_1 gpc163 (
      {stage1_18[7]},
      {stage2_18[3]}
   );
   gpc1_1 gpc164 (
      {stage1_18[8]},
      {stage2_18[4]}
   );
   gpc1_1 gpc165 (
      {stage1_19[0]},
      {stage2_19[2]}
   );
   gpc1_1 gpc166 (
      {stage1_19[1]},
      {stage2_19[3]}
   );
   gpc1_1 gpc167 (
      {stage1_19[2]},
      {stage2_19[4]}
   );
   gpc1_1 gpc168 (
      {stage1_19[3]},
      {stage2_19[5]}
   );
   gpc1_1 gpc169 (
      {stage1_19[4]},
      {stage2_19[6]}
   );
   gpc1_1 gpc170 (
      {stage1_19[5]},
      {stage2_19[7]}
   );
   gpc1_1 gpc171 (
      {stage1_20[0]},
      {stage2_20[1]}
   );
   gpc1_1 gpc172 (
      {stage1_20[1]},
      {stage2_20[2]}
   );
   gpc1_1 gpc173 (
      {stage1_20[2]},
      {stage2_20[3]}
   );
   gpc1_1 gpc174 (
      {stage1_20[3]},
      {stage2_20[4]}
   );
   gpc1_1 gpc175 (
      {stage1_20[4]},
      {stage2_20[5]}
   );
   gpc1_1 gpc176 (
      {stage1_20[5]},
      {stage2_20[6]}
   );
   gpc1_1 gpc177 (
      {stage1_20[6]},
      {stage2_20[7]}
   );
   gpc1_1 gpc178 (
      {stage1_20[7]},
      {stage2_20[8]}
   );
   gpc1_1 gpc179 (
      {stage1_21[0]},
      {stage2_21[0]}
   );
   gpc1_1 gpc180 (
      {stage1_21[1]},
      {stage2_21[1]}
   );
   gpc1_1 gpc181 (
      {stage1_21[2]},
      {stage2_21[2]}
   );
   gpc1_1 gpc182 (
      {stage1_21[3]},
      {stage2_21[3]}
   );
   gpc1_1 gpc183 (
      {stage1_22[0]},
      {stage2_22[0]}
   );
   gpc1_1 gpc184 (
      {stage1_22[1]},
      {stage2_22[1]}
   );
   gpc1_1 gpc185 (
      {stage1_22[2]},
      {stage2_22[2]}
   );
   gpc1_1 gpc186 (
      {stage1_22[3]},
      {stage2_22[3]}
   );
   gpc1_1 gpc187 (
      {stage1_22[4]},
      {stage2_22[4]}
   );
   gpc1_1 gpc188 (
      {stage1_22[5]},
      {stage2_22[5]}
   );
   gpc1_1 gpc189 (
      {stage1_22[6]},
      {stage2_22[6]}
   );
   gpc1_1 gpc190 (
      {stage1_22[7]},
      {stage2_22[7]}
   );
   gpc1_1 gpc191 (
      {stage1_23[0]},
      {stage2_23[0]}
   );
   gpc1_1 gpc192 (
      {stage1_23[1]},
      {stage2_23[1]}
   );
   gpc1_1 gpc193 (
      {stage1_23[2]},
      {stage2_23[2]}
   );
   gpc1_1 gpc194 (
      {stage1_23[3]},
      {stage2_23[3]}
   );
   gpc1_1 gpc195 (
      {stage1_23[4]},
      {stage2_23[4]}
   );
   gpc1_1 gpc196 (
      {stage1_23[5]},
      {stage2_23[5]}
   );
   gpc1_1 gpc197 (
      {stage1_23[6]},
      {stage2_23[6]}
   );
   gpc1_1 gpc198 (
      {stage1_24[0]},
      {stage2_24[0]}
   );
   gpc1_1 gpc199 (
      {stage1_24[1]},
      {stage2_24[1]}
   );
   gpc1_1 gpc200 (
      {stage1_24[2]},
      {stage2_24[2]}
   );
   gpc1_1 gpc201 (
      {stage1_24[3]},
      {stage2_24[3]}
   );
   gpc1_1 gpc202 (
      {stage1_24[4]},
      {stage2_24[4]}
   );
   gpc1_1 gpc203 (
      {stage1_25[0]},
      {stage2_25[0]}
   );
   gpc1_1 gpc204 (
      {stage1_25[1]},
      {stage2_25[1]}
   );
   gpc1_1 gpc205 (
      {stage1_25[2]},
      {stage2_25[2]}
   );
   gpc1_1 gpc206 (
      {stage1_25[3]},
      {stage2_25[3]}
   );
   gpc1_1 gpc207 (
      {stage1_26[0]},
      {stage2_26[0]}
   );
   gpc1_1 gpc208 (
      {stage1_26[1]},
      {stage2_26[1]}
   );
   gpc1_1 gpc209 (
      {stage1_26[2]},
      {stage2_26[2]}
   );
   gpc1_1 gpc210 (
      {stage1_27[0]},
      {stage2_27[0]}
   );
   gpc1_1 gpc211 (
      {stage1_27[1]},
      {stage2_27[1]}
   );
   gpc1_1 gpc212 (
      {stage1_28[0]},
      {stage2_28[0]}
   );
   gpc1253_5 gpc213 (
      {stage2_6[0], stage2_6[1], 1'b0},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0], stage2_8[1]},
      {stage2_9[0]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[0]}
   );
   gpc615_5 gpc214 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[0]}
   );
   gpc606_5 gpc215 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[0],stage3_15[1],stage3_14[1]}
   );
   gpc615_5 gpc216 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[0]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[1]}
   );
   gpc1_1 gpc217 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc218 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc219 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc220 (
      {stage2_3[0]},
      {stage3_3[0]}
   );
   gpc1_1 gpc221 (
      {stage2_4[0]},
      {stage3_4[0]}
   );
   gpc1_1 gpc222 (
      {stage2_5[0]},
      {stage3_5[0]}
   );
   gpc1_1 gpc223 (
      {stage2_10[0]},
      {stage3_10[1]}
   );
   gpc1_1 gpc224 (
      {stage2_10[1]},
      {stage3_10[2]}
   );
   gpc1_1 gpc225 (
      {stage2_11[5]},
      {stage3_11[1]}
   );
   gpc1_1 gpc226 (
      {stage2_11[6]},
      {stage3_11[2]}
   );
   gpc1_1 gpc227 (
      {stage2_11[7]},
      {stage3_11[3]}
   );
   gpc1_1 gpc228 (
      {stage2_11[8]},
      {stage3_11[4]}
   );
   gpc1_1 gpc229 (
      {stage2_12[1]},
      {stage3_12[1]}
   );
   gpc1_1 gpc230 (
      {stage2_14[6]},
      {stage3_14[2]}
   );
   gpc1_1 gpc231 (
      {stage2_14[7]},
      {stage3_14[3]}
   );
   gpc1_1 gpc232 (
      {stage2_15[0]},
      {stage3_15[2]}
   );
   gpc1_1 gpc233 (
      {stage2_15[1]},
      {stage3_15[3]}
   );
   gpc1_1 gpc234 (
      {stage2_15[2]},
      {stage3_15[4]}
   );
   gpc1_1 gpc235 (
      {stage2_16[6]},
      {stage3_16[1]}
   );
   gpc1_1 gpc236 (
      {stage2_16[7]},
      {stage3_16[2]}
   );
   gpc1_1 gpc237 (
      {stage2_16[8]},
      {stage3_16[3]}
   );
   gpc1_1 gpc238 (
      {stage2_16[9]},
      {stage3_16[4]}
   );
   gpc1_1 gpc239 (
      {stage2_16[10]},
      {stage3_16[5]}
   );
   gpc1_1 gpc240 (
      {stage2_17[0]},
      {stage3_17[1]}
   );
   gpc1_1 gpc241 (
      {stage2_17[1]},
      {stage3_17[2]}
   );
   gpc1_1 gpc242 (
      {stage2_17[2]},
      {stage3_17[3]}
   );
   gpc1_1 gpc243 (
      {stage2_17[3]},
      {stage3_17[4]}
   );
   gpc1_1 gpc244 (
      {stage2_17[4]},
      {stage3_17[5]}
   );
   gpc1_1 gpc245 (
      {stage2_17[5]},
      {stage3_17[6]}
   );
   gpc1_1 gpc246 (
      {stage2_19[1]},
      {stage3_19[1]}
   );
   gpc1_1 gpc247 (
      {stage2_19[2]},
      {stage3_19[2]}
   );
   gpc1_1 gpc248 (
      {stage2_19[3]},
      {stage3_19[3]}
   );
   gpc1_1 gpc249 (
      {stage2_19[4]},
      {stage3_19[4]}
   );
   gpc1_1 gpc250 (
      {stage2_19[5]},
      {stage3_19[5]}
   );
   gpc1_1 gpc251 (
      {stage2_19[6]},
      {stage3_19[6]}
   );
   gpc1_1 gpc252 (
      {stage2_19[7]},
      {stage3_19[7]}
   );
   gpc1_1 gpc253 (
      {stage2_20[6]},
      {stage3_20[1]}
   );
   gpc1_1 gpc254 (
      {stage2_20[7]},
      {stage3_20[2]}
   );
   gpc1_1 gpc255 (
      {stage2_20[8]},
      {stage3_20[3]}
   );
   gpc1_1 gpc256 (
      {stage2_21[0]},
      {stage3_21[1]}
   );
   gpc1_1 gpc257 (
      {stage2_21[1]},
      {stage3_21[2]}
   );
   gpc1_1 gpc258 (
      {stage2_21[2]},
      {stage3_21[3]}
   );
   gpc1_1 gpc259 (
      {stage2_21[3]},
      {stage3_21[4]}
   );
   gpc1_1 gpc260 (
      {stage2_22[0]},
      {stage3_22[1]}
   );
   gpc1_1 gpc261 (
      {stage2_22[1]},
      {stage3_22[2]}
   );
   gpc1_1 gpc262 (
      {stage2_22[2]},
      {stage3_22[3]}
   );
   gpc1_1 gpc263 (
      {stage2_22[3]},
      {stage3_22[4]}
   );
   gpc1_1 gpc264 (
      {stage2_22[4]},
      {stage3_22[5]}
   );
   gpc1_1 gpc265 (
      {stage2_22[5]},
      {stage3_22[6]}
   );
   gpc1_1 gpc266 (
      {stage2_22[6]},
      {stage3_22[7]}
   );
   gpc1_1 gpc267 (
      {stage2_22[7]},
      {stage3_22[8]}
   );
   gpc1_1 gpc268 (
      {stage2_23[0]},
      {stage3_23[0]}
   );
   gpc1_1 gpc269 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc270 (
      {stage2_23[2]},
      {stage3_23[2]}
   );
   gpc1_1 gpc271 (
      {stage2_23[3]},
      {stage3_23[3]}
   );
   gpc1_1 gpc272 (
      {stage2_23[4]},
      {stage3_23[4]}
   );
   gpc1_1 gpc273 (
      {stage2_23[5]},
      {stage3_23[5]}
   );
   gpc1_1 gpc274 (
      {stage2_23[6]},
      {stage3_23[6]}
   );
   gpc1_1 gpc275 (
      {stage2_24[0]},
      {stage3_24[0]}
   );
   gpc1_1 gpc276 (
      {stage2_24[1]},
      {stage3_24[1]}
   );
   gpc1_1 gpc277 (
      {stage2_24[2]},
      {stage3_24[2]}
   );
   gpc1_1 gpc278 (
      {stage2_24[3]},
      {stage3_24[3]}
   );
   gpc1_1 gpc279 (
      {stage2_24[4]},
      {stage3_24[4]}
   );
   gpc1_1 gpc280 (
      {stage2_25[0]},
      {stage3_25[0]}
   );
   gpc1_1 gpc281 (
      {stage2_25[1]},
      {stage3_25[1]}
   );
   gpc1_1 gpc282 (
      {stage2_25[2]},
      {stage3_25[2]}
   );
   gpc1_1 gpc283 (
      {stage2_25[3]},
      {stage3_25[3]}
   );
   gpc1_1 gpc284 (
      {stage2_26[0]},
      {stage3_26[0]}
   );
   gpc1_1 gpc285 (
      {stage2_26[1]},
      {stage3_26[1]}
   );
   gpc1_1 gpc286 (
      {stage2_26[2]},
      {stage3_26[2]}
   );
   gpc1_1 gpc287 (
      {stage2_27[0]},
      {stage3_27[0]}
   );
   gpc1_1 gpc288 (
      {stage2_27[1]},
      {stage3_27[1]}
   );
   gpc1_1 gpc289 (
      {stage2_28[0]},
      {stage3_28[0]}
   );
   gpc1253_5 gpc290 (
      {stage3_10[0], stage3_10[1], stage3_10[2]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4]},
      {stage3_12[0], stage3_12[1]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[0]}
   );
   gpc615_5 gpc291 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[0]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[0]}
   );
   gpc207_4 gpc292 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_21[0], stage3_21[1]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[1]}
   );
   gpc1_1 gpc293 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc294 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc295 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc296 (
      {stage3_3[0]},
      {stage4_3[0]}
   );
   gpc1_1 gpc297 (
      {stage3_4[0]},
      {stage4_4[0]}
   );
   gpc1_1 gpc298 (
      {stage3_5[0]},
      {stage4_5[0]}
   );
   gpc1_1 gpc299 (
      {stage3_6[0]},
      {stage4_6[0]}
   );
   gpc1_1 gpc300 (
      {stage3_7[0]},
      {stage4_7[0]}
   );
   gpc1_1 gpc301 (
      {stage3_8[0]},
      {stage4_8[0]}
   );
   gpc1_1 gpc302 (
      {stage3_9[0]},
      {stage4_9[0]}
   );
   gpc1_1 gpc303 (
      {stage3_14[0]},
      {stage4_14[1]}
   );
   gpc1_1 gpc304 (
      {stage3_14[1]},
      {stage4_14[2]}
   );
   gpc1_1 gpc305 (
      {stage3_14[2]},
      {stage4_14[3]}
   );
   gpc1_1 gpc306 (
      {stage3_14[3]},
      {stage4_14[4]}
   );
   gpc1_1 gpc307 (
      {stage3_16[1]},
      {stage4_16[1]}
   );
   gpc1_1 gpc308 (
      {stage3_16[2]},
      {stage4_16[2]}
   );
   gpc1_1 gpc309 (
      {stage3_16[3]},
      {stage4_16[3]}
   );
   gpc1_1 gpc310 (
      {stage3_16[4]},
      {stage4_16[4]}
   );
   gpc1_1 gpc311 (
      {stage3_16[5]},
      {stage4_16[5]}
   );
   gpc1_1 gpc312 (
      {stage3_17[6]},
      {stage4_17[1]}
   );
   gpc1_1 gpc313 (
      {stage3_18[0]},
      {stage4_18[1]}
   );
   gpc1_1 gpc314 (
      {stage3_18[1]},
      {stage4_18[2]}
   );
   gpc1_1 gpc315 (
      {stage3_19[7]},
      {stage4_19[2]}
   );
   gpc1_1 gpc316 (
      {stage3_20[0]},
      {stage4_20[1]}
   );
   gpc1_1 gpc317 (
      {stage3_20[1]},
      {stage4_20[2]}
   );
   gpc1_1 gpc318 (
      {stage3_20[2]},
      {stage4_20[3]}
   );
   gpc1_1 gpc319 (
      {stage3_20[3]},
      {stage4_20[4]}
   );
   gpc1_1 gpc320 (
      {stage3_21[2]},
      {stage4_21[1]}
   );
   gpc1_1 gpc321 (
      {stage3_21[3]},
      {stage4_21[2]}
   );
   gpc1_1 gpc322 (
      {stage3_21[4]},
      {stage4_21[3]}
   );
   gpc1_1 gpc323 (
      {stage3_22[0]},
      {stage4_22[1]}
   );
   gpc1_1 gpc324 (
      {stage3_22[1]},
      {stage4_22[2]}
   );
   gpc1_1 gpc325 (
      {stage3_22[2]},
      {stage4_22[3]}
   );
   gpc1_1 gpc326 (
      {stage3_22[3]},
      {stage4_22[4]}
   );
   gpc1_1 gpc327 (
      {stage3_22[4]},
      {stage4_22[5]}
   );
   gpc1_1 gpc328 (
      {stage3_22[5]},
      {stage4_22[6]}
   );
   gpc1_1 gpc329 (
      {stage3_22[6]},
      {stage4_22[7]}
   );
   gpc1_1 gpc330 (
      {stage3_22[7]},
      {stage4_22[8]}
   );
   gpc1_1 gpc331 (
      {stage3_22[8]},
      {stage4_22[9]}
   );
   gpc1_1 gpc332 (
      {stage3_23[0]},
      {stage4_23[0]}
   );
   gpc1_1 gpc333 (
      {stage3_23[1]},
      {stage4_23[1]}
   );
   gpc1_1 gpc334 (
      {stage3_23[2]},
      {stage4_23[2]}
   );
   gpc1_1 gpc335 (
      {stage3_23[3]},
      {stage4_23[3]}
   );
   gpc1_1 gpc336 (
      {stage3_23[4]},
      {stage4_23[4]}
   );
   gpc1_1 gpc337 (
      {stage3_23[5]},
      {stage4_23[5]}
   );
   gpc1_1 gpc338 (
      {stage3_23[6]},
      {stage4_23[6]}
   );
   gpc1_1 gpc339 (
      {stage3_24[0]},
      {stage4_24[0]}
   );
   gpc1_1 gpc340 (
      {stage3_24[1]},
      {stage4_24[1]}
   );
   gpc1_1 gpc341 (
      {stage3_24[2]},
      {stage4_24[2]}
   );
   gpc1_1 gpc342 (
      {stage3_24[3]},
      {stage4_24[3]}
   );
   gpc1_1 gpc343 (
      {stage3_24[4]},
      {stage4_24[4]}
   );
   gpc1_1 gpc344 (
      {stage3_25[0]},
      {stage4_25[0]}
   );
   gpc1_1 gpc345 (
      {stage3_25[1]},
      {stage4_25[1]}
   );
   gpc1_1 gpc346 (
      {stage3_25[2]},
      {stage4_25[2]}
   );
   gpc1_1 gpc347 (
      {stage3_25[3]},
      {stage4_25[3]}
   );
   gpc1_1 gpc348 (
      {stage3_26[0]},
      {stage4_26[0]}
   );
   gpc1_1 gpc349 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
   gpc1_1 gpc350 (
      {stage3_26[2]},
      {stage4_26[2]}
   );
   gpc1_1 gpc351 (
      {stage3_27[0]},
      {stage4_27[0]}
   );
   gpc1_1 gpc352 (
      {stage3_27[1]},
      {stage4_27[1]}
   );
   gpc1_1 gpc353 (
      {stage3_28[0]},
      {stage4_28[0]}
   );
   gpc615_5 gpc354 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0]}
   );
   gpc615_5 gpc355 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4]},
      {stage4_21[0]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[0]}
   );
   gpc1415_5 gpc356 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4]},
      {stage4_24[0]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[1]}
   );
   gpc1_1 gpc357 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc358 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc359 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc360 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc361 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc362 (
      {stage4_5[0]},
      {stage5_5[0]}
   );
   gpc1_1 gpc363 (
      {stage4_6[0]},
      {stage5_6[0]}
   );
   gpc1_1 gpc364 (
      {stage4_7[0]},
      {stage5_7[0]}
   );
   gpc1_1 gpc365 (
      {stage4_8[0]},
      {stage5_8[0]}
   );
   gpc1_1 gpc366 (
      {stage4_9[0]},
      {stage5_9[0]}
   );
   gpc1_1 gpc367 (
      {stage4_10[0]},
      {stage5_10[0]}
   );
   gpc1_1 gpc368 (
      {stage4_11[0]},
      {stage5_11[0]}
   );
   gpc1_1 gpc369 (
      {stage4_12[0]},
      {stage5_12[0]}
   );
   gpc1_1 gpc370 (
      {stage4_13[0]},
      {stage5_13[0]}
   );
   gpc1_1 gpc371 (
      {stage4_17[0]},
      {stage5_17[1]}
   );
   gpc1_1 gpc372 (
      {stage4_17[1]},
      {stage5_17[2]}
   );
   gpc1_1 gpc373 (
      {stage4_18[0]},
      {stage5_18[1]}
   );
   gpc1_1 gpc374 (
      {stage4_18[1]},
      {stage5_18[2]}
   );
   gpc1_1 gpc375 (
      {stage4_18[2]},
      {stage5_18[3]}
   );
   gpc1_1 gpc376 (
      {stage4_19[0]},
      {stage5_19[0]}
   );
   gpc1_1 gpc377 (
      {stage4_19[1]},
      {stage5_19[1]}
   );
   gpc1_1 gpc378 (
      {stage4_19[2]},
      {stage5_19[2]}
   );
   gpc1_1 gpc379 (
      {stage4_21[1]},
      {stage5_21[1]}
   );
   gpc1_1 gpc380 (
      {stage4_21[2]},
      {stage5_21[2]}
   );
   gpc1_1 gpc381 (
      {stage4_21[3]},
      {stage5_21[3]}
   );
   gpc1_1 gpc382 (
      {stage4_22[6]},
      {stage5_22[1]}
   );
   gpc1_1 gpc383 (
      {stage4_22[7]},
      {stage5_22[2]}
   );
   gpc1_1 gpc384 (
      {stage4_22[8]},
      {stage5_22[3]}
   );
   gpc1_1 gpc385 (
      {stage4_22[9]},
      {stage5_22[4]}
   );
   gpc1_1 gpc386 (
      {stage4_23[5]},
      {stage5_23[2]}
   );
   gpc1_1 gpc387 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc388 (
      {stage4_24[1]},
      {stage5_24[2]}
   );
   gpc1_1 gpc389 (
      {stage4_24[2]},
      {stage5_24[3]}
   );
   gpc1_1 gpc390 (
      {stage4_24[3]},
      {stage5_24[4]}
   );
   gpc1_1 gpc391 (
      {stage4_24[4]},
      {stage5_24[5]}
   );
   gpc1_1 gpc392 (
      {stage4_26[1]},
      {stage5_26[1]}
   );
   gpc1_1 gpc393 (
      {stage4_26[2]},
      {stage5_26[2]}
   );
   gpc1_1 gpc394 (
      {stage4_27[0]},
      {stage5_27[1]}
   );
   gpc1_1 gpc395 (
      {stage4_27[1]},
      {stage5_27[2]}
   );
   gpc1_1 gpc396 (
      {stage4_28[0]},
      {stage5_28[0]}
   );
   gpc1343_5 gpc397 (
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[0]}
   );
   gpc615_5 gpc398 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[0],stage6_22[0]}
   );
   gpc1_1 gpc399 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc400 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc401 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc402 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc403 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc404 (
      {stage5_5[0]},
      {stage6_5[0]}
   );
   gpc1_1 gpc405 (
      {stage5_6[0]},
      {stage6_6[0]}
   );
   gpc1_1 gpc406 (
      {stage5_7[0]},
      {stage6_7[0]}
   );
   gpc1_1 gpc407 (
      {stage5_8[0]},
      {stage6_8[0]}
   );
   gpc1_1 gpc408 (
      {stage5_9[0]},
      {stage6_9[0]}
   );
   gpc1_1 gpc409 (
      {stage5_10[0]},
      {stage6_10[0]}
   );
   gpc1_1 gpc410 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc411 (
      {stage5_12[0]},
      {stage6_12[0]}
   );
   gpc1_1 gpc412 (
      {stage5_13[0]},
      {stage6_13[0]}
   );
   gpc1_1 gpc413 (
      {stage5_14[0]},
      {stage6_14[0]}
   );
   gpc1_1 gpc414 (
      {stage5_15[0]},
      {stage6_15[0]}
   );
   gpc1_1 gpc415 (
      {stage5_16[0]},
      {stage6_16[0]}
   );
   gpc1_1 gpc416 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc417 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc418 (
      {stage5_21[2]},
      {stage6_21[3]}
   );
   gpc1_1 gpc419 (
      {stage5_21[3]},
      {stage6_21[4]}
   );
   gpc1_1 gpc420 (
      {stage5_23[1]},
      {stage6_23[1]}
   );
   gpc1_1 gpc421 (
      {stage5_23[2]},
      {stage6_23[2]}
   );
   gpc1_1 gpc422 (
      {stage5_23[3]},
      {stage6_23[3]}
   );
   gpc1_1 gpc423 (
      {stage5_25[0]},
      {stage6_25[1]}
   );
   gpc1_1 gpc424 (
      {stage5_26[0]},
      {stage6_26[1]}
   );
   gpc1_1 gpc425 (
      {stage5_26[1]},
      {stage6_26[2]}
   );
   gpc1_1 gpc426 (
      {stage5_26[2]},
      {stage6_26[3]}
   );
   gpc1_1 gpc427 (
      {stage5_27[0]},
      {stage6_27[0]}
   );
   gpc1_1 gpc428 (
      {stage5_27[1]},
      {stage6_27[1]}
   );
   gpc1_1 gpc429 (
      {stage5_27[2]},
      {stage6_27[2]}
   );
   gpc1_1 gpc430 (
      {stage5_28[0]},
      {stage6_28[0]}
   );
   gpc1415_5 gpc431 (
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4]},
      {stage6_22[0]},
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[0],stage7_22[0],stage7_21[0]}
   );
   gpc1_1 gpc432 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc433 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc434 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc435 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc436 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc437 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc438 (
      {stage6_6[0]},
      {stage7_6[0]}
   );
   gpc1_1 gpc439 (
      {stage6_7[0]},
      {stage7_7[0]}
   );
   gpc1_1 gpc440 (
      {stage6_8[0]},
      {stage7_8[0]}
   );
   gpc1_1 gpc441 (
      {stage6_9[0]},
      {stage7_9[0]}
   );
   gpc1_1 gpc442 (
      {stage6_10[0]},
      {stage7_10[0]}
   );
   gpc1_1 gpc443 (
      {stage6_11[0]},
      {stage7_11[0]}
   );
   gpc1_1 gpc444 (
      {stage6_12[0]},
      {stage7_12[0]}
   );
   gpc1_1 gpc445 (
      {stage6_13[0]},
      {stage7_13[0]}
   );
   gpc1_1 gpc446 (
      {stage6_14[0]},
      {stage7_14[0]}
   );
   gpc1_1 gpc447 (
      {stage6_15[0]},
      {stage7_15[0]}
   );
   gpc1_1 gpc448 (
      {stage6_16[0]},
      {stage7_16[0]}
   );
   gpc1_1 gpc449 (
      {stage6_17[0]},
      {stage7_17[0]}
   );
   gpc1_1 gpc450 (
      {stage6_18[0]},
      {stage7_18[0]}
   );
   gpc1_1 gpc451 (
      {stage6_19[0]},
      {stage7_19[0]}
   );
   gpc1_1 gpc452 (
      {stage6_20[0]},
      {stage7_20[0]}
   );
   gpc1_1 gpc453 (
      {stage6_25[0]},
      {stage7_25[1]}
   );
   gpc1_1 gpc454 (
      {stage6_25[1]},
      {stage7_25[2]}
   );
   gpc1_1 gpc455 (
      {stage6_26[0]},
      {stage7_26[0]}
   );
   gpc1_1 gpc456 (
      {stage6_26[1]},
      {stage7_26[1]}
   );
   gpc1_1 gpc457 (
      {stage6_26[2]},
      {stage7_26[2]}
   );
   gpc1_1 gpc458 (
      {stage6_26[3]},
      {stage7_26[3]}
   );
   gpc1_1 gpc459 (
      {stage6_27[0]},
      {stage7_27[0]}
   );
   gpc1_1 gpc460 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc461 (
      {stage6_27[2]},
      {stage7_27[2]}
   );
   gpc1_1 gpc462 (
      {stage6_28[0]},
      {stage7_28[0]}
   );
   gpc1343_5 gpc463 (
      {stage7_25[0], stage7_25[1], stage7_25[2]},
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3]},
      {stage7_27[0], stage7_27[1], stage7_27[2]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[0],stage8_27[0],stage8_26[0],stage8_25[0]}
   );
   gpc1_1 gpc464 (
      {stage7_0[0]},
      {stage8_0[0]}
   );
   gpc1_1 gpc465 (
      {stage7_1[0]},
      {stage8_1[0]}
   );
   gpc1_1 gpc466 (
      {stage7_2[0]},
      {stage8_2[0]}
   );
   gpc1_1 gpc467 (
      {stage7_3[0]},
      {stage8_3[0]}
   );
   gpc1_1 gpc468 (
      {stage7_4[0]},
      {stage8_4[0]}
   );
   gpc1_1 gpc469 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc470 (
      {stage7_6[0]},
      {stage8_6[0]}
   );
   gpc1_1 gpc471 (
      {stage7_7[0]},
      {stage8_7[0]}
   );
   gpc1_1 gpc472 (
      {stage7_8[0]},
      {stage8_8[0]}
   );
   gpc1_1 gpc473 (
      {stage7_9[0]},
      {stage8_9[0]}
   );
   gpc1_1 gpc474 (
      {stage7_10[0]},
      {stage8_10[0]}
   );
   gpc1_1 gpc475 (
      {stage7_11[0]},
      {stage8_11[0]}
   );
   gpc1_1 gpc476 (
      {stage7_12[0]},
      {stage8_12[0]}
   );
   gpc1_1 gpc477 (
      {stage7_13[0]},
      {stage8_13[0]}
   );
   gpc1_1 gpc478 (
      {stage7_14[0]},
      {stage8_14[0]}
   );
   gpc1_1 gpc479 (
      {stage7_15[0]},
      {stage8_15[0]}
   );
   gpc1_1 gpc480 (
      {stage7_16[0]},
      {stage8_16[0]}
   );
   gpc1_1 gpc481 (
      {stage7_17[0]},
      {stage8_17[0]}
   );
   gpc1_1 gpc482 (
      {stage7_18[0]},
      {stage8_18[0]}
   );
   gpc1_1 gpc483 (
      {stage7_19[0]},
      {stage8_19[0]}
   );
   gpc1_1 gpc484 (
      {stage7_20[0]},
      {stage8_20[0]}
   );
   gpc1_1 gpc485 (
      {stage7_21[0]},
      {stage8_21[0]}
   );
   gpc1_1 gpc486 (
      {stage7_22[0]},
      {stage8_22[0]}
   );
   gpc1_1 gpc487 (
      {stage7_23[0]},
      {stage8_23[0]}
   );
   gpc1_1 gpc488 (
      {stage7_24[0]},
      {stage8_24[0]}
   );
   gpc1_1 gpc489 (
      {stage8_0[0]},
      {stage9_0[0]}
   );
   gpc1_1 gpc490 (
      {stage8_1[0]},
      {stage9_1[0]}
   );
   gpc1_1 gpc491 (
      {stage8_2[0]},
      {stage9_2[0]}
   );
   gpc1_1 gpc492 (
      {stage8_3[0]},
      {stage9_3[0]}
   );
   gpc1_1 gpc493 (
      {stage8_4[0]},
      {stage9_4[0]}
   );
   gpc1_1 gpc494 (
      {stage8_5[0]},
      {stage9_5[0]}
   );
   gpc1_1 gpc495 (
      {stage8_6[0]},
      {stage9_6[0]}
   );
   gpc1_1 gpc496 (
      {stage8_7[0]},
      {stage9_7[0]}
   );
   gpc1_1 gpc497 (
      {stage8_8[0]},
      {stage9_8[0]}
   );
   gpc1_1 gpc498 (
      {stage8_9[0]},
      {stage9_9[0]}
   );
   gpc1_1 gpc499 (
      {stage8_10[0]},
      {stage9_10[0]}
   );
   gpc1_1 gpc500 (
      {stage8_11[0]},
      {stage9_11[0]}
   );
   gpc1_1 gpc501 (
      {stage8_12[0]},
      {stage9_12[0]}
   );
   gpc1_1 gpc502 (
      {stage8_13[0]},
      {stage9_13[0]}
   );
   gpc1_1 gpc503 (
      {stage8_14[0]},
      {stage9_14[0]}
   );
   gpc1_1 gpc504 (
      {stage8_15[0]},
      {stage9_15[0]}
   );
   gpc1_1 gpc505 (
      {stage8_16[0]},
      {stage9_16[0]}
   );
   gpc1_1 gpc506 (
      {stage8_17[0]},
      {stage9_17[0]}
   );
   gpc1_1 gpc507 (
      {stage8_18[0]},
      {stage9_18[0]}
   );
   gpc1_1 gpc508 (
      {stage8_19[0]},
      {stage9_19[0]}
   );
   gpc1_1 gpc509 (
      {stage8_20[0]},
      {stage9_20[0]}
   );
   gpc1_1 gpc510 (
      {stage8_21[0]},
      {stage9_21[0]}
   );
   gpc1_1 gpc511 (
      {stage8_22[0]},
      {stage9_22[0]}
   );
   gpc1_1 gpc512 (
      {stage8_23[0]},
      {stage9_23[0]}
   );
   gpc1_1 gpc513 (
      {stage8_24[0]},
      {stage9_24[0]}
   );
   gpc1_1 gpc514 (
      {stage8_25[0]},
      {stage9_25[0]}
   );
   gpc1_1 gpc515 (
      {stage8_26[0]},
      {stage9_26[0]}
   );
   gpc1_1 gpc516 (
      {stage8_27[0]},
      {stage9_27[0]}
   );
   gpc1_1 gpc517 (
      {stage8_28[0]},
      {stage9_28[0]}
   );
   gpc1_1 gpc518 (
      {stage8_29[0]},
      {stage9_29[0]}
   );
endmodule
