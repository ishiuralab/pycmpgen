module compressor2_1_162_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, input in_data128, input in_data129, input in_data130, input in_data131, input in_data132, input in_data133, input in_data134, input in_data135, input in_data136, input in_data137, input in_data138, input in_data139, input in_data140, input in_data141, input in_data142, input in_data143, input in_data144, input in_data145, input in_data146, input in_data147, input in_data148, input in_data149, input in_data150, input in_data151, input in_data152, input in_data153, input in_data154, input in_data155, input in_data156, input in_data157, input in_data158, input in_data159, input in_data160, input in_data161, output [23:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    reg [15:0] src128;
    reg [15:0] src129;
    reg [15:0] src130;
    reg [15:0] src131;
    reg [15:0] src132;
    reg [15:0] src133;
    reg [15:0] src134;
    reg [15:0] src135;
    reg [15:0] src136;
    reg [15:0] src137;
    reg [15:0] src138;
    reg [15:0] src139;
    reg [15:0] src140;
    reg [15:0] src141;
    reg [15:0] src142;
    reg [15:0] src143;
    reg [15:0] src144;
    reg [15:0] src145;
    reg [15:0] src146;
    reg [15:0] src147;
    reg [15:0] src148;
    reg [15:0] src149;
    reg [15:0] src150;
    reg [15:0] src151;
    reg [15:0] src152;
    reg [15:0] src153;
    reg [15:0] src154;
    reg [15:0] src155;
    reg [15:0] src156;
    reg [15:0] src157;
    reg [15:0] src158;
    reg [15:0] src159;
    reg [15:0] src160;
    reg [15:0] src161;
    compressor2_1_162_16 compressor2_1_162_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .src128(src128), .src129(src129), .src130(src130), .src131(src131), .src132(src132), .src133(src133), .src134(src134), .src135(src135), .src136(src136), .src137(src137), .src138(src138), .src139(src139), .src140(src140), .src141(src141), .src142(src142), .src143(src143), .src144(src144), .src145(src145), .src146(src146), .src147(src147), .src148(src148), .src149(src149), .src150(src150), .src151(src151), .src152(src152), .src153(src153), .src154(src154), .src155(src155), .src156(src156), .src157(src157), .src158(src158), .src159(src159), .src160(src160), .src161(src161), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
        src128 <= 0;
        src129 <= 0;
        src130 <= 0;
        src131 <= 0;
        src132 <= 0;
        src133 <= 0;
        src134 <= 0;
        src135 <= 0;
        src136 <= 0;
        src137 <= 0;
        src138 <= 0;
        src139 <= 0;
        src140 <= 0;
        src141 <= 0;
        src142 <= 0;
        src143 <= 0;
        src144 <= 0;
        src145 <= 0;
        src146 <= 0;
        src147 <= 0;
        src148 <= 0;
        src149 <= 0;
        src150 <= 0;
        src151 <= 0;
        src152 <= 0;
        src153 <= 0;
        src154 <= 0;
        src155 <= 0;
        src156 <= 0;
        src157 <= 0;
        src158 <= 0;
        src159 <= 0;
        src160 <= 0;
        src161 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
        src32 <= {src32[14:0], in_data32};
        src33 <= {src33[14:0], in_data33};
        src34 <= {src34[14:0], in_data34};
        src35 <= {src35[14:0], in_data35};
        src36 <= {src36[14:0], in_data36};
        src37 <= {src37[14:0], in_data37};
        src38 <= {src38[14:0], in_data38};
        src39 <= {src39[14:0], in_data39};
        src40 <= {src40[14:0], in_data40};
        src41 <= {src41[14:0], in_data41};
        src42 <= {src42[14:0], in_data42};
        src43 <= {src43[14:0], in_data43};
        src44 <= {src44[14:0], in_data44};
        src45 <= {src45[14:0], in_data45};
        src46 <= {src46[14:0], in_data46};
        src47 <= {src47[14:0], in_data47};
        src48 <= {src48[14:0], in_data48};
        src49 <= {src49[14:0], in_data49};
        src50 <= {src50[14:0], in_data50};
        src51 <= {src51[14:0], in_data51};
        src52 <= {src52[14:0], in_data52};
        src53 <= {src53[14:0], in_data53};
        src54 <= {src54[14:0], in_data54};
        src55 <= {src55[14:0], in_data55};
        src56 <= {src56[14:0], in_data56};
        src57 <= {src57[14:0], in_data57};
        src58 <= {src58[14:0], in_data58};
        src59 <= {src59[14:0], in_data59};
        src60 <= {src60[14:0], in_data60};
        src61 <= {src61[14:0], in_data61};
        src62 <= {src62[14:0], in_data62};
        src63 <= {src63[14:0], in_data63};
        src64 <= {src64[14:0], in_data64};
        src65 <= {src65[14:0], in_data65};
        src66 <= {src66[14:0], in_data66};
        src67 <= {src67[14:0], in_data67};
        src68 <= {src68[14:0], in_data68};
        src69 <= {src69[14:0], in_data69};
        src70 <= {src70[14:0], in_data70};
        src71 <= {src71[14:0], in_data71};
        src72 <= {src72[14:0], in_data72};
        src73 <= {src73[14:0], in_data73};
        src74 <= {src74[14:0], in_data74};
        src75 <= {src75[14:0], in_data75};
        src76 <= {src76[14:0], in_data76};
        src77 <= {src77[14:0], in_data77};
        src78 <= {src78[14:0], in_data78};
        src79 <= {src79[14:0], in_data79};
        src80 <= {src80[14:0], in_data80};
        src81 <= {src81[14:0], in_data81};
        src82 <= {src82[14:0], in_data82};
        src83 <= {src83[14:0], in_data83};
        src84 <= {src84[14:0], in_data84};
        src85 <= {src85[14:0], in_data85};
        src86 <= {src86[14:0], in_data86};
        src87 <= {src87[14:0], in_data87};
        src88 <= {src88[14:0], in_data88};
        src89 <= {src89[14:0], in_data89};
        src90 <= {src90[14:0], in_data90};
        src91 <= {src91[14:0], in_data91};
        src92 <= {src92[14:0], in_data92};
        src93 <= {src93[14:0], in_data93};
        src94 <= {src94[14:0], in_data94};
        src95 <= {src95[14:0], in_data95};
        src96 <= {src96[14:0], in_data96};
        src97 <= {src97[14:0], in_data97};
        src98 <= {src98[14:0], in_data98};
        src99 <= {src99[14:0], in_data99};
        src100 <= {src100[14:0], in_data100};
        src101 <= {src101[14:0], in_data101};
        src102 <= {src102[14:0], in_data102};
        src103 <= {src103[14:0], in_data103};
        src104 <= {src104[14:0], in_data104};
        src105 <= {src105[14:0], in_data105};
        src106 <= {src106[14:0], in_data106};
        src107 <= {src107[14:0], in_data107};
        src108 <= {src108[14:0], in_data108};
        src109 <= {src109[14:0], in_data109};
        src110 <= {src110[14:0], in_data110};
        src111 <= {src111[14:0], in_data111};
        src112 <= {src112[14:0], in_data112};
        src113 <= {src113[14:0], in_data113};
        src114 <= {src114[14:0], in_data114};
        src115 <= {src115[14:0], in_data115};
        src116 <= {src116[14:0], in_data116};
        src117 <= {src117[14:0], in_data117};
        src118 <= {src118[14:0], in_data118};
        src119 <= {src119[14:0], in_data119};
        src120 <= {src120[14:0], in_data120};
        src121 <= {src121[14:0], in_data121};
        src122 <= {src122[14:0], in_data122};
        src123 <= {src123[14:0], in_data123};
        src124 <= {src124[14:0], in_data124};
        src125 <= {src125[14:0], in_data125};
        src126 <= {src126[14:0], in_data126};
        src127 <= {src127[14:0], in_data127};
        src128 <= {src128[14:0], in_data128};
        src129 <= {src129[14:0], in_data129};
        src130 <= {src130[14:0], in_data130};
        src131 <= {src131[14:0], in_data131};
        src132 <= {src132[14:0], in_data132};
        src133 <= {src133[14:0], in_data133};
        src134 <= {src134[14:0], in_data134};
        src135 <= {src135[14:0], in_data135};
        src136 <= {src136[14:0], in_data136};
        src137 <= {src137[14:0], in_data137};
        src138 <= {src138[14:0], in_data138};
        src139 <= {src139[14:0], in_data139};
        src140 <= {src140[14:0], in_data140};
        src141 <= {src141[14:0], in_data141};
        src142 <= {src142[14:0], in_data142};
        src143 <= {src143[14:0], in_data143};
        src144 <= {src144[14:0], in_data144};
        src145 <= {src145[14:0], in_data145};
        src146 <= {src146[14:0], in_data146};
        src147 <= {src147[14:0], in_data147};
        src148 <= {src148[14:0], in_data148};
        src149 <= {src149[14:0], in_data149};
        src150 <= {src150[14:0], in_data150};
        src151 <= {src151[14:0], in_data151};
        src152 <= {src152[14:0], in_data152};
        src153 <= {src153[14:0], in_data153};
        src154 <= {src154[14:0], in_data154};
        src155 <= {src155[14:0], in_data155};
        src156 <= {src156[14:0], in_data156};
        src157 <= {src157[14:0], in_data157};
        src158 <= {src158[14:0], in_data158};
        src159 <= {src159[14:0], in_data159};
        src160 <= {src160[14:0], in_data160};
        src161 <= {src161[14:0], in_data161};
    end
endmodule

module compressor2_1_162_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    input [15:0]src64,
    input [15:0]src65,
    input [15:0]src66,
    input [15:0]src67,
    input [15:0]src68,
    input [15:0]src69,
    input [15:0]src70,
    input [15:0]src71,
    input [15:0]src72,
    input [15:0]src73,
    input [15:0]src74,
    input [15:0]src75,
    input [15:0]src76,
    input [15:0]src77,
    input [15:0]src78,
    input [15:0]src79,
    input [15:0]src80,
    input [15:0]src81,
    input [15:0]src82,
    input [15:0]src83,
    input [15:0]src84,
    input [15:0]src85,
    input [15:0]src86,
    input [15:0]src87,
    input [15:0]src88,
    input [15:0]src89,
    input [15:0]src90,
    input [15:0]src91,
    input [15:0]src92,
    input [15:0]src93,
    input [15:0]src94,
    input [15:0]src95,
    input [15:0]src96,
    input [15:0]src97,
    input [15:0]src98,
    input [15:0]src99,
    input [15:0]src100,
    input [15:0]src101,
    input [15:0]src102,
    input [15:0]src103,
    input [15:0]src104,
    input [15:0]src105,
    input [15:0]src106,
    input [15:0]src107,
    input [15:0]src108,
    input [15:0]src109,
    input [15:0]src110,
    input [15:0]src111,
    input [15:0]src112,
    input [15:0]src113,
    input [15:0]src114,
    input [15:0]src115,
    input [15:0]src116,
    input [15:0]src117,
    input [15:0]src118,
    input [15:0]src119,
    input [15:0]src120,
    input [15:0]src121,
    input [15:0]src122,
    input [15:0]src123,
    input [15:0]src124,
    input [15:0]src125,
    input [15:0]src126,
    input [15:0]src127,
    input [15:0]src128,
    input [15:0]src129,
    input [15:0]src130,
    input [15:0]src131,
    input [15:0]src132,
    input [15:0]src133,
    input [15:0]src134,
    input [15:0]src135,
    input [15:0]src136,
    input [15:0]src137,
    input [15:0]src138,
    input [15:0]src139,
    input [15:0]src140,
    input [15:0]src141,
    input [15:0]src142,
    input [15:0]src143,
    input [15:0]src144,
    input [15:0]src145,
    input [15:0]src146,
    input [15:0]src147,
    input [15:0]src148,
    input [15:0]src149,
    input [15:0]src150,
    input [15:0]src151,
    input [15:0]src152,
    input [15:0]src153,
    input [15:0]src154,
    input [15:0]src155,
    input [15:0]src156,
    input [15:0]src157,
    input [15:0]src158,
    input [15:0]src159,
    input [15:0]src160,
    input [15:0]src161,
    output [23:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [23:0] out;
    compressor compressor_inst(
        .src0({src161[0], src160[0], src159[0], src158[0], src157[0], src156[0], src155[0], src154[0], src153[0], src152[0], src151[0], src150[0], src149[0], src148[0], src147[0], src146[0], src145[0], src144[0], src143[0], src142[0], src141[0], src140[0], src139[0], src138[0], src137[0], src136[0], src135[0], src134[0], src133[0], src132[0], src131[0], src130[0], src129[0], src128[0], src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src161[1], src160[1], src159[1], src158[1], src157[1], src156[1], src155[1], src154[1], src153[1], src152[1], src151[1], src150[1], src149[1], src148[1], src147[1], src146[1], src145[1], src144[1], src143[1], src142[1], src141[1], src140[1], src139[1], src138[1], src137[1], src136[1], src135[1], src134[1], src133[1], src132[1], src131[1], src130[1], src129[1], src128[1], src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src161[2], src160[2], src159[2], src158[2], src157[2], src156[2], src155[2], src154[2], src153[2], src152[2], src151[2], src150[2], src149[2], src148[2], src147[2], src146[2], src145[2], src144[2], src143[2], src142[2], src141[2], src140[2], src139[2], src138[2], src137[2], src136[2], src135[2], src134[2], src133[2], src132[2], src131[2], src130[2], src129[2], src128[2], src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src161[3], src160[3], src159[3], src158[3], src157[3], src156[3], src155[3], src154[3], src153[3], src152[3], src151[3], src150[3], src149[3], src148[3], src147[3], src146[3], src145[3], src144[3], src143[3], src142[3], src141[3], src140[3], src139[3], src138[3], src137[3], src136[3], src135[3], src134[3], src133[3], src132[3], src131[3], src130[3], src129[3], src128[3], src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src161[4], src160[4], src159[4], src158[4], src157[4], src156[4], src155[4], src154[4], src153[4], src152[4], src151[4], src150[4], src149[4], src148[4], src147[4], src146[4], src145[4], src144[4], src143[4], src142[4], src141[4], src140[4], src139[4], src138[4], src137[4], src136[4], src135[4], src134[4], src133[4], src132[4], src131[4], src130[4], src129[4], src128[4], src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src161[5], src160[5], src159[5], src158[5], src157[5], src156[5], src155[5], src154[5], src153[5], src152[5], src151[5], src150[5], src149[5], src148[5], src147[5], src146[5], src145[5], src144[5], src143[5], src142[5], src141[5], src140[5], src139[5], src138[5], src137[5], src136[5], src135[5], src134[5], src133[5], src132[5], src131[5], src130[5], src129[5], src128[5], src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src161[6], src160[6], src159[6], src158[6], src157[6], src156[6], src155[6], src154[6], src153[6], src152[6], src151[6], src150[6], src149[6], src148[6], src147[6], src146[6], src145[6], src144[6], src143[6], src142[6], src141[6], src140[6], src139[6], src138[6], src137[6], src136[6], src135[6], src134[6], src133[6], src132[6], src131[6], src130[6], src129[6], src128[6], src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src161[7], src160[7], src159[7], src158[7], src157[7], src156[7], src155[7], src154[7], src153[7], src152[7], src151[7], src150[7], src149[7], src148[7], src147[7], src146[7], src145[7], src144[7], src143[7], src142[7], src141[7], src140[7], src139[7], src138[7], src137[7], src136[7], src135[7], src134[7], src133[7], src132[7], src131[7], src130[7], src129[7], src128[7], src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src161[8], src160[8], src159[8], src158[8], src157[8], src156[8], src155[8], src154[8], src153[8], src152[8], src151[8], src150[8], src149[8], src148[8], src147[8], src146[8], src145[8], src144[8], src143[8], src142[8], src141[8], src140[8], src139[8], src138[8], src137[8], src136[8], src135[8], src134[8], src133[8], src132[8], src131[8], src130[8], src129[8], src128[8], src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src161[9], src160[9], src159[9], src158[9], src157[9], src156[9], src155[9], src154[9], src153[9], src152[9], src151[9], src150[9], src149[9], src148[9], src147[9], src146[9], src145[9], src144[9], src143[9], src142[9], src141[9], src140[9], src139[9], src138[9], src137[9], src136[9], src135[9], src134[9], src133[9], src132[9], src131[9], src130[9], src129[9], src128[9], src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src161[10], src160[10], src159[10], src158[10], src157[10], src156[10], src155[10], src154[10], src153[10], src152[10], src151[10], src150[10], src149[10], src148[10], src147[10], src146[10], src145[10], src144[10], src143[10], src142[10], src141[10], src140[10], src139[10], src138[10], src137[10], src136[10], src135[10], src134[10], src133[10], src132[10], src131[10], src130[10], src129[10], src128[10], src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src161[11], src160[11], src159[11], src158[11], src157[11], src156[11], src155[11], src154[11], src153[11], src152[11], src151[11], src150[11], src149[11], src148[11], src147[11], src146[11], src145[11], src144[11], src143[11], src142[11], src141[11], src140[11], src139[11], src138[11], src137[11], src136[11], src135[11], src134[11], src133[11], src132[11], src131[11], src130[11], src129[11], src128[11], src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src161[12], src160[12], src159[12], src158[12], src157[12], src156[12], src155[12], src154[12], src153[12], src152[12], src151[12], src150[12], src149[12], src148[12], src147[12], src146[12], src145[12], src144[12], src143[12], src142[12], src141[12], src140[12], src139[12], src138[12], src137[12], src136[12], src135[12], src134[12], src133[12], src132[12], src131[12], src130[12], src129[12], src128[12], src127[12], src126[12], src125[12], src124[12], src123[12], src122[12], src121[12], src120[12], src119[12], src118[12], src117[12], src116[12], src115[12], src114[12], src113[12], src112[12], src111[12], src110[12], src109[12], src108[12], src107[12], src106[12], src105[12], src104[12], src103[12], src102[12], src101[12], src100[12], src99[12], src98[12], src97[12], src96[12], src95[12], src94[12], src93[12], src92[12], src91[12], src90[12], src89[12], src88[12], src87[12], src86[12], src85[12], src84[12], src83[12], src82[12], src81[12], src80[12], src79[12], src78[12], src77[12], src76[12], src75[12], src74[12], src73[12], src72[12], src71[12], src70[12], src69[12], src68[12], src67[12], src66[12], src65[12], src64[12], src63[12], src62[12], src61[12], src60[12], src59[12], src58[12], src57[12], src56[12], src55[12], src54[12], src53[12], src52[12], src51[12], src50[12], src49[12], src48[12], src47[12], src46[12], src45[12], src44[12], src43[12], src42[12], src41[12], src40[12], src39[12], src38[12], src37[12], src36[12], src35[12], src34[12], src33[12], src32[12], src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src161[13], src160[13], src159[13], src158[13], src157[13], src156[13], src155[13], src154[13], src153[13], src152[13], src151[13], src150[13], src149[13], src148[13], src147[13], src146[13], src145[13], src144[13], src143[13], src142[13], src141[13], src140[13], src139[13], src138[13], src137[13], src136[13], src135[13], src134[13], src133[13], src132[13], src131[13], src130[13], src129[13], src128[13], src127[13], src126[13], src125[13], src124[13], src123[13], src122[13], src121[13], src120[13], src119[13], src118[13], src117[13], src116[13], src115[13], src114[13], src113[13], src112[13], src111[13], src110[13], src109[13], src108[13], src107[13], src106[13], src105[13], src104[13], src103[13], src102[13], src101[13], src100[13], src99[13], src98[13], src97[13], src96[13], src95[13], src94[13], src93[13], src92[13], src91[13], src90[13], src89[13], src88[13], src87[13], src86[13], src85[13], src84[13], src83[13], src82[13], src81[13], src80[13], src79[13], src78[13], src77[13], src76[13], src75[13], src74[13], src73[13], src72[13], src71[13], src70[13], src69[13], src68[13], src67[13], src66[13], src65[13], src64[13], src63[13], src62[13], src61[13], src60[13], src59[13], src58[13], src57[13], src56[13], src55[13], src54[13], src53[13], src52[13], src51[13], src50[13], src49[13], src48[13], src47[13], src46[13], src45[13], src44[13], src43[13], src42[13], src41[13], src40[13], src39[13], src38[13], src37[13], src36[13], src35[13], src34[13], src33[13], src32[13], src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src161[14], src160[14], src159[14], src158[14], src157[14], src156[14], src155[14], src154[14], src153[14], src152[14], src151[14], src150[14], src149[14], src148[14], src147[14], src146[14], src145[14], src144[14], src143[14], src142[14], src141[14], src140[14], src139[14], src138[14], src137[14], src136[14], src135[14], src134[14], src133[14], src132[14], src131[14], src130[14], src129[14], src128[14], src127[14], src126[14], src125[14], src124[14], src123[14], src122[14], src121[14], src120[14], src119[14], src118[14], src117[14], src116[14], src115[14], src114[14], src113[14], src112[14], src111[14], src110[14], src109[14], src108[14], src107[14], src106[14], src105[14], src104[14], src103[14], src102[14], src101[14], src100[14], src99[14], src98[14], src97[14], src96[14], src95[14], src94[14], src93[14], src92[14], src91[14], src90[14], src89[14], src88[14], src87[14], src86[14], src85[14], src84[14], src83[14], src82[14], src81[14], src80[14], src79[14], src78[14], src77[14], src76[14], src75[14], src74[14], src73[14], src72[14], src71[14], src70[14], src69[14], src68[14], src67[14], src66[14], src65[14], src64[14], src63[14], src62[14], src61[14], src60[14], src59[14], src58[14], src57[14], src56[14], src55[14], src54[14], src53[14], src52[14], src51[14], src50[14], src49[14], src48[14], src47[14], src46[14], src45[14], src44[14], src43[14], src42[14], src41[14], src40[14], src39[14], src38[14], src37[14], src36[14], src35[14], src34[14], src33[14], src32[14], src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src161[15], src160[15], src159[15], src158[15], src157[15], src156[15], src155[15], src154[15], src153[15], src152[15], src151[15], src150[15], src149[15], src148[15], src147[15], src146[15], src145[15], src144[15], src143[15], src142[15], src141[15], src140[15], src139[15], src138[15], src137[15], src136[15], src135[15], src134[15], src133[15], src132[15], src131[15], src130[15], src129[15], src128[15], src127[15], src126[15], src125[15], src124[15], src123[15], src122[15], src121[15], src120[15], src119[15], src118[15], src117[15], src116[15], src115[15], src114[15], src113[15], src112[15], src111[15], src110[15], src109[15], src108[15], src107[15], src106[15], src105[15], src104[15], src103[15], src102[15], src101[15], src100[15], src99[15], src98[15], src97[15], src96[15], src95[15], src94[15], src93[15], src92[15], src91[15], src90[15], src89[15], src88[15], src87[15], src86[15], src85[15], src84[15], src83[15], src82[15], src81[15], src80[15], src79[15], src78[15], src77[15], src76[15], src75[15], src74[15], src73[15], src72[15], src71[15], src70[15], src69[15], src68[15], src67[15], src66[15], src65[15], src64[15], src63[15], src62[15], src61[15], src60[15], src59[15], src58[15], src57[15], src56[15], src55[15], src54[15], src53[15], src52[15], src51[15], src50[15], src49[15], src48[15], src47[15], src46[15], src45[15], src44[15], src43[15], src42[15], src41[15], src40[15], src39[15], src38[15], src37[15], src36[15], src35[15], src34[15], src33[15], src32[15], src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    rowadder2_1_23 rowadder2_1inst(
        .src0({comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[23:0];
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [32:0] stage1_0;
   wire [47:0] stage1_1;
   wire [63:0] stage1_2;
   wire [91:0] stage1_3;
   wire [74:0] stage1_4;
   wire [70:0] stage1_5;
   wire [59:0] stage1_6;
   wire [53:0] stage1_7;
   wire [89:0] stage1_8;
   wire [82:0] stage1_9;
   wire [60:0] stage1_10;
   wire [57:0] stage1_11;
   wire [72:0] stage1_12;
   wire [77:0] stage1_13;
   wire [77:0] stage1_14;
   wire [53:0] stage1_15;
   wire [48:0] stage1_16;
   wire [27:0] stage1_17;
   wire [10:0] stage2_0;
   wire [29:0] stage2_1;
   wire [15:0] stage2_2;
   wire [36:0] stage2_3;
   wire [29:0] stage2_4;
   wire [29:0] stage2_5;
   wire [29:0] stage2_6;
   wire [38:0] stage2_7;
   wire [29:0] stage2_8;
   wire [51:0] stage2_9;
   wire [25:0] stage2_10;
   wire [28:0] stage2_11;
   wire [33:0] stage2_12;
   wire [26:0] stage2_13;
   wire [29:0] stage2_14;
   wire [50:0] stage2_15;
   wire [17:0] stage2_16;
   wire [34:0] stage2_17;
   wire [8:0] stage2_18;
   wire [0:0] stage2_19;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [18:0] stage3_2;
   wire [13:0] stage3_3;
   wire [14:0] stage3_4;
   wire [11:0] stage3_5;
   wire [10:0] stage3_6;
   wire [13:0] stage3_7;
   wire [16:0] stage3_8;
   wire [19:0] stage3_9;
   wire [14:0] stage3_10;
   wire [12:0] stage3_11;
   wire [15:0] stage3_12;
   wire [15:0] stage3_13;
   wire [9:0] stage3_14;
   wire [17:0] stage3_15;
   wire [14:0] stage3_16;
   wire [10:0] stage3_17;
   wire [10:0] stage3_18;
   wire [7:0] stage3_19;
   wire [0:0] stage3_20;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [10:0] stage4_2;
   wire [5:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [6:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [6:0] stage4_9;
   wire [9:0] stage4_10;
   wire [11:0] stage4_11;
   wire [6:0] stage4_12;
   wire [5:0] stage4_13;
   wire [7:0] stage4_14;
   wire [3:0] stage4_15;
   wire [5:0] stage4_16;
   wire [10:0] stage4_17;
   wire [6:0] stage4_18;
   wire [8:0] stage4_19;
   wire [2:0] stage4_20;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [4:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [2:0] stage5_8;
   wire [4:0] stage5_9;
   wire [3:0] stage5_10;
   wire [3:0] stage5_11;
   wire [5:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [2:0] stage5_15;
   wire [1:0] stage5_16;
   wire [4:0] stage5_17;
   wire [2:0] stage5_18;
   wire [9:0] stage5_19;
   wire [1:0] stage5_20;
   wire [0:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[8]},
      {stage0_3[16]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[9]},
      {stage0_3[17]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[10]},
      {stage0_3[18]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[11]},
      {stage0_3[19]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[12]},
      {stage0_3[20]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[13]},
      {stage0_3[21]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27]},
      {stage1_5[0],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[1],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[2],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[3],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[4],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[5],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[6],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[7],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[8],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[9],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[10],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[11],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[12],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[13],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[14],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[15],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[16],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[17],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc606_5 gpc49 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[18],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc606_5 gpc50 (
      {stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[19],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc606_5 gpc51 (
      {stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[20],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc606_5 gpc52 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[21],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc606_5 gpc53 (
      {stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[22],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[6],stage1_5[23],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[7],stage1_5[24],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[8],stage1_5[25],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[9],stage1_5[26],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[10],stage1_5[27],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[11],stage1_5[28],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[12],stage1_5[29],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[13],stage1_5[30],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[14],stage1_5[31],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[15],stage1_5[32],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[16],stage1_5[33],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[17],stage1_5[34],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[18],stage1_5[35],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[19],stage1_5[36],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[20],stage1_5[37],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[21],stage1_5[38],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[22],stage1_5[39],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[23],stage1_5[40],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[24],stage1_5[41],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[25],stage1_5[42],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[20],stage1_6[26],stage1_5[43],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[21],stage1_7[21],stage1_6[27],stage1_5[44]}
   );
   gpc606_5 gpc76 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[22],stage1_7[22],stage1_6[28],stage1_5[45]}
   );
   gpc606_5 gpc77 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[23],stage1_7[23],stage1_6[29],stage1_5[46]}
   );
   gpc606_5 gpc78 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[24],stage1_7[24],stage1_6[30],stage1_5[47]}
   );
   gpc606_5 gpc79 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[25],stage1_7[25],stage1_6[31],stage1_5[48]}
   );
   gpc606_5 gpc80 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[26],stage1_7[26],stage1_6[32],stage1_5[49]}
   );
   gpc606_5 gpc81 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[27],stage1_7[27],stage1_6[33],stage1_5[50]}
   );
   gpc606_5 gpc82 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[28],stage1_7[28],stage1_6[34],stage1_5[51]}
   );
   gpc606_5 gpc83 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[29],stage1_7[29],stage1_6[35],stage1_5[52]}
   );
   gpc606_5 gpc84 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[30],stage1_7[30],stage1_6[36],stage1_5[53]}
   );
   gpc606_5 gpc85 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[31],stage1_7[31],stage1_6[37],stage1_5[54]}
   );
   gpc606_5 gpc86 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[32],stage1_7[32],stage1_6[38],stage1_5[55]}
   );
   gpc606_5 gpc87 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[33],stage1_7[33],stage1_6[39],stage1_5[56]}
   );
   gpc606_5 gpc88 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[34],stage1_7[34],stage1_6[40],stage1_5[57]}
   );
   gpc606_5 gpc89 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[35],stage1_7[35],stage1_6[41],stage1_5[58]}
   );
   gpc606_5 gpc90 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[36],stage1_7[36],stage1_6[42],stage1_5[59]}
   );
   gpc606_5 gpc91 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[37],stage1_7[37],stage1_6[43],stage1_5[60]}
   );
   gpc606_5 gpc92 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[38],stage1_7[38],stage1_6[44],stage1_5[61]}
   );
   gpc606_5 gpc93 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[39],stage1_7[39],stage1_6[45],stage1_5[62]}
   );
   gpc606_5 gpc94 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[40],stage1_7[40],stage1_6[46],stage1_5[63]}
   );
   gpc606_5 gpc95 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[41],stage1_7[41],stage1_6[47],stage1_5[64]}
   );
   gpc606_5 gpc96 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[42],stage1_7[42],stage1_6[48],stage1_5[65]}
   );
   gpc606_5 gpc97 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[43],stage1_7[43],stage1_6[49],stage1_5[66]}
   );
   gpc606_5 gpc98 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[44],stage1_7[44],stage1_6[50],stage1_5[67]}
   );
   gpc606_5 gpc99 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[45],stage1_7[45],stage1_6[51],stage1_5[68]}
   );
   gpc606_5 gpc100 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[46],stage1_7[46],stage1_6[52],stage1_5[69]}
   );
   gpc606_5 gpc101 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[47],stage1_7[47],stage1_6[53],stage1_5[70]}
   );
   gpc606_5 gpc102 (
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[48],stage1_7[48],stage1_6[54]}
   );
   gpc606_5 gpc103 (
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[49],stage1_7[49],stage1_6[55]}
   );
   gpc606_5 gpc104 (
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[50],stage1_7[50],stage1_6[56]}
   );
   gpc606_5 gpc105 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[51],stage1_7[51],stage1_6[57]}
   );
   gpc606_5 gpc106 (
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[52],stage1_7[52],stage1_6[58]}
   );
   gpc606_5 gpc107 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[53],stage1_7[53],stage1_6[59]}
   );
   gpc606_5 gpc108 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[6],stage1_9[33],stage1_8[54]}
   );
   gpc606_5 gpc109 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[7],stage1_9[34],stage1_8[55]}
   );
   gpc606_5 gpc110 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[8],stage1_9[35],stage1_8[56]}
   );
   gpc606_5 gpc111 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[9],stage1_9[36],stage1_8[57]}
   );
   gpc606_5 gpc112 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[10],stage1_9[37],stage1_8[58]}
   );
   gpc606_5 gpc113 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[11],stage1_9[38],stage1_8[59]}
   );
   gpc615_5 gpc114 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_9[0]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[12],stage1_9[39],stage1_8[60]}
   );
   gpc615_5 gpc115 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_9[1]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[13],stage1_9[40],stage1_8[61]}
   );
   gpc615_5 gpc116 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86]},
      {stage0_9[2]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[14],stage1_9[41],stage1_8[62]}
   );
   gpc615_5 gpc117 (
      {stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_9[3]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[15],stage1_9[42],stage1_8[63]}
   );
   gpc615_5 gpc118 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_9[4]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[16],stage1_9[43],stage1_8[64]}
   );
   gpc615_5 gpc119 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_9[5]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[17],stage1_9[44],stage1_8[65]}
   );
   gpc615_5 gpc120 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_9[6]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[18],stage1_9[45],stage1_8[66]}
   );
   gpc615_5 gpc121 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_9[7]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[19],stage1_9[46],stage1_8[67]}
   );
   gpc615_5 gpc122 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_9[8]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[20],stage1_9[47],stage1_8[68]}
   );
   gpc615_5 gpc123 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_9[9]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[21],stage1_9[48],stage1_8[69]}
   );
   gpc615_5 gpc124 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_9[10]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[22],stage1_9[49],stage1_8[70]}
   );
   gpc615_5 gpc125 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_9[11]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[23],stage1_9[50],stage1_8[71]}
   );
   gpc615_5 gpc126 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_9[12]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[24],stage1_9[51],stage1_8[72]}
   );
   gpc615_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_9[13]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[25],stage1_9[52],stage1_8[73]}
   );
   gpc615_5 gpc128 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_9[14]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[26],stage1_9[53],stage1_8[74]}
   );
   gpc606_5 gpc129 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[27],stage1_9[54]}
   );
   gpc606_5 gpc130 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[28],stage1_9[55]}
   );
   gpc606_5 gpc131 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[29],stage1_9[56]}
   );
   gpc606_5 gpc132 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[30],stage1_9[57]}
   );
   gpc606_5 gpc133 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[31],stage1_9[58]}
   );
   gpc606_5 gpc134 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[32],stage1_9[59]}
   );
   gpc606_5 gpc135 (
      {stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[33],stage1_9[60]}
   );
   gpc606_5 gpc136 (
      {stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[34],stage1_9[61]}
   );
   gpc606_5 gpc137 (
      {stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[35],stage1_9[62]}
   );
   gpc606_5 gpc138 (
      {stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[36],stage1_9[63]}
   );
   gpc606_5 gpc139 (
      {stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[37],stage1_9[64]}
   );
   gpc606_5 gpc140 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[38],stage1_9[65]}
   );
   gpc606_5 gpc141 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[39],stage1_9[66]}
   );
   gpc606_5 gpc142 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[40],stage1_9[67]}
   );
   gpc606_5 gpc143 (
      {stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[41],stage1_9[68]}
   );
   gpc606_5 gpc144 (
      {stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[42],stage1_9[69]}
   );
   gpc606_5 gpc145 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[43],stage1_9[70]}
   );
   gpc606_5 gpc146 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[44],stage1_9[71]}
   );
   gpc606_5 gpc147 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[45],stage1_9[72]}
   );
   gpc606_5 gpc148 (
      {stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[46],stage1_9[73]}
   );
   gpc606_5 gpc149 (
      {stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[47],stage1_9[74]}
   );
   gpc606_5 gpc150 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[42],stage1_11[42],stage1_10[48],stage1_9[75]}
   );
   gpc615_5 gpc151 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[126]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[43],stage1_11[43],stage1_10[49],stage1_9[76]}
   );
   gpc615_5 gpc152 (
      {stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_10[127]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[44],stage1_11[44],stage1_10[50],stage1_9[77]}
   );
   gpc615_5 gpc153 (
      {stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131], stage0_10[132]},
      {stage0_11[144]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[24],stage1_12[45],stage1_11[45],stage1_10[51]}
   );
   gpc615_5 gpc154 (
      {stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage0_11[145]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[25],stage1_12[46],stage1_11[46],stage1_10[52]}
   );
   gpc615_5 gpc155 (
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142]},
      {stage0_11[146]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[26],stage1_12[47],stage1_11[47],stage1_10[53]}
   );
   gpc615_5 gpc156 (
      {stage0_10[143], stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147]},
      {stage0_11[147]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[27],stage1_12[48],stage1_11[48],stage1_10[54]}
   );
   gpc615_5 gpc157 (
      {stage0_10[148], stage0_10[149], stage0_10[150], stage0_10[151], stage0_10[152]},
      {stage0_11[148]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[28],stage1_12[49],stage1_11[49],stage1_10[55]}
   );
   gpc615_5 gpc158 (
      {stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_11[149]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[29],stage1_12[50],stage1_11[50],stage1_10[56]}
   );
   gpc606_5 gpc159 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[30],stage1_12[51],stage1_11[51]}
   );
   gpc606_5 gpc160 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[7],stage1_13[31],stage1_12[52]}
   );
   gpc606_5 gpc161 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[8],stage1_13[32],stage1_12[53]}
   );
   gpc606_5 gpc162 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[9],stage1_13[33],stage1_12[54]}
   );
   gpc606_5 gpc163 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[10],stage1_13[34],stage1_12[55]}
   );
   gpc606_5 gpc164 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[11],stage1_13[35],stage1_12[56]}
   );
   gpc606_5 gpc165 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[12],stage1_13[36],stage1_12[57]}
   );
   gpc606_5 gpc166 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[13],stage1_13[37],stage1_12[58]}
   );
   gpc606_5 gpc167 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[14],stage1_13[38],stage1_12[59]}
   );
   gpc606_5 gpc168 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[15],stage1_13[39],stage1_12[60]}
   );
   gpc606_5 gpc169 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[10],stage1_14[16],stage1_13[40],stage1_12[61]}
   );
   gpc606_5 gpc170 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[11],stage1_14[17],stage1_13[41],stage1_12[62]}
   );
   gpc606_5 gpc171 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[12],stage1_14[18],stage1_13[42],stage1_12[63]}
   );
   gpc606_5 gpc172 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[13],stage1_14[19],stage1_13[43],stage1_12[64]}
   );
   gpc606_5 gpc173 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[14],stage1_14[20],stage1_13[44],stage1_12[65]}
   );
   gpc606_5 gpc174 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[15],stage1_14[21],stage1_13[45],stage1_12[66]}
   );
   gpc606_5 gpc175 (
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[16],stage1_14[22],stage1_13[46],stage1_12[67]}
   );
   gpc606_5 gpc176 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[17],stage1_14[23],stage1_13[47],stage1_12[68]}
   );
   gpc606_5 gpc177 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[18],stage1_14[24],stage1_13[48],stage1_12[69]}
   );
   gpc606_5 gpc178 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[19],stage1_14[25],stage1_13[49],stage1_12[70]}
   );
   gpc606_5 gpc179 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[20],stage1_14[26],stage1_13[50],stage1_12[71]}
   );
   gpc606_5 gpc180 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[21],stage1_14[27],stage1_13[51],stage1_12[72]}
   );
   gpc606_5 gpc181 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[21],stage1_15[22],stage1_14[28],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[22],stage1_15[23],stage1_14[29],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[23],stage1_15[24],stage1_14[30],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[24],stage1_15[25],stage1_14[31],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[25],stage1_15[26],stage1_14[32],stage1_13[56]}
   );
   gpc606_5 gpc186 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[26],stage1_15[27],stage1_14[33],stage1_13[57]}
   );
   gpc606_5 gpc187 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[27],stage1_15[28],stage1_14[34],stage1_13[58]}
   );
   gpc606_5 gpc188 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[28],stage1_15[29],stage1_14[35],stage1_13[59]}
   );
   gpc606_5 gpc189 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[29],stage1_15[30],stage1_14[36],stage1_13[60]}
   );
   gpc606_5 gpc190 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[30],stage1_15[31],stage1_14[37],stage1_13[61]}
   );
   gpc606_5 gpc191 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[31],stage1_15[32],stage1_14[38],stage1_13[62]}
   );
   gpc606_5 gpc192 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[32],stage1_15[33],stage1_14[39],stage1_13[63]}
   );
   gpc606_5 gpc193 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[33],stage1_15[34],stage1_14[40],stage1_13[64]}
   );
   gpc606_5 gpc194 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[34],stage1_15[35],stage1_14[41],stage1_13[65]}
   );
   gpc606_5 gpc195 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[35],stage1_15[36],stage1_14[42],stage1_13[66]}
   );
   gpc606_5 gpc196 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[36],stage1_15[37],stage1_14[43],stage1_13[67]}
   );
   gpc606_5 gpc197 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[37],stage1_15[38],stage1_14[44],stage1_13[68]}
   );
   gpc606_5 gpc198 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[38],stage1_15[39],stage1_14[45],stage1_13[69]}
   );
   gpc606_5 gpc199 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[39],stage1_15[40],stage1_14[46],stage1_13[70]}
   );
   gpc606_5 gpc200 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[40],stage1_15[41],stage1_14[47],stage1_13[71]}
   );
   gpc606_5 gpc201 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[41],stage1_15[42],stage1_14[48],stage1_13[72]}
   );
   gpc606_5 gpc202 (
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[42],stage1_15[43],stage1_14[49],stage1_13[73]}
   );
   gpc606_5 gpc203 (
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[43],stage1_15[44],stage1_14[50],stage1_13[74]}
   );
   gpc606_5 gpc204 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[44],stage1_15[45],stage1_14[51],stage1_13[75]}
   );
   gpc606_5 gpc205 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[45],stage1_15[46],stage1_14[52],stage1_13[76]}
   );
   gpc606_5 gpc206 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[46],stage1_15[47],stage1_14[53],stage1_13[77]}
   );
   gpc117_4 gpc207 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[156]},
      {1'b0},
      {stage1_17[26],stage1_16[47],stage1_15[48],stage1_14[54]}
   );
   gpc117_4 gpc208 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage0_15[157]},
      {1'b0},
      {stage1_17[27],stage1_16[48],stage1_15[49],stage1_14[55]}
   );
   gpc1_1 gpc209 (
      {stage0_0[160]},
      {stage1_0[31]}
   );
   gpc1_1 gpc210 (
      {stage0_0[161]},
      {stage1_0[32]}
   );
   gpc1_1 gpc211 (
      {stage0_2[152]},
      {stage1_2[54]}
   );
   gpc1_1 gpc212 (
      {stage0_2[153]},
      {stage1_2[55]}
   );
   gpc1_1 gpc213 (
      {stage0_2[154]},
      {stage1_2[56]}
   );
   gpc1_1 gpc214 (
      {stage0_2[155]},
      {stage1_2[57]}
   );
   gpc1_1 gpc215 (
      {stage0_2[156]},
      {stage1_2[58]}
   );
   gpc1_1 gpc216 (
      {stage0_2[157]},
      {stage1_2[59]}
   );
   gpc1_1 gpc217 (
      {stage0_2[158]},
      {stage1_2[60]}
   );
   gpc1_1 gpc218 (
      {stage0_2[159]},
      {stage1_2[61]}
   );
   gpc1_1 gpc219 (
      {stage0_2[160]},
      {stage1_2[62]}
   );
   gpc1_1 gpc220 (
      {stage0_2[161]},
      {stage1_2[63]}
   );
   gpc1_1 gpc221 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc222 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc223 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc224 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc225 (
      {stage0_3[128]},
      {stage1_3[58]}
   );
   gpc1_1 gpc226 (
      {stage0_3[129]},
      {stage1_3[59]}
   );
   gpc1_1 gpc227 (
      {stage0_3[130]},
      {stage1_3[60]}
   );
   gpc1_1 gpc228 (
      {stage0_3[131]},
      {stage1_3[61]}
   );
   gpc1_1 gpc229 (
      {stage0_3[132]},
      {stage1_3[62]}
   );
   gpc1_1 gpc230 (
      {stage0_3[133]},
      {stage1_3[63]}
   );
   gpc1_1 gpc231 (
      {stage0_3[134]},
      {stage1_3[64]}
   );
   gpc1_1 gpc232 (
      {stage0_3[135]},
      {stage1_3[65]}
   );
   gpc1_1 gpc233 (
      {stage0_3[136]},
      {stage1_3[66]}
   );
   gpc1_1 gpc234 (
      {stage0_3[137]},
      {stage1_3[67]}
   );
   gpc1_1 gpc235 (
      {stage0_3[138]},
      {stage1_3[68]}
   );
   gpc1_1 gpc236 (
      {stage0_3[139]},
      {stage1_3[69]}
   );
   gpc1_1 gpc237 (
      {stage0_3[140]},
      {stage1_3[70]}
   );
   gpc1_1 gpc238 (
      {stage0_3[141]},
      {stage1_3[71]}
   );
   gpc1_1 gpc239 (
      {stage0_3[142]},
      {stage1_3[72]}
   );
   gpc1_1 gpc240 (
      {stage0_3[143]},
      {stage1_3[73]}
   );
   gpc1_1 gpc241 (
      {stage0_3[144]},
      {stage1_3[74]}
   );
   gpc1_1 gpc242 (
      {stage0_3[145]},
      {stage1_3[75]}
   );
   gpc1_1 gpc243 (
      {stage0_3[146]},
      {stage1_3[76]}
   );
   gpc1_1 gpc244 (
      {stage0_3[147]},
      {stage1_3[77]}
   );
   gpc1_1 gpc245 (
      {stage0_3[148]},
      {stage1_3[78]}
   );
   gpc1_1 gpc246 (
      {stage0_3[149]},
      {stage1_3[79]}
   );
   gpc1_1 gpc247 (
      {stage0_3[150]},
      {stage1_3[80]}
   );
   gpc1_1 gpc248 (
      {stage0_3[151]},
      {stage1_3[81]}
   );
   gpc1_1 gpc249 (
      {stage0_3[152]},
      {stage1_3[82]}
   );
   gpc1_1 gpc250 (
      {stage0_3[153]},
      {stage1_3[83]}
   );
   gpc1_1 gpc251 (
      {stage0_3[154]},
      {stage1_3[84]}
   );
   gpc1_1 gpc252 (
      {stage0_3[155]},
      {stage1_3[85]}
   );
   gpc1_1 gpc253 (
      {stage0_3[156]},
      {stage1_3[86]}
   );
   gpc1_1 gpc254 (
      {stage0_3[157]},
      {stage1_3[87]}
   );
   gpc1_1 gpc255 (
      {stage0_3[158]},
      {stage1_3[88]}
   );
   gpc1_1 gpc256 (
      {stage0_3[159]},
      {stage1_3[89]}
   );
   gpc1_1 gpc257 (
      {stage0_3[160]},
      {stage1_3[90]}
   );
   gpc1_1 gpc258 (
      {stage0_3[161]},
      {stage1_3[91]}
   );
   gpc1_1 gpc259 (
      {stage0_8[147]},
      {stage1_8[75]}
   );
   gpc1_1 gpc260 (
      {stage0_8[148]},
      {stage1_8[76]}
   );
   gpc1_1 gpc261 (
      {stage0_8[149]},
      {stage1_8[77]}
   );
   gpc1_1 gpc262 (
      {stage0_8[150]},
      {stage1_8[78]}
   );
   gpc1_1 gpc263 (
      {stage0_8[151]},
      {stage1_8[79]}
   );
   gpc1_1 gpc264 (
      {stage0_8[152]},
      {stage1_8[80]}
   );
   gpc1_1 gpc265 (
      {stage0_8[153]},
      {stage1_8[81]}
   );
   gpc1_1 gpc266 (
      {stage0_8[154]},
      {stage1_8[82]}
   );
   gpc1_1 gpc267 (
      {stage0_8[155]},
      {stage1_8[83]}
   );
   gpc1_1 gpc268 (
      {stage0_8[156]},
      {stage1_8[84]}
   );
   gpc1_1 gpc269 (
      {stage0_8[157]},
      {stage1_8[85]}
   );
   gpc1_1 gpc270 (
      {stage0_8[158]},
      {stage1_8[86]}
   );
   gpc1_1 gpc271 (
      {stage0_8[159]},
      {stage1_8[87]}
   );
   gpc1_1 gpc272 (
      {stage0_8[160]},
      {stage1_8[88]}
   );
   gpc1_1 gpc273 (
      {stage0_8[161]},
      {stage1_8[89]}
   );
   gpc1_1 gpc274 (
      {stage0_9[157]},
      {stage1_9[78]}
   );
   gpc1_1 gpc275 (
      {stage0_9[158]},
      {stage1_9[79]}
   );
   gpc1_1 gpc276 (
      {stage0_9[159]},
      {stage1_9[80]}
   );
   gpc1_1 gpc277 (
      {stage0_9[160]},
      {stage1_9[81]}
   );
   gpc1_1 gpc278 (
      {stage0_9[161]},
      {stage1_9[82]}
   );
   gpc1_1 gpc279 (
      {stage0_10[158]},
      {stage1_10[57]}
   );
   gpc1_1 gpc280 (
      {stage0_10[159]},
      {stage1_10[58]}
   );
   gpc1_1 gpc281 (
      {stage0_10[160]},
      {stage1_10[59]}
   );
   gpc1_1 gpc282 (
      {stage0_10[161]},
      {stage1_10[60]}
   );
   gpc1_1 gpc283 (
      {stage0_11[156]},
      {stage1_11[52]}
   );
   gpc1_1 gpc284 (
      {stage0_11[157]},
      {stage1_11[53]}
   );
   gpc1_1 gpc285 (
      {stage0_11[158]},
      {stage1_11[54]}
   );
   gpc1_1 gpc286 (
      {stage0_11[159]},
      {stage1_11[55]}
   );
   gpc1_1 gpc287 (
      {stage0_11[160]},
      {stage1_11[56]}
   );
   gpc1_1 gpc288 (
      {stage0_11[161]},
      {stage1_11[57]}
   );
   gpc1_1 gpc289 (
      {stage0_14[140]},
      {stage1_14[56]}
   );
   gpc1_1 gpc290 (
      {stage0_14[141]},
      {stage1_14[57]}
   );
   gpc1_1 gpc291 (
      {stage0_14[142]},
      {stage1_14[58]}
   );
   gpc1_1 gpc292 (
      {stage0_14[143]},
      {stage1_14[59]}
   );
   gpc1_1 gpc293 (
      {stage0_14[144]},
      {stage1_14[60]}
   );
   gpc1_1 gpc294 (
      {stage0_14[145]},
      {stage1_14[61]}
   );
   gpc1_1 gpc295 (
      {stage0_14[146]},
      {stage1_14[62]}
   );
   gpc1_1 gpc296 (
      {stage0_14[147]},
      {stage1_14[63]}
   );
   gpc1_1 gpc297 (
      {stage0_14[148]},
      {stage1_14[64]}
   );
   gpc1_1 gpc298 (
      {stage0_14[149]},
      {stage1_14[65]}
   );
   gpc1_1 gpc299 (
      {stage0_14[150]},
      {stage1_14[66]}
   );
   gpc1_1 gpc300 (
      {stage0_14[151]},
      {stage1_14[67]}
   );
   gpc1_1 gpc301 (
      {stage0_14[152]},
      {stage1_14[68]}
   );
   gpc1_1 gpc302 (
      {stage0_14[153]},
      {stage1_14[69]}
   );
   gpc1_1 gpc303 (
      {stage0_14[154]},
      {stage1_14[70]}
   );
   gpc1_1 gpc304 (
      {stage0_14[155]},
      {stage1_14[71]}
   );
   gpc1_1 gpc305 (
      {stage0_14[156]},
      {stage1_14[72]}
   );
   gpc1_1 gpc306 (
      {stage0_14[157]},
      {stage1_14[73]}
   );
   gpc1_1 gpc307 (
      {stage0_14[158]},
      {stage1_14[74]}
   );
   gpc1_1 gpc308 (
      {stage0_14[159]},
      {stage1_14[75]}
   );
   gpc1_1 gpc309 (
      {stage0_14[160]},
      {stage1_14[76]}
   );
   gpc1_1 gpc310 (
      {stage0_14[161]},
      {stage1_14[77]}
   );
   gpc1_1 gpc311 (
      {stage0_15[158]},
      {stage1_15[50]}
   );
   gpc1_1 gpc312 (
      {stage0_15[159]},
      {stage1_15[51]}
   );
   gpc1_1 gpc313 (
      {stage0_15[160]},
      {stage1_15[52]}
   );
   gpc1_1 gpc314 (
      {stage0_15[161]},
      {stage1_15[53]}
   );
   gpc606_5 gpc315 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc316 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc317 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[0]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc318 (
      {stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21]},
      {stage1_1[1]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc319 (
      {stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[2]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc320 (
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc321 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc322 (
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc323 (
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc615_5 gpc324 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34]},
      {stage1_3[24]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc325 (
      {stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage1_3[25]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc326 (
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage1_3[26]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc327 (
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_3[27]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc328 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage1_3[28]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc329 (
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_3[29]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc330 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], 1'b0},
      {stage1_3[30]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc331 (
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc332 (
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc333 (
      {stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc334 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc335 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc336 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[16],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc337 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[17],stage2_4[22],stage2_3[22]}
   );
   gpc615_5 gpc338 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[49]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[14],stage2_5[18],stage2_4[23],stage2_3[23]}
   );
   gpc615_5 gpc339 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[50]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[15],stage2_5[19],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc340 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[51]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[16],stage2_5[20],stage2_4[25],stage2_3[25]}
   );
   gpc606_5 gpc341 (
      {stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[10],stage2_6[17],stage2_5[21],stage2_4[26]}
   );
   gpc606_5 gpc342 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[11],stage2_6[18],stage2_5[22],stage2_4[27]}
   );
   gpc606_5 gpc343 (
      {stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[12],stage2_6[19],stage2_5[23],stage2_4[28]}
   );
   gpc615_5 gpc344 (
      {stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_5[60]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[13],stage2_6[20],stage2_5[24],stage2_4[29]}
   );
   gpc606_5 gpc345 (
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[14],stage2_6[21],stage2_5[25]}
   );
   gpc606_5 gpc346 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[5],stage2_7[15],stage2_6[22]}
   );
   gpc606_5 gpc347 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[6],stage2_7[16],stage2_6[23]}
   );
   gpc606_5 gpc348 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[7],stage2_7[17],stage2_6[24]}
   );
   gpc606_5 gpc349 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[4],stage2_8[8],stage2_7[18],stage2_6[25]}
   );
   gpc615_5 gpc350 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52]},
      {stage1_7[6]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[5],stage2_8[9],stage2_7[19],stage2_6[26]}
   );
   gpc615_5 gpc351 (
      {stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57]},
      {stage1_7[7]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[6],stage2_8[10],stage2_7[20],stage2_6[27]}
   );
   gpc615_5 gpc352 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[7],stage2_8[11],stage2_7[21]}
   );
   gpc615_5 gpc353 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[8],stage2_8[12],stage2_7[22]}
   );
   gpc615_5 gpc354 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[9],stage2_8[13],stage2_7[23]}
   );
   gpc615_5 gpc355 (
      {stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[10],stage2_8[14],stage2_7[24]}
   );
   gpc615_5 gpc356 (
      {stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32]},
      {stage1_8[40]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[10],stage2_9[11],stage2_8[15],stage2_7[25]}
   );
   gpc615_5 gpc357 (
      {stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage1_8[41]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[11],stage2_9[12],stage2_8[16],stage2_7[26]}
   );
   gpc615_5 gpc358 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage1_8[42]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[12],stage2_9[13],stage2_8[17],stage2_7[27]}
   );
   gpc606_5 gpc359 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[7],stage2_10[13],stage2_9[14],stage2_8[18]}
   );
   gpc606_5 gpc360 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[8],stage2_10[14],stage2_9[15],stage2_8[19]}
   );
   gpc606_5 gpc361 (
      {stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[9],stage2_10[15],stage2_9[16],stage2_8[20]}
   );
   gpc606_5 gpc362 (
      {stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[10],stage2_10[16],stage2_9[17],stage2_8[21]}
   );
   gpc606_5 gpc363 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[11],stage2_10[17],stage2_9[18],stage2_8[22]}
   );
   gpc606_5 gpc364 (
      {stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[12],stage2_10[18],stage2_9[19],stage2_8[23]}
   );
   gpc606_5 gpc365 (
      {stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[13],stage2_10[19],stage2_9[20],stage2_8[24]}
   );
   gpc606_5 gpc366 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[7],stage2_11[14],stage2_10[20],stage2_9[21]}
   );
   gpc606_5 gpc367 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[8],stage2_11[15],stage2_10[21],stage2_9[22]}
   );
   gpc615_5 gpc368 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46]},
      {stage1_11[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[9],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc369 (
      {stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51]},
      {stage1_11[13]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[10],stage2_11[17],stage2_10[23]}
   );
   gpc615_5 gpc370 (
      {stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_11[14]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[11],stage2_11[18],stage2_10[24]}
   );
   gpc615_5 gpc371 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], 1'b0},
      {stage1_11[15]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[5],stage2_12[12],stage2_11[19],stage2_10[25]}
   );
   gpc1343_5 gpc372 (
      {stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27]},
      {stage1_13[0], stage1_13[1], stage1_13[2]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[4],stage2_13[6],stage2_12[13],stage2_11[20]}
   );
   gpc615_5 gpc373 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage1_12[28]},
      {stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage2_15[1],stage2_14[5],stage2_13[7],stage2_12[14],stage2_11[21]}
   );
   gpc615_5 gpc374 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[29]},
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage2_15[2],stage2_14[6],stage2_13[8],stage2_12[15],stage2_11[22]}
   );
   gpc615_5 gpc375 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[30]},
      {stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20]},
      {stage2_15[3],stage2_14[7],stage2_13[9],stage2_12[16],stage2_11[23]}
   );
   gpc615_5 gpc376 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[31]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[4],stage2_14[8],stage2_13[10],stage2_12[17],stage2_11[24]}
   );
   gpc615_5 gpc377 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[32]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[5],stage2_14[9],stage2_13[11],stage2_12[18],stage2_11[25]}
   );
   gpc615_5 gpc378 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[33]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[6],stage2_14[10],stage2_13[12],stage2_12[19],stage2_11[26]}
   );
   gpc615_5 gpc379 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[34]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[7],stage2_14[11],stage2_13[13],stage2_12[20],stage2_11[27]}
   );
   gpc615_5 gpc380 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], 1'b0},
      {stage1_12[35]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[8],stage2_14[12],stage2_13[14],stage2_12[21],stage2_11[28]}
   );
   gpc606_5 gpc381 (
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[9],stage2_14[13],stage2_13[15],stage2_12[22]}
   );
   gpc606_5 gpc382 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[10],stage2_14[14],stage2_13[16],stage2_12[23]}
   );
   gpc606_5 gpc383 (
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[11],stage2_14[15],stage2_13[17],stage2_12[24]}
   );
   gpc606_5 gpc384 (
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[12],stage2_14[16],stage2_13[18],stage2_12[25]}
   );
   gpc606_5 gpc385 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[13],stage2_14[17],stage2_13[19],stage2_12[26]}
   );
   gpc606_5 gpc386 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[18],stage2_13[20]}
   );
   gpc606_5 gpc387 (
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[19],stage2_13[21]}
   );
   gpc606_5 gpc388 (
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[20],stage2_13[22]}
   );
   gpc606_5 gpc389 (
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[21],stage2_13[23]}
   );
   gpc606_5 gpc390 (
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[22]}
   );
   gpc606_5 gpc391 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[23]}
   );
   gpc606_5 gpc392 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[24]}
   );
   gpc606_5 gpc393 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[25]}
   );
   gpc606_5 gpc394 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[26]}
   );
   gpc606_5 gpc395 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23],stage2_14[27]}
   );
   gpc606_5 gpc396 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24],stage2_14[28]}
   );
   gpc615_5 gpc397 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[24]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[11],stage2_16[16],stage2_15[25],stage2_14[29]}
   );
   gpc615_5 gpc398 (
      {stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[48]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[8],stage2_17[12],stage2_16[17],stage2_15[26]}
   );
   gpc1_1 gpc399 (
      {stage1_0[27]},
      {stage2_0[5]}
   );
   gpc1_1 gpc400 (
      {stage1_0[28]},
      {stage2_0[6]}
   );
   gpc1_1 gpc401 (
      {stage1_0[29]},
      {stage2_0[7]}
   );
   gpc1_1 gpc402 (
      {stage1_0[30]},
      {stage2_0[8]}
   );
   gpc1_1 gpc403 (
      {stage1_0[31]},
      {stage2_0[9]}
   );
   gpc1_1 gpc404 (
      {stage1_0[32]},
      {stage2_0[10]}
   );
   gpc1_1 gpc405 (
      {stage1_1[27]},
      {stage2_1[9]}
   );
   gpc1_1 gpc406 (
      {stage1_1[28]},
      {stage2_1[10]}
   );
   gpc1_1 gpc407 (
      {stage1_1[29]},
      {stage2_1[11]}
   );
   gpc1_1 gpc408 (
      {stage1_1[30]},
      {stage2_1[12]}
   );
   gpc1_1 gpc409 (
      {stage1_1[31]},
      {stage2_1[13]}
   );
   gpc1_1 gpc410 (
      {stage1_1[32]},
      {stage2_1[14]}
   );
   gpc1_1 gpc411 (
      {stage1_1[33]},
      {stage2_1[15]}
   );
   gpc1_1 gpc412 (
      {stage1_1[34]},
      {stage2_1[16]}
   );
   gpc1_1 gpc413 (
      {stage1_1[35]},
      {stage2_1[17]}
   );
   gpc1_1 gpc414 (
      {stage1_1[36]},
      {stage2_1[18]}
   );
   gpc1_1 gpc415 (
      {stage1_1[37]},
      {stage2_1[19]}
   );
   gpc1_1 gpc416 (
      {stage1_1[38]},
      {stage2_1[20]}
   );
   gpc1_1 gpc417 (
      {stage1_1[39]},
      {stage2_1[21]}
   );
   gpc1_1 gpc418 (
      {stage1_1[40]},
      {stage2_1[22]}
   );
   gpc1_1 gpc419 (
      {stage1_1[41]},
      {stage2_1[23]}
   );
   gpc1_1 gpc420 (
      {stage1_1[42]},
      {stage2_1[24]}
   );
   gpc1_1 gpc421 (
      {stage1_1[43]},
      {stage2_1[25]}
   );
   gpc1_1 gpc422 (
      {stage1_1[44]},
      {stage2_1[26]}
   );
   gpc1_1 gpc423 (
      {stage1_1[45]},
      {stage2_1[27]}
   );
   gpc1_1 gpc424 (
      {stage1_1[46]},
      {stage2_1[28]}
   );
   gpc1_1 gpc425 (
      {stage1_1[47]},
      {stage2_1[29]}
   );
   gpc1_1 gpc426 (
      {stage1_3[81]},
      {stage2_3[26]}
   );
   gpc1_1 gpc427 (
      {stage1_3[82]},
      {stage2_3[27]}
   );
   gpc1_1 gpc428 (
      {stage1_3[83]},
      {stage2_3[28]}
   );
   gpc1_1 gpc429 (
      {stage1_3[84]},
      {stage2_3[29]}
   );
   gpc1_1 gpc430 (
      {stage1_3[85]},
      {stage2_3[30]}
   );
   gpc1_1 gpc431 (
      {stage1_3[86]},
      {stage2_3[31]}
   );
   gpc1_1 gpc432 (
      {stage1_3[87]},
      {stage2_3[32]}
   );
   gpc1_1 gpc433 (
      {stage1_3[88]},
      {stage2_3[33]}
   );
   gpc1_1 gpc434 (
      {stage1_3[89]},
      {stage2_3[34]}
   );
   gpc1_1 gpc435 (
      {stage1_3[90]},
      {stage2_3[35]}
   );
   gpc1_1 gpc436 (
      {stage1_3[91]},
      {stage2_3[36]}
   );
   gpc1_1 gpc437 (
      {stage1_5[67]},
      {stage2_5[26]}
   );
   gpc1_1 gpc438 (
      {stage1_5[68]},
      {stage2_5[27]}
   );
   gpc1_1 gpc439 (
      {stage1_5[69]},
      {stage2_5[28]}
   );
   gpc1_1 gpc440 (
      {stage1_5[70]},
      {stage2_5[29]}
   );
   gpc1_1 gpc441 (
      {stage1_6[58]},
      {stage2_6[28]}
   );
   gpc1_1 gpc442 (
      {stage1_6[59]},
      {stage2_6[29]}
   );
   gpc1_1 gpc443 (
      {stage1_7[43]},
      {stage2_7[28]}
   );
   gpc1_1 gpc444 (
      {stage1_7[44]},
      {stage2_7[29]}
   );
   gpc1_1 gpc445 (
      {stage1_7[45]},
      {stage2_7[30]}
   );
   gpc1_1 gpc446 (
      {stage1_7[46]},
      {stage2_7[31]}
   );
   gpc1_1 gpc447 (
      {stage1_7[47]},
      {stage2_7[32]}
   );
   gpc1_1 gpc448 (
      {stage1_7[48]},
      {stage2_7[33]}
   );
   gpc1_1 gpc449 (
      {stage1_7[49]},
      {stage2_7[34]}
   );
   gpc1_1 gpc450 (
      {stage1_7[50]},
      {stage2_7[35]}
   );
   gpc1_1 gpc451 (
      {stage1_7[51]},
      {stage2_7[36]}
   );
   gpc1_1 gpc452 (
      {stage1_7[52]},
      {stage2_7[37]}
   );
   gpc1_1 gpc453 (
      {stage1_7[53]},
      {stage2_7[38]}
   );
   gpc1_1 gpc454 (
      {stage1_8[85]},
      {stage2_8[25]}
   );
   gpc1_1 gpc455 (
      {stage1_8[86]},
      {stage2_8[26]}
   );
   gpc1_1 gpc456 (
      {stage1_8[87]},
      {stage2_8[27]}
   );
   gpc1_1 gpc457 (
      {stage1_8[88]},
      {stage2_8[28]}
   );
   gpc1_1 gpc458 (
      {stage1_8[89]},
      {stage2_8[29]}
   );
   gpc1_1 gpc459 (
      {stage1_9[54]},
      {stage2_9[23]}
   );
   gpc1_1 gpc460 (
      {stage1_9[55]},
      {stage2_9[24]}
   );
   gpc1_1 gpc461 (
      {stage1_9[56]},
      {stage2_9[25]}
   );
   gpc1_1 gpc462 (
      {stage1_9[57]},
      {stage2_9[26]}
   );
   gpc1_1 gpc463 (
      {stage1_9[58]},
      {stage2_9[27]}
   );
   gpc1_1 gpc464 (
      {stage1_9[59]},
      {stage2_9[28]}
   );
   gpc1_1 gpc465 (
      {stage1_9[60]},
      {stage2_9[29]}
   );
   gpc1_1 gpc466 (
      {stage1_9[61]},
      {stage2_9[30]}
   );
   gpc1_1 gpc467 (
      {stage1_9[62]},
      {stage2_9[31]}
   );
   gpc1_1 gpc468 (
      {stage1_9[63]},
      {stage2_9[32]}
   );
   gpc1_1 gpc469 (
      {stage1_9[64]},
      {stage2_9[33]}
   );
   gpc1_1 gpc470 (
      {stage1_9[65]},
      {stage2_9[34]}
   );
   gpc1_1 gpc471 (
      {stage1_9[66]},
      {stage2_9[35]}
   );
   gpc1_1 gpc472 (
      {stage1_9[67]},
      {stage2_9[36]}
   );
   gpc1_1 gpc473 (
      {stage1_9[68]},
      {stage2_9[37]}
   );
   gpc1_1 gpc474 (
      {stage1_9[69]},
      {stage2_9[38]}
   );
   gpc1_1 gpc475 (
      {stage1_9[70]},
      {stage2_9[39]}
   );
   gpc1_1 gpc476 (
      {stage1_9[71]},
      {stage2_9[40]}
   );
   gpc1_1 gpc477 (
      {stage1_9[72]},
      {stage2_9[41]}
   );
   gpc1_1 gpc478 (
      {stage1_9[73]},
      {stage2_9[42]}
   );
   gpc1_1 gpc479 (
      {stage1_9[74]},
      {stage2_9[43]}
   );
   gpc1_1 gpc480 (
      {stage1_9[75]},
      {stage2_9[44]}
   );
   gpc1_1 gpc481 (
      {stage1_9[76]},
      {stage2_9[45]}
   );
   gpc1_1 gpc482 (
      {stage1_9[77]},
      {stage2_9[46]}
   );
   gpc1_1 gpc483 (
      {stage1_9[78]},
      {stage2_9[47]}
   );
   gpc1_1 gpc484 (
      {stage1_9[79]},
      {stage2_9[48]}
   );
   gpc1_1 gpc485 (
      {stage1_9[80]},
      {stage2_9[49]}
   );
   gpc1_1 gpc486 (
      {stage1_9[81]},
      {stage2_9[50]}
   );
   gpc1_1 gpc487 (
      {stage1_9[82]},
      {stage2_9[51]}
   );
   gpc1_1 gpc488 (
      {stage1_12[66]},
      {stage2_12[27]}
   );
   gpc1_1 gpc489 (
      {stage1_12[67]},
      {stage2_12[28]}
   );
   gpc1_1 gpc490 (
      {stage1_12[68]},
      {stage2_12[29]}
   );
   gpc1_1 gpc491 (
      {stage1_12[69]},
      {stage2_12[30]}
   );
   gpc1_1 gpc492 (
      {stage1_12[70]},
      {stage2_12[31]}
   );
   gpc1_1 gpc493 (
      {stage1_12[71]},
      {stage2_12[32]}
   );
   gpc1_1 gpc494 (
      {stage1_12[72]},
      {stage2_12[33]}
   );
   gpc1_1 gpc495 (
      {stage1_13[75]},
      {stage2_13[24]}
   );
   gpc1_1 gpc496 (
      {stage1_13[76]},
      {stage2_13[25]}
   );
   gpc1_1 gpc497 (
      {stage1_13[77]},
      {stage2_13[26]}
   );
   gpc1_1 gpc498 (
      {stage1_15[30]},
      {stage2_15[27]}
   );
   gpc1_1 gpc499 (
      {stage1_15[31]},
      {stage2_15[28]}
   );
   gpc1_1 gpc500 (
      {stage1_15[32]},
      {stage2_15[29]}
   );
   gpc1_1 gpc501 (
      {stage1_15[33]},
      {stage2_15[30]}
   );
   gpc1_1 gpc502 (
      {stage1_15[34]},
      {stage2_15[31]}
   );
   gpc1_1 gpc503 (
      {stage1_15[35]},
      {stage2_15[32]}
   );
   gpc1_1 gpc504 (
      {stage1_15[36]},
      {stage2_15[33]}
   );
   gpc1_1 gpc505 (
      {stage1_15[37]},
      {stage2_15[34]}
   );
   gpc1_1 gpc506 (
      {stage1_15[38]},
      {stage2_15[35]}
   );
   gpc1_1 gpc507 (
      {stage1_15[39]},
      {stage2_15[36]}
   );
   gpc1_1 gpc508 (
      {stage1_15[40]},
      {stage2_15[37]}
   );
   gpc1_1 gpc509 (
      {stage1_15[41]},
      {stage2_15[38]}
   );
   gpc1_1 gpc510 (
      {stage1_15[42]},
      {stage2_15[39]}
   );
   gpc1_1 gpc511 (
      {stage1_15[43]},
      {stage2_15[40]}
   );
   gpc1_1 gpc512 (
      {stage1_15[44]},
      {stage2_15[41]}
   );
   gpc1_1 gpc513 (
      {stage1_15[45]},
      {stage2_15[42]}
   );
   gpc1_1 gpc514 (
      {stage1_15[46]},
      {stage2_15[43]}
   );
   gpc1_1 gpc515 (
      {stage1_15[47]},
      {stage2_15[44]}
   );
   gpc1_1 gpc516 (
      {stage1_15[48]},
      {stage2_15[45]}
   );
   gpc1_1 gpc517 (
      {stage1_15[49]},
      {stage2_15[46]}
   );
   gpc1_1 gpc518 (
      {stage1_15[50]},
      {stage2_15[47]}
   );
   gpc1_1 gpc519 (
      {stage1_15[51]},
      {stage2_15[48]}
   );
   gpc1_1 gpc520 (
      {stage1_15[52]},
      {stage2_15[49]}
   );
   gpc1_1 gpc521 (
      {stage1_15[53]},
      {stage2_15[50]}
   );
   gpc1_1 gpc522 (
      {stage1_17[6]},
      {stage2_17[13]}
   );
   gpc1_1 gpc523 (
      {stage1_17[7]},
      {stage2_17[14]}
   );
   gpc1_1 gpc524 (
      {stage1_17[8]},
      {stage2_17[15]}
   );
   gpc1_1 gpc525 (
      {stage1_17[9]},
      {stage2_17[16]}
   );
   gpc1_1 gpc526 (
      {stage1_17[10]},
      {stage2_17[17]}
   );
   gpc1_1 gpc527 (
      {stage1_17[11]},
      {stage2_17[18]}
   );
   gpc1_1 gpc528 (
      {stage1_17[12]},
      {stage2_17[19]}
   );
   gpc1_1 gpc529 (
      {stage1_17[13]},
      {stage2_17[20]}
   );
   gpc1_1 gpc530 (
      {stage1_17[14]},
      {stage2_17[21]}
   );
   gpc1_1 gpc531 (
      {stage1_17[15]},
      {stage2_17[22]}
   );
   gpc1_1 gpc532 (
      {stage1_17[16]},
      {stage2_17[23]}
   );
   gpc1_1 gpc533 (
      {stage1_17[17]},
      {stage2_17[24]}
   );
   gpc1_1 gpc534 (
      {stage1_17[18]},
      {stage2_17[25]}
   );
   gpc1_1 gpc535 (
      {stage1_17[19]},
      {stage2_17[26]}
   );
   gpc1_1 gpc536 (
      {stage1_17[20]},
      {stage2_17[27]}
   );
   gpc1_1 gpc537 (
      {stage1_17[21]},
      {stage2_17[28]}
   );
   gpc1_1 gpc538 (
      {stage1_17[22]},
      {stage2_17[29]}
   );
   gpc1_1 gpc539 (
      {stage1_17[23]},
      {stage2_17[30]}
   );
   gpc1_1 gpc540 (
      {stage1_17[24]},
      {stage2_17[31]}
   );
   gpc1_1 gpc541 (
      {stage1_17[25]},
      {stage2_17[32]}
   );
   gpc1_1 gpc542 (
      {stage1_17[26]},
      {stage2_17[33]}
   );
   gpc1_1 gpc543 (
      {stage1_17[27]},
      {stage2_17[34]}
   );
   gpc1163_5 gpc544 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc545 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc546 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc547 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc548 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc615_5 gpc549 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc550 (
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage2_4[1]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc606_5 gpc551 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc552 (
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc553 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[4],stage3_6[4],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc554 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[5],stage3_6[5],stage3_5[8],stage3_4[10]}
   );
   gpc606_5 gpc555 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[4],stage3_7[6],stage3_6[6],stage3_5[9]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[5],stage3_7[7],stage3_6[7],stage3_5[10]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[6],stage3_7[8],stage3_6[8],stage3_5[11]}
   );
   gpc615_5 gpc558 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28]},
      {stage2_7[18]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[7],stage3_7[9],stage3_6[9]}
   );
   gpc615_5 gpc559 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[4],stage3_8[8],stage3_7[10]}
   );
   gpc615_5 gpc560 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[5],stage3_8[9],stage3_7[11]}
   );
   gpc615_5 gpc561 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[6],stage3_8[10],stage3_7[12]}
   );
   gpc615_5 gpc562 (
      {stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[7],stage3_8[11],stage3_7[13]}
   );
   gpc606_5 gpc563 (
      {stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[8],stage3_8[12]}
   );
   gpc606_5 gpc564 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[9],stage3_8[13]}
   );
   gpc606_5 gpc565 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[10],stage3_8[14]}
   );
   gpc606_5 gpc566 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[11]}
   );
   gpc606_5 gpc567 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[12]}
   );
   gpc606_5 gpc568 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[13]}
   );
   gpc615_5 gpc569 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46]},
      {stage2_10[18]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[6],stage3_11[10],stage3_10[11],stage3_9[14]}
   );
   gpc615_5 gpc570 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[7],stage3_11[11],stage3_10[12]}
   );
   gpc615_5 gpc571 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], 1'b0},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[5],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc572 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[6],stage3_12[9]}
   );
   gpc606_5 gpc573 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[2],stage3_14[3],stage3_13[7],stage3_12[10]}
   );
   gpc606_5 gpc574 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[3],stage3_14[4],stage3_13[8],stage3_12[11]}
   );
   gpc606_5 gpc575 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[4],stage3_14[5],stage3_13[9],stage3_12[12]}
   );
   gpc606_5 gpc576 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[5],stage3_14[6],stage3_13[10]}
   );
   gpc606_5 gpc577 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[5],stage3_15[6],stage3_14[7],stage3_13[11]}
   );
   gpc606_5 gpc578 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[6],stage3_15[7],stage3_14[8],stage3_13[12]}
   );
   gpc606_5 gpc579 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[7],stage3_15[8],stage3_14[9]}
   );
   gpc615_5 gpc580 (
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[8],stage3_15[9]}
   );
   gpc615_5 gpc581 (
      {stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[9],stage3_15[10]}
   );
   gpc615_5 gpc582 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[6],stage3_16[10],stage3_15[11]}
   );
   gpc615_5 gpc583 (
      {stage2_15[33], stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[7],stage3_16[11],stage3_15[12]}
   );
   gpc615_5 gpc584 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[8],stage3_16[12],stage3_15[13]}
   );
   gpc615_5 gpc585 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[11]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], 1'b0},
      {stage3_19[5],stage3_18[6],stage3_17[9],stage3_16[13],stage3_15[14]}
   );
   gpc606_5 gpc586 (
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[6],stage3_18[7],stage3_17[10],stage3_16[14]}
   );
   gpc1_1 gpc587 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc588 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc589 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc590 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc591 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc592 (
      {stage2_2[2]},
      {stage3_2[5]}
   );
   gpc1_1 gpc593 (
      {stage2_2[3]},
      {stage3_2[6]}
   );
   gpc1_1 gpc594 (
      {stage2_2[4]},
      {stage3_2[7]}
   );
   gpc1_1 gpc595 (
      {stage2_2[5]},
      {stage3_2[8]}
   );
   gpc1_1 gpc596 (
      {stage2_2[6]},
      {stage3_2[9]}
   );
   gpc1_1 gpc597 (
      {stage2_2[7]},
      {stage3_2[10]}
   );
   gpc1_1 gpc598 (
      {stage2_2[8]},
      {stage3_2[11]}
   );
   gpc1_1 gpc599 (
      {stage2_2[9]},
      {stage3_2[12]}
   );
   gpc1_1 gpc600 (
      {stage2_2[10]},
      {stage3_2[13]}
   );
   gpc1_1 gpc601 (
      {stage2_2[11]},
      {stage3_2[14]}
   );
   gpc1_1 gpc602 (
      {stage2_2[12]},
      {stage3_2[15]}
   );
   gpc1_1 gpc603 (
      {stage2_2[13]},
      {stage3_2[16]}
   );
   gpc1_1 gpc604 (
      {stage2_2[14]},
      {stage3_2[17]}
   );
   gpc1_1 gpc605 (
      {stage2_2[15]},
      {stage3_2[18]}
   );
   gpc1_1 gpc606 (
      {stage2_3[30]},
      {stage3_3[7]}
   );
   gpc1_1 gpc607 (
      {stage2_3[31]},
      {stage3_3[8]}
   );
   gpc1_1 gpc608 (
      {stage2_3[32]},
      {stage3_3[9]}
   );
   gpc1_1 gpc609 (
      {stage2_3[33]},
      {stage3_3[10]}
   );
   gpc1_1 gpc610 (
      {stage2_3[34]},
      {stage3_3[11]}
   );
   gpc1_1 gpc611 (
      {stage2_3[35]},
      {stage3_3[12]}
   );
   gpc1_1 gpc612 (
      {stage2_3[36]},
      {stage3_3[13]}
   );
   gpc1_1 gpc613 (
      {stage2_4[26]},
      {stage3_4[11]}
   );
   gpc1_1 gpc614 (
      {stage2_4[27]},
      {stage3_4[12]}
   );
   gpc1_1 gpc615 (
      {stage2_4[28]},
      {stage3_4[13]}
   );
   gpc1_1 gpc616 (
      {stage2_4[29]},
      {stage3_4[14]}
   );
   gpc1_1 gpc617 (
      {stage2_6[29]},
      {stage3_6[10]}
   );
   gpc1_1 gpc618 (
      {stage2_8[28]},
      {stage3_8[15]}
   );
   gpc1_1 gpc619 (
      {stage2_8[29]},
      {stage3_8[16]}
   );
   gpc1_1 gpc620 (
      {stage2_9[47]},
      {stage3_9[15]}
   );
   gpc1_1 gpc621 (
      {stage2_9[48]},
      {stage3_9[16]}
   );
   gpc1_1 gpc622 (
      {stage2_9[49]},
      {stage3_9[17]}
   );
   gpc1_1 gpc623 (
      {stage2_9[50]},
      {stage3_9[18]}
   );
   gpc1_1 gpc624 (
      {stage2_9[51]},
      {stage3_9[19]}
   );
   gpc1_1 gpc625 (
      {stage2_10[24]},
      {stage3_10[13]}
   );
   gpc1_1 gpc626 (
      {stage2_10[25]},
      {stage3_10[14]}
   );
   gpc1_1 gpc627 (
      {stage2_12[31]},
      {stage3_12[13]}
   );
   gpc1_1 gpc628 (
      {stage2_12[32]},
      {stage3_12[14]}
   );
   gpc1_1 gpc629 (
      {stage2_12[33]},
      {stage3_12[15]}
   );
   gpc1_1 gpc630 (
      {stage2_13[24]},
      {stage3_13[13]}
   );
   gpc1_1 gpc631 (
      {stage2_13[25]},
      {stage3_13[14]}
   );
   gpc1_1 gpc632 (
      {stage2_13[26]},
      {stage3_13[15]}
   );
   gpc1_1 gpc633 (
      {stage2_15[48]},
      {stage3_15[15]}
   );
   gpc1_1 gpc634 (
      {stage2_15[49]},
      {stage3_15[16]}
   );
   gpc1_1 gpc635 (
      {stage2_15[50]},
      {stage3_15[17]}
   );
   gpc1_1 gpc636 (
      {stage2_18[6]},
      {stage3_18[8]}
   );
   gpc1_1 gpc637 (
      {stage2_18[7]},
      {stage3_18[9]}
   );
   gpc1_1 gpc638 (
      {stage2_18[8]},
      {stage3_18[10]}
   );
   gpc1_1 gpc639 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc615_5 gpc640 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc641 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[1]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc615_5 gpc642 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[2],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc643 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[3],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc644 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[2],stage4_6[4]}
   );
   gpc615_5 gpc645 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[3],stage4_6[5]}
   );
   gpc615_5 gpc646 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage3_8[12]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[4]}
   );
   gpc615_5 gpc647 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[13]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc648 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc649 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3],stage4_10[5]}
   );
   gpc606_5 gpc650 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4],stage4_10[6]}
   );
   gpc606_5 gpc651 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc615_5 gpc652 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[0]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[4]}
   );
   gpc615_5 gpc653 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[1]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[5]}
   );
   gpc606_5 gpc654 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[3],stage4_16[3],stage4_15[3],stage4_14[5]}
   );
   gpc1163_5 gpc655 (
      {stage3_16[6], stage3_16[7], stage3_16[8]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[4],stage4_16[4]}
   );
   gpc606_5 gpc656 (
      {stage3_16[9], stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14]},
      {stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[5],stage4_16[5]}
   );
   gpc1_1 gpc657 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc658 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc659 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc660 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc661 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc662 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc663 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc664 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc665 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc666 (
      {stage3_1[2]},
      {stage4_1[2]}
   );
   gpc1_1 gpc667 (
      {stage3_1[3]},
      {stage4_1[3]}
   );
   gpc1_1 gpc668 (
      {stage3_1[4]},
      {stage4_1[4]}
   );
   gpc1_1 gpc669 (
      {stage3_2[10]},
      {stage4_2[2]}
   );
   gpc1_1 gpc670 (
      {stage3_2[11]},
      {stage4_2[3]}
   );
   gpc1_1 gpc671 (
      {stage3_2[12]},
      {stage4_2[4]}
   );
   gpc1_1 gpc672 (
      {stage3_2[13]},
      {stage4_2[5]}
   );
   gpc1_1 gpc673 (
      {stage3_2[14]},
      {stage4_2[6]}
   );
   gpc1_1 gpc674 (
      {stage3_2[15]},
      {stage4_2[7]}
   );
   gpc1_1 gpc675 (
      {stage3_2[16]},
      {stage4_2[8]}
   );
   gpc1_1 gpc676 (
      {stage3_2[17]},
      {stage4_2[9]}
   );
   gpc1_1 gpc677 (
      {stage3_2[18]},
      {stage4_2[10]}
   );
   gpc1_1 gpc678 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc679 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc680 (
      {stage3_4[14]},
      {stage4_4[4]}
   );
   gpc1_1 gpc681 (
      {stage3_6[10]},
      {stage4_6[6]}
   );
   gpc1_1 gpc682 (
      {stage3_7[12]},
      {stage4_7[6]}
   );
   gpc1_1 gpc683 (
      {stage3_7[13]},
      {stage4_7[7]}
   );
   gpc1_1 gpc684 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc685 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc686 (
      {stage3_8[16]},
      {stage4_8[6]}
   );
   gpc1_1 gpc687 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc688 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc689 (
      {stage3_10[12]},
      {stage4_10[7]}
   );
   gpc1_1 gpc690 (
      {stage3_10[13]},
      {stage4_10[8]}
   );
   gpc1_1 gpc691 (
      {stage3_10[14]},
      {stage4_10[9]}
   );
   gpc1_1 gpc692 (
      {stage3_11[6]},
      {stage4_11[5]}
   );
   gpc1_1 gpc693 (
      {stage3_11[7]},
      {stage4_11[6]}
   );
   gpc1_1 gpc694 (
      {stage3_11[8]},
      {stage4_11[7]}
   );
   gpc1_1 gpc695 (
      {stage3_11[9]},
      {stage4_11[8]}
   );
   gpc1_1 gpc696 (
      {stage3_11[10]},
      {stage4_11[9]}
   );
   gpc1_1 gpc697 (
      {stage3_11[11]},
      {stage4_11[10]}
   );
   gpc1_1 gpc698 (
      {stage3_11[12]},
      {stage4_11[11]}
   );
   gpc1_1 gpc699 (
      {stage3_12[12]},
      {stage4_12[3]}
   );
   gpc1_1 gpc700 (
      {stage3_12[13]},
      {stage4_12[4]}
   );
   gpc1_1 gpc701 (
      {stage3_12[14]},
      {stage4_12[5]}
   );
   gpc1_1 gpc702 (
      {stage3_12[15]},
      {stage4_12[6]}
   );
   gpc1_1 gpc703 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc704 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc705 (
      {stage3_17[6]},
      {stage4_17[6]}
   );
   gpc1_1 gpc706 (
      {stage3_17[7]},
      {stage4_17[7]}
   );
   gpc1_1 gpc707 (
      {stage3_17[8]},
      {stage4_17[8]}
   );
   gpc1_1 gpc708 (
      {stage3_17[9]},
      {stage4_17[9]}
   );
   gpc1_1 gpc709 (
      {stage3_17[10]},
      {stage4_17[10]}
   );
   gpc1_1 gpc710 (
      {stage3_18[7]},
      {stage4_18[3]}
   );
   gpc1_1 gpc711 (
      {stage3_18[8]},
      {stage4_18[4]}
   );
   gpc1_1 gpc712 (
      {stage3_18[9]},
      {stage4_18[5]}
   );
   gpc1_1 gpc713 (
      {stage3_18[10]},
      {stage4_18[6]}
   );
   gpc1_1 gpc714 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc715 (
      {stage3_19[2]},
      {stage4_19[3]}
   );
   gpc1_1 gpc716 (
      {stage3_19[3]},
      {stage4_19[4]}
   );
   gpc1_1 gpc717 (
      {stage3_19[4]},
      {stage4_19[5]}
   );
   gpc1_1 gpc718 (
      {stage3_19[5]},
      {stage4_19[6]}
   );
   gpc1_1 gpc719 (
      {stage3_19[6]},
      {stage4_19[7]}
   );
   gpc1_1 gpc720 (
      {stage3_19[7]},
      {stage4_19[8]}
   );
   gpc1_1 gpc721 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc606_5 gpc722 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc615_5 gpc723 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1343_5 gpc724 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0], stage4_8[1], stage4_8[2]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0]}
   );
   gpc1343_5 gpc725 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc1343_5 gpc726 (
      {stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc2116_5 gpc727 (
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9]},
      {stage4_11[3]},
      {stage4_12[1]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc207_4 gpc728 (
      {stage4_11[4], stage4_11[5], stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10]},
      {stage4_13[2], stage4_13[3]},
      {stage5_14[1],stage5_13[2],stage5_12[2],stage5_11[2]}
   );
   gpc623_5 gpc729 (
      {stage4_12[2], stage4_12[3], stage4_12[4]},
      {stage4_13[4], stage4_13[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[3],stage5_12[3]}
   );
   gpc1163_5 gpc730 (
      {stage4_15[0], stage4_15[1], stage4_15[2]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0]},
      {stage4_18[0]},
      {stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1]}
   );
   gpc207_4 gpc731 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6], stage4_17[7]},
      {stage4_19[0], stage4_19[1]},
      {stage5_20[0],stage5_19[1],stage5_18[1],stage5_17[1]}
   );
   gpc1406_5 gpc732 (
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], 1'b0},
      {1'b0},
      {stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[2]}
   );
   gpc1_1 gpc733 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc734 (
      {stage4_2[7]},
      {stage5_2[2]}
   );
   gpc1_1 gpc735 (
      {stage4_2[8]},
      {stage5_2[3]}
   );
   gpc1_1 gpc736 (
      {stage4_2[9]},
      {stage5_2[4]}
   );
   gpc1_1 gpc737 (
      {stage4_2[10]},
      {stage5_2[5]}
   );
   gpc1_1 gpc738 (
      {stage4_4[0]},
      {stage5_4[2]}
   );
   gpc1_1 gpc739 (
      {stage4_4[1]},
      {stage5_4[3]}
   );
   gpc1_1 gpc740 (
      {stage4_4[2]},
      {stage5_4[4]}
   );
   gpc1_1 gpc741 (
      {stage4_4[3]},
      {stage5_4[5]}
   );
   gpc1_1 gpc742 (
      {stage4_4[4]},
      {stage5_4[6]}
   );
   gpc1_1 gpc743 (
      {stage4_5[0]},
      {stage5_5[1]}
   );
   gpc1_1 gpc744 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc745 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc746 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc747 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc748 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc749 (
      {stage4_9[5]},
      {stage5_9[3]}
   );
   gpc1_1 gpc750 (
      {stage4_9[6]},
      {stage5_9[4]}
   );
   gpc1_1 gpc751 (
      {stage4_11[11]},
      {stage5_11[3]}
   );
   gpc1_1 gpc752 (
      {stage4_12[5]},
      {stage5_12[4]}
   );
   gpc1_1 gpc753 (
      {stage4_12[6]},
      {stage5_12[5]}
   );
   gpc1_1 gpc754 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc755 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc756 (
      {stage4_15[3]},
      {stage5_15[2]}
   );
   gpc1_1 gpc757 (
      {stage4_17[8]},
      {stage5_17[2]}
   );
   gpc1_1 gpc758 (
      {stage4_17[9]},
      {stage5_17[3]}
   );
   gpc1_1 gpc759 (
      {stage4_17[10]},
      {stage5_17[4]}
   );
   gpc1_1 gpc760 (
      {stage4_19[2]},
      {stage5_19[3]}
   );
   gpc1_1 gpc761 (
      {stage4_19[3]},
      {stage5_19[4]}
   );
   gpc1_1 gpc762 (
      {stage4_19[4]},
      {stage5_19[5]}
   );
   gpc1_1 gpc763 (
      {stage4_19[5]},
      {stage5_19[6]}
   );
   gpc1_1 gpc764 (
      {stage4_19[6]},
      {stage5_19[7]}
   );
   gpc1_1 gpc765 (
      {stage4_19[7]},
      {stage5_19[8]}
   );
   gpc1_1 gpc766 (
      {stage4_19[8]},
      {stage5_19[9]}
   );
   gpc615_5 gpc767 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc768 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0]},
      {stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc769 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc1163_5 gpc770 (
      {stage5_11[1], stage5_11[2], stage5_11[3]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_13[0]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1343_5 gpc771 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc772 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], 1'b0},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1]}
   );
   gpc1343_5 gpc773 (
      {stage5_18[0], stage5_18[1], stage5_18[2]},
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9]},
      {stage5_20[0], stage5_20[1], 1'b0},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[1]}
   );
   gpc1_1 gpc774 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc775 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc776 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc777 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc778 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc779 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc780 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc781 (
      {stage5_7[1]},
      {stage6_7[1]}
   );
   gpc1_1 gpc782 (
      {stage5_9[4]},
      {stage6_9[1]}
   );
   gpc1_1 gpc783 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc784 (
      {stage5_16[1]},
      {stage6_16[1]}
   );
   gpc1_1 gpc785 (
      {stage5_22[0]},
      {stage6_22[1]}
   );
endmodule
module rowadder2_1_23(input [22:0] src0, input [22:0] src1, output [23:0] dst0);
    wire [22:0] gene;
    wire [22:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[22:20]}),
        .S({1'h0, prop[22:20]})
    );
    assign dst0 = {carryout[22], out[22:0]};
endmodule


module comp2_1test_162_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    reg [15:0] src128;
    reg [15:0] src129;
    reg [15:0] src130;
    reg [15:0] src131;
    reg [15:0] src132;
    reg [15:0] src133;
    reg [15:0] src134;
    reg [15:0] src135;
    reg [15:0] src136;
    reg [15:0] src137;
    reg [15:0] src138;
    reg [15:0] src139;
    reg [15:0] src140;
    reg [15:0] src141;
    reg [15:0] src142;
    reg [15:0] src143;
    reg [15:0] src144;
    reg [15:0] src145;
    reg [15:0] src146;
    reg [15:0] src147;
    reg [15:0] src148;
    reg [15:0] src149;
    reg [15:0] src150;
    reg [15:0] src151;
    reg [15:0] src152;
    reg [15:0] src153;
    reg [15:0] src154;
    reg [15:0] src155;
    reg [15:0] src156;
    reg [15:0] src157;
    reg [15:0] src158;
    reg [15:0] src159;
    reg [15:0] src160;
    reg [15:0] src161;
    reg [23:0] exp;
    wire [23:0] dst;
    assign test = dst == exp;
    compressor2_1_162_16 compressor2_1_162_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .src128(src128),
        .src129(src129),
        .src130(src130),
        .src131(src131),
        .src132(src132),
        .src133(src133),
        .src134(src134),
        .src135(src135),
        .src136(src136),
        .src137(src137),
        .src138(src138),
        .src139(src139),
        .src140(src140),
        .src141(src141),
        .src142(src142),
        .src143(src143),
        .src144(src144),
        .src145(src145),
        .src146(src146),
        .src147(src147),
        .src148(src148),
        .src149(src149),
        .src150(src150),
        .src151(src151),
        .src152(src152),
        .src153(src153),
        .src154(src154),
        .src155(src155),
        .src156(src156),
        .src157(src157),
        .src158(src158),
        .src159(src159),
        .src160(src160),
        .src161(src161),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, src128, src129, src130, src131, src132, src133, src134, src135, src136, src137, src138, src139, src140, src141, src142, src143, src144, src145, src146, src147, src148, src149, src150, src151, src152, src153, src154, src155, src156, src157, src158, src159, src160, src161, dst, exp, test);
        src0 <= 16'h20ad;
        src1 <= 16'h9172;
        src2 <= 16'h6cdc;
        src3 <= 16'ha34f;
        src4 <= 16'h6fea;
        src5 <= 16'hf368;
        src6 <= 16'h44b1;
        src7 <= 16'ha2f1;
        src8 <= 16'he0b0;
        src9 <= 16'hc150;
        src10 <= 16'h4433;
        src11 <= 16'h6e61;
        src12 <= 16'hd4b8;
        src13 <= 16'h9b01;
        src14 <= 16'h7df8;
        src15 <= 16'h4dbf;
        src16 <= 16'hf085;
        src17 <= 16'hee18;
        src18 <= 16'h2070;
        src19 <= 16'h5a24;
        src20 <= 16'h3ded;
        src21 <= 16'h2d21;
        src22 <= 16'hbb20;
        src23 <= 16'h309a;
        src24 <= 16'h767f;
        src25 <= 16'h33d3;
        src26 <= 16'h513e;
        src27 <= 16'hbbb;
        src28 <= 16'h9423;
        src29 <= 16'h3f3d;
        src30 <= 16'hdd10;
        src31 <= 16'h14a;
        src32 <= 16'ha5e5;
        src33 <= 16'hae74;
        src34 <= 16'hb3a3;
        src35 <= 16'he75e;
        src36 <= 16'h43bc;
        src37 <= 16'hcb66;
        src38 <= 16'hfbce;
        src39 <= 16'h6fe9;
        src40 <= 16'h23d3;
        src41 <= 16'hcbdc;
        src42 <= 16'hf922;
        src43 <= 16'h985d;
        src44 <= 16'hc50a;
        src45 <= 16'h335;
        src46 <= 16'h3ad2;
        src47 <= 16'hc2e6;
        src48 <= 16'hba98;
        src49 <= 16'hb3cd;
        src50 <= 16'h4235;
        src51 <= 16'hcbcf;
        src52 <= 16'h450c;
        src53 <= 16'h54e0;
        src54 <= 16'ha82d;
        src55 <= 16'h9df2;
        src56 <= 16'h3d0d;
        src57 <= 16'h790;
        src58 <= 16'h32f4;
        src59 <= 16'hb6e0;
        src60 <= 16'h6935;
        src61 <= 16'h242c;
        src62 <= 16'hccec;
        src63 <= 16'h97b8;
        src64 <= 16'h428f;
        src65 <= 16'h6e77;
        src66 <= 16'h7e59;
        src67 <= 16'h7138;
        src68 <= 16'h3df4;
        src69 <= 16'h7bf0;
        src70 <= 16'hbe8c;
        src71 <= 16'h4e18;
        src72 <= 16'hffb0;
        src73 <= 16'h9481;
        src74 <= 16'h600e;
        src75 <= 16'h3586;
        src76 <= 16'h1a80;
        src77 <= 16'hf131;
        src78 <= 16'h7752;
        src79 <= 16'h46a1;
        src80 <= 16'hb1fc;
        src81 <= 16'h6064;
        src82 <= 16'h4d4b;
        src83 <= 16'hecb5;
        src84 <= 16'hb7fb;
        src85 <= 16'h6a35;
        src86 <= 16'h7efc;
        src87 <= 16'hc79b;
        src88 <= 16'h8d9c;
        src89 <= 16'h5728;
        src90 <= 16'h4a09;
        src91 <= 16'h2823;
        src92 <= 16'hf400;
        src93 <= 16'h89f4;
        src94 <= 16'h3da;
        src95 <= 16'ha13a;
        src96 <= 16'h4cb9;
        src97 <= 16'h57d;
        src98 <= 16'h2cff;
        src99 <= 16'h4219;
        src100 <= 16'hdd57;
        src101 <= 16'h3d48;
        src102 <= 16'hb7e3;
        src103 <= 16'h1c5c;
        src104 <= 16'ha8ba;
        src105 <= 16'h4ddd;
        src106 <= 16'h9c70;
        src107 <= 16'h7a66;
        src108 <= 16'h83a5;
        src109 <= 16'he429;
        src110 <= 16'h75e9;
        src111 <= 16'he7fa;
        src112 <= 16'hbbc3;
        src113 <= 16'h19c0;
        src114 <= 16'h63d9;
        src115 <= 16'h8084;
        src116 <= 16'h7ea8;
        src117 <= 16'hd650;
        src118 <= 16'h24eb;
        src119 <= 16'ha769;
        src120 <= 16'h86dd;
        src121 <= 16'ha410;
        src122 <= 16'h9c58;
        src123 <= 16'h9d2d;
        src124 <= 16'hbf20;
        src125 <= 16'h515;
        src126 <= 16'h2985;
        src127 <= 16'h4ba5;
        src128 <= 16'h7a19;
        src129 <= 16'he849;
        src130 <= 16'h77d3;
        src131 <= 16'he2df;
        src132 <= 16'h5ec8;
        src133 <= 16'h556;
        src134 <= 16'hf2f0;
        src135 <= 16'ha64;
        src136 <= 16'hcf5;
        src137 <= 16'h7453;
        src138 <= 16'h3451;
        src139 <= 16'hfb92;
        src140 <= 16'h9b65;
        src141 <= 16'hca3a;
        src142 <= 16'h99eb;
        src143 <= 16'h8728;
        src144 <= 16'h50d1;
        src145 <= 16'h1f54;
        src146 <= 16'h5a81;
        src147 <= 16'h212d;
        src148 <= 16'h6180;
        src149 <= 16'hfd6f;
        src150 <= 16'h5688;
        src151 <= 16'hab4a;
        src152 <= 16'hab1e;
        src153 <= 16'h6386;
        src154 <= 16'h73bf;
        src155 <= 16'hd4df;
        src156 <= 16'h371;
        src157 <= 16'h1308;
        src158 <= 16'h12cf;
        src159 <= 16'h78ce;
        src160 <= 16'hb1b5;
        src161 <= 16'h7803;
        exp <= 24'h4e8077;
        #1
        src0 <= 16'h6c7d;
        src1 <= 16'h4851;
        src2 <= 16'hb25b;
        src3 <= 16'hb859;
        src4 <= 16'h5811;
        src5 <= 16'hd807;
        src6 <= 16'hc575;
        src7 <= 16'hb114;
        src8 <= 16'ha1ea;
        src9 <= 16'hca0c;
        src10 <= 16'h93e7;
        src11 <= 16'h2145;
        src12 <= 16'h1bef;
        src13 <= 16'hd400;
        src14 <= 16'hd880;
        src15 <= 16'h204d;
        src16 <= 16'h5012;
        src17 <= 16'hc63e;
        src18 <= 16'h1895;
        src19 <= 16'hd8c8;
        src20 <= 16'had3b;
        src21 <= 16'h3480;
        src22 <= 16'he3f;
        src23 <= 16'hd36f;
        src24 <= 16'hc293;
        src25 <= 16'hce32;
        src26 <= 16'h4508;
        src27 <= 16'he9c3;
        src28 <= 16'hd445;
        src29 <= 16'hf334;
        src30 <= 16'h299d;
        src31 <= 16'h9926;
        src32 <= 16'h321b;
        src33 <= 16'h9a52;
        src34 <= 16'h962d;
        src35 <= 16'h5109;
        src36 <= 16'hd687;
        src37 <= 16'h166f;
        src38 <= 16'h6d55;
        src39 <= 16'h8f58;
        src40 <= 16'hf031;
        src41 <= 16'h48e1;
        src42 <= 16'he839;
        src43 <= 16'h2571;
        src44 <= 16'ha075;
        src45 <= 16'hca62;
        src46 <= 16'h2aca;
        src47 <= 16'hc94c;
        src48 <= 16'h28b;
        src49 <= 16'h347c;
        src50 <= 16'hc081;
        src51 <= 16'hc58f;
        src52 <= 16'h7cbd;
        src53 <= 16'h6aa9;
        src54 <= 16'ha667;
        src55 <= 16'hc82;
        src56 <= 16'hdba2;
        src57 <= 16'hab65;
        src58 <= 16'h57e4;
        src59 <= 16'h14f8;
        src60 <= 16'h93a4;
        src61 <= 16'hadbd;
        src62 <= 16'h9e45;
        src63 <= 16'h53bd;
        src64 <= 16'h75b7;
        src65 <= 16'h2aa0;
        src66 <= 16'h890e;
        src67 <= 16'h7fa7;
        src68 <= 16'h87de;
        src69 <= 16'h2dab;
        src70 <= 16'h441b;
        src71 <= 16'h6a39;
        src72 <= 16'h79b4;
        src73 <= 16'h666a;
        src74 <= 16'h42ba;
        src75 <= 16'hc2c2;
        src76 <= 16'h65b6;
        src77 <= 16'h737d;
        src78 <= 16'h2555;
        src79 <= 16'h12f2;
        src80 <= 16'h44d6;
        src81 <= 16'h68f;
        src82 <= 16'h908d;
        src83 <= 16'h25f1;
        src84 <= 16'h6aa0;
        src85 <= 16'h102a;
        src86 <= 16'hebbe;
        src87 <= 16'h9217;
        src88 <= 16'h7297;
        src89 <= 16'h98ee;
        src90 <= 16'h6119;
        src91 <= 16'h3837;
        src92 <= 16'hab;
        src93 <= 16'hb4a3;
        src94 <= 16'h1fa1;
        src95 <= 16'ha003;
        src96 <= 16'hfb11;
        src97 <= 16'h3fec;
        src98 <= 16'h82be;
        src99 <= 16'h76d3;
        src100 <= 16'h974d;
        src101 <= 16'h107b;
        src102 <= 16'hf237;
        src103 <= 16'hdf9c;
        src104 <= 16'hf18d;
        src105 <= 16'h9f5b;
        src106 <= 16'h5da4;
        src107 <= 16'h973f;
        src108 <= 16'h84b6;
        src109 <= 16'h68fa;
        src110 <= 16'h5394;
        src111 <= 16'h1333;
        src112 <= 16'ha7c1;
        src113 <= 16'h2937;
        src114 <= 16'ha657;
        src115 <= 16'h1aba;
        src116 <= 16'h1821;
        src117 <= 16'hec9a;
        src118 <= 16'hf073;
        src119 <= 16'heec2;
        src120 <= 16'ha660;
        src121 <= 16'h61e0;
        src122 <= 16'hb692;
        src123 <= 16'h98b2;
        src124 <= 16'h2a95;
        src125 <= 16'he070;
        src126 <= 16'h41bd;
        src127 <= 16'h1278;
        src128 <= 16'h653a;
        src129 <= 16'hcf2b;
        src130 <= 16'h8dda;
        src131 <= 16'h9678;
        src132 <= 16'h2732;
        src133 <= 16'h39ba;
        src134 <= 16'he999;
        src135 <= 16'hd3af;
        src136 <= 16'hdf47;
        src137 <= 16'ha690;
        src138 <= 16'h362d;
        src139 <= 16'h9fdb;
        src140 <= 16'h7fd1;
        src141 <= 16'hf255;
        src142 <= 16'h74be;
        src143 <= 16'ha539;
        src144 <= 16'h78a4;
        src145 <= 16'h4dd3;
        src146 <= 16'h9630;
        src147 <= 16'h98dc;
        src148 <= 16'hdaf9;
        src149 <= 16'h1250;
        src150 <= 16'hba3c;
        src151 <= 16'h8e4f;
        src152 <= 16'hb0a0;
        src153 <= 16'ha394;
        src154 <= 16'h353b;
        src155 <= 16'h3e13;
        src156 <= 16'h8538;
        src157 <= 16'hbef;
        src158 <= 16'h455a;
        src159 <= 16'h9e60;
        src160 <= 16'hbbeb;
        src161 <= 16'h9173;
        exp <= 24'h5087e5;
        #1
        src0 <= 16'h6ce9;
        src1 <= 16'h55fc;
        src2 <= 16'hd503;
        src3 <= 16'h2db2;
        src4 <= 16'h666c;
        src5 <= 16'h262;
        src6 <= 16'h8e40;
        src7 <= 16'h5c62;
        src8 <= 16'hc1c2;
        src9 <= 16'h45f7;
        src10 <= 16'h3bc5;
        src11 <= 16'h5a6a;
        src12 <= 16'ha4cf;
        src13 <= 16'hf436;
        src14 <= 16'hf3e5;
        src15 <= 16'h807f;
        src16 <= 16'h3881;
        src17 <= 16'h225d;
        src18 <= 16'h7ffa;
        src19 <= 16'h8d4f;
        src20 <= 16'he0fa;
        src21 <= 16'h712f;
        src22 <= 16'h2ee;
        src23 <= 16'habb7;
        src24 <= 16'h4852;
        src25 <= 16'heee3;
        src26 <= 16'h8836;
        src27 <= 16'hb068;
        src28 <= 16'h3b1f;
        src29 <= 16'hb4ea;
        src30 <= 16'h1ac0;
        src31 <= 16'h6675;
        src32 <= 16'h5927;
        src33 <= 16'h4ca3;
        src34 <= 16'h43b8;
        src35 <= 16'h6424;
        src36 <= 16'h86a7;
        src37 <= 16'hbe0c;
        src38 <= 16'h7425;
        src39 <= 16'h6879;
        src40 <= 16'hc95a;
        src41 <= 16'h5b2e;
        src42 <= 16'hc6e0;
        src43 <= 16'h2383;
        src44 <= 16'h6bd4;
        src45 <= 16'h5912;
        src46 <= 16'he980;
        src47 <= 16'h398f;
        src48 <= 16'h21b6;
        src49 <= 16'hb6b9;
        src50 <= 16'hd12;
        src51 <= 16'h20c5;
        src52 <= 16'h8c2a;
        src53 <= 16'h4d27;
        src54 <= 16'he3d8;
        src55 <= 16'h560b;
        src56 <= 16'h62d7;
        src57 <= 16'hedbe;
        src58 <= 16'he6e7;
        src59 <= 16'h8caf;
        src60 <= 16'hece1;
        src61 <= 16'h2c2;
        src62 <= 16'h22b4;
        src63 <= 16'h8942;
        src64 <= 16'hfc73;
        src65 <= 16'h1964;
        src66 <= 16'h4081;
        src67 <= 16'h90e6;
        src68 <= 16'hf499;
        src69 <= 16'he386;
        src70 <= 16'h133b;
        src71 <= 16'h2093;
        src72 <= 16'h4e55;
        src73 <= 16'h9fe4;
        src74 <= 16'h1817;
        src75 <= 16'heb25;
        src76 <= 16'hc921;
        src77 <= 16'hb713;
        src78 <= 16'hffde;
        src79 <= 16'h8a27;
        src80 <= 16'h9a67;
        src81 <= 16'hdb3b;
        src82 <= 16'h162b;
        src83 <= 16'hd202;
        src84 <= 16'h7342;
        src85 <= 16'hb632;
        src86 <= 16'hef0a;
        src87 <= 16'h390f;
        src88 <= 16'ha167;
        src89 <= 16'h4dd3;
        src90 <= 16'hd9b7;
        src91 <= 16'hbd86;
        src92 <= 16'hd66b;
        src93 <= 16'ha795;
        src94 <= 16'h730f;
        src95 <= 16'h3613;
        src96 <= 16'hfffe;
        src97 <= 16'hcfc6;
        src98 <= 16'hb898;
        src99 <= 16'h1712;
        src100 <= 16'h64ff;
        src101 <= 16'h6f43;
        src102 <= 16'h76d1;
        src103 <= 16'hf659;
        src104 <= 16'h6562;
        src105 <= 16'h564d;
        src106 <= 16'h81ea;
        src107 <= 16'ha9b7;
        src108 <= 16'hcb7c;
        src109 <= 16'hbfff;
        src110 <= 16'h9d6c;
        src111 <= 16'hfeed;
        src112 <= 16'h8866;
        src113 <= 16'h277c;
        src114 <= 16'h8c4;
        src115 <= 16'h824;
        src116 <= 16'h59b9;
        src117 <= 16'ha57a;
        src118 <= 16'h51e3;
        src119 <= 16'hab5;
        src120 <= 16'hc00d;
        src121 <= 16'hb30a;
        src122 <= 16'h9982;
        src123 <= 16'h2d6a;
        src124 <= 16'h4478;
        src125 <= 16'h743c;
        src126 <= 16'hf4fc;
        src127 <= 16'h4256;
        src128 <= 16'h9648;
        src129 <= 16'h1de1;
        src130 <= 16'ha9b;
        src131 <= 16'h1976;
        src132 <= 16'he9d4;
        src133 <= 16'h64c7;
        src134 <= 16'hf94d;
        src135 <= 16'h936;
        src136 <= 16'hedf6;
        src137 <= 16'hd14f;
        src138 <= 16'hc926;
        src139 <= 16'h4101;
        src140 <= 16'hf6d3;
        src141 <= 16'h4cbf;
        src142 <= 16'hb84e;
        src143 <= 16'h3bf9;
        src144 <= 16'h9b60;
        src145 <= 16'hdbc3;
        src146 <= 16'h4575;
        src147 <= 16'hfd5c;
        src148 <= 16'he744;
        src149 <= 16'h5eb0;
        src150 <= 16'h92d8;
        src151 <= 16'h4a43;
        src152 <= 16'he7cf;
        src153 <= 16'h578;
        src154 <= 16'hfe1b;
        src155 <= 16'hee9a;
        src156 <= 16'hc22d;
        src157 <= 16'h9057;
        src158 <= 16'hd10b;
        src159 <= 16'h7d61;
        src160 <= 16'h1589;
        src161 <= 16'he915;
        exp <= 24'h53f10a;
        #1
        src0 <= 16'h814b;
        src1 <= 16'hb0da;
        src2 <= 16'he9d4;
        src3 <= 16'h5095;
        src4 <= 16'h8d95;
        src5 <= 16'hffa4;
        src6 <= 16'heae;
        src7 <= 16'h178a;
        src8 <= 16'hc4bb;
        src9 <= 16'hd701;
        src10 <= 16'hb51f;
        src11 <= 16'hc3ff;
        src12 <= 16'h27ca;
        src13 <= 16'h7c7;
        src14 <= 16'h988e;
        src15 <= 16'h233a;
        src16 <= 16'hc2;
        src17 <= 16'h7166;
        src18 <= 16'h790c;
        src19 <= 16'h8a59;
        src20 <= 16'h936b;
        src21 <= 16'h8fa9;
        src22 <= 16'h40be;
        src23 <= 16'h282b;
        src24 <= 16'ha876;
        src25 <= 16'hc189;
        src26 <= 16'hd2ec;
        src27 <= 16'h6fc1;
        src28 <= 16'h48a;
        src29 <= 16'hf86b;
        src30 <= 16'hc489;
        src31 <= 16'h5ce;
        src32 <= 16'h401e;
        src33 <= 16'h4fd3;
        src34 <= 16'h1de5;
        src35 <= 16'h9853;
        src36 <= 16'h3cdf;
        src37 <= 16'h34ed;
        src38 <= 16'h41a7;
        src39 <= 16'h6cdb;
        src40 <= 16'he12e;
        src41 <= 16'ha907;
        src42 <= 16'h605d;
        src43 <= 16'he035;
        src44 <= 16'h9297;
        src45 <= 16'h21f;
        src46 <= 16'h82fe;
        src47 <= 16'h9605;
        src48 <= 16'h8624;
        src49 <= 16'hcfc7;
        src50 <= 16'h20a7;
        src51 <= 16'h4514;
        src52 <= 16'hac4c;
        src53 <= 16'h8bb4;
        src54 <= 16'ha0c8;
        src55 <= 16'ha3b4;
        src56 <= 16'h9ee8;
        src57 <= 16'hebd0;
        src58 <= 16'h7105;
        src59 <= 16'h9727;
        src60 <= 16'hfa06;
        src61 <= 16'he4d5;
        src62 <= 16'h1b55;
        src63 <= 16'h7d6e;
        src64 <= 16'had82;
        src65 <= 16'h6484;
        src66 <= 16'hdc8c;
        src67 <= 16'h989f;
        src68 <= 16'h1c50;
        src69 <= 16'h59da;
        src70 <= 16'hd521;
        src71 <= 16'h2dd0;
        src72 <= 16'h1761;
        src73 <= 16'h2477;
        src74 <= 16'h9a1c;
        src75 <= 16'h1ed;
        src76 <= 16'hc228;
        src77 <= 16'h9b29;
        src78 <= 16'h31f2;
        src79 <= 16'h91e1;
        src80 <= 16'h5f8c;
        src81 <= 16'h368c;
        src82 <= 16'h59d3;
        src83 <= 16'h899e;
        src84 <= 16'hcf43;
        src85 <= 16'h35de;
        src86 <= 16'hf20f;
        src87 <= 16'h6b61;
        src88 <= 16'h949c;
        src89 <= 16'hb560;
        src90 <= 16'h595f;
        src91 <= 16'h1fcf;
        src92 <= 16'haff6;
        src93 <= 16'h26e8;
        src94 <= 16'hcf72;
        src95 <= 16'hb7d7;
        src96 <= 16'ha86c;
        src97 <= 16'h314a;
        src98 <= 16'h3f56;
        src99 <= 16'hed96;
        src100 <= 16'h9d26;
        src101 <= 16'h1f62;
        src102 <= 16'h68e4;
        src103 <= 16'h51fd;
        src104 <= 16'h5c81;
        src105 <= 16'hfa9f;
        src106 <= 16'h632b;
        src107 <= 16'hd1e7;
        src108 <= 16'hb034;
        src109 <= 16'hb5ff;
        src110 <= 16'hba02;
        src111 <= 16'h1e7;
        src112 <= 16'h3fc6;
        src113 <= 16'h7a5b;
        src114 <= 16'h8e6b;
        src115 <= 16'h51aa;
        src116 <= 16'h3cce;
        src117 <= 16'h78af;
        src118 <= 16'ha74c;
        src119 <= 16'h2a52;
        src120 <= 16'h2c44;
        src121 <= 16'hc9db;
        src122 <= 16'hfc6e;
        src123 <= 16'h73f8;
        src124 <= 16'hecf3;
        src125 <= 16'h4c6c;
        src126 <= 16'hdc6a;
        src127 <= 16'h21f4;
        src128 <= 16'hbe67;
        src129 <= 16'h7880;
        src130 <= 16'h5bbf;
        src131 <= 16'hf3;
        src132 <= 16'h6377;
        src133 <= 16'he1ca;
        src134 <= 16'hea73;
        src135 <= 16'h843a;
        src136 <= 16'hff7c;
        src137 <= 16'h4594;
        src138 <= 16'hb029;
        src139 <= 16'h4771;
        src140 <= 16'hc94f;
        src141 <= 16'h9f8b;
        src142 <= 16'he530;
        src143 <= 16'hba6f;
        src144 <= 16'h1bd0;
        src145 <= 16'h7359;
        src146 <= 16'h6c7e;
        src147 <= 16'hee22;
        src148 <= 16'h4c8;
        src149 <= 16'h46f2;
        src150 <= 16'h36b6;
        src151 <= 16'heda2;
        src152 <= 16'h248a;
        src153 <= 16'hb99d;
        src154 <= 16'he0a1;
        src155 <= 16'he62;
        src156 <= 16'h6160;
        src157 <= 16'had9b;
        src158 <= 16'hca6a;
        src159 <= 16'h9216;
        src160 <= 16'h762e;
        src161 <= 16'h5f54;
        exp <= 24'h508ea3;
        #1
        src0 <= 16'hcb60;
        src1 <= 16'h6414;
        src2 <= 16'hf7af;
        src3 <= 16'ha961;
        src4 <= 16'hcd14;
        src5 <= 16'hebef;
        src6 <= 16'h1821;
        src7 <= 16'ha289;
        src8 <= 16'h7d56;
        src9 <= 16'hd858;
        src10 <= 16'h4a60;
        src11 <= 16'hd9e7;
        src12 <= 16'h9dab;
        src13 <= 16'h2f2a;
        src14 <= 16'h5fb3;
        src15 <= 16'h1d5e;
        src16 <= 16'h75e2;
        src17 <= 16'h2ace;
        src18 <= 16'h5faf;
        src19 <= 16'hff47;
        src20 <= 16'h26fd;
        src21 <= 16'ha786;
        src22 <= 16'h3d5d;
        src23 <= 16'h1b91;
        src24 <= 16'hc047;
        src25 <= 16'h6a4a;
        src26 <= 16'hbcd7;
        src27 <= 16'hce1a;
        src28 <= 16'h60bc;
        src29 <= 16'h716c;
        src30 <= 16'h23f;
        src31 <= 16'h2268;
        src32 <= 16'h9614;
        src33 <= 16'h44ca;
        src34 <= 16'h1c3e;
        src35 <= 16'h5f1a;
        src36 <= 16'hc5b0;
        src37 <= 16'h73ad;
        src38 <= 16'h8eb3;
        src39 <= 16'h80b6;
        src40 <= 16'h9993;
        src41 <= 16'h9cc4;
        src42 <= 16'hf57e;
        src43 <= 16'h4dc5;
        src44 <= 16'ha8aa;
        src45 <= 16'hbff4;
        src46 <= 16'h13f;
        src47 <= 16'h4448;
        src48 <= 16'hf635;
        src49 <= 16'h3d56;
        src50 <= 16'h9af0;
        src51 <= 16'h45c0;
        src52 <= 16'h82cf;
        src53 <= 16'h79d3;
        src54 <= 16'h29bb;
        src55 <= 16'h9706;
        src56 <= 16'h9920;
        src57 <= 16'h4868;
        src58 <= 16'hc072;
        src59 <= 16'hb5ff;
        src60 <= 16'hef1;
        src61 <= 16'ha102;
        src62 <= 16'h6fbb;
        src63 <= 16'h165d;
        src64 <= 16'h3597;
        src65 <= 16'h20fc;
        src66 <= 16'h7633;
        src67 <= 16'h56dd;
        src68 <= 16'h35f4;
        src69 <= 16'h336e;
        src70 <= 16'h10f8;
        src71 <= 16'hfbac;
        src72 <= 16'he8c4;
        src73 <= 16'h2633;
        src74 <= 16'hd0e9;
        src75 <= 16'ha853;
        src76 <= 16'h5ddd;
        src77 <= 16'h5bfe;
        src78 <= 16'h1c4a;
        src79 <= 16'hbf92;
        src80 <= 16'ha3cc;
        src81 <= 16'hfe89;
        src82 <= 16'hd5d7;
        src83 <= 16'ha35a;
        src84 <= 16'h41f7;
        src85 <= 16'hf3a1;
        src86 <= 16'h3d4d;
        src87 <= 16'hdb56;
        src88 <= 16'heea7;
        src89 <= 16'h94df;
        src90 <= 16'h9f70;
        src91 <= 16'hea58;
        src92 <= 16'h18fe;
        src93 <= 16'h699b;
        src94 <= 16'h2887;
        src95 <= 16'he133;
        src96 <= 16'hc051;
        src97 <= 16'h2388;
        src98 <= 16'ha33f;
        src99 <= 16'hd47d;
        src100 <= 16'hde1a;
        src101 <= 16'hfcd4;
        src102 <= 16'h5a4f;
        src103 <= 16'h572e;
        src104 <= 16'hecec;
        src105 <= 16'hfc50;
        src106 <= 16'he9e7;
        src107 <= 16'hcf18;
        src108 <= 16'ha3d1;
        src109 <= 16'h50d1;
        src110 <= 16'h356d;
        src111 <= 16'h94cf;
        src112 <= 16'h8b5c;
        src113 <= 16'hb7cb;
        src114 <= 16'h64af;
        src115 <= 16'h51a4;
        src116 <= 16'hc647;
        src117 <= 16'he000;
        src118 <= 16'hfa87;
        src119 <= 16'h3bfb;
        src120 <= 16'ha847;
        src121 <= 16'h335f;
        src122 <= 16'hbea1;
        src123 <= 16'h5695;
        src124 <= 16'h529a;
        src125 <= 16'hf993;
        src126 <= 16'hf425;
        src127 <= 16'hcec8;
        src128 <= 16'h9927;
        src129 <= 16'h139d;
        src130 <= 16'hafac;
        src131 <= 16'h723d;
        src132 <= 16'he9b;
        src133 <= 16'h3289;
        src134 <= 16'hffa6;
        src135 <= 16'haa85;
        src136 <= 16'h2374;
        src137 <= 16'hcc37;
        src138 <= 16'he4b0;
        src139 <= 16'h416d;
        src140 <= 16'h57c7;
        src141 <= 16'h2dac;
        src142 <= 16'h73ee;
        src143 <= 16'ha74e;
        src144 <= 16'h3bbb;
        src145 <= 16'hdefb;
        src146 <= 16'h4b11;
        src147 <= 16'h963c;
        src148 <= 16'h1dac;
        src149 <= 16'h53a;
        src150 <= 16'h720b;
        src151 <= 16'hc293;
        src152 <= 16'h2e57;
        src153 <= 16'h991f;
        src154 <= 16'hf30d;
        src155 <= 16'h6117;
        src156 <= 16'hc4cd;
        src157 <= 16'h9591;
        src158 <= 16'h4085;
        src159 <= 16'h70cb;
        src160 <= 16'hdb3c;
        src161 <= 16'h1fe0;
        exp <= 24'h53c276;
        #1
        src0 <= 16'h403d;
        src1 <= 16'h850d;
        src2 <= 16'h78c9;
        src3 <= 16'h9736;
        src4 <= 16'h7afd;
        src5 <= 16'h19f8;
        src6 <= 16'hf0d3;
        src7 <= 16'h9aac;
        src8 <= 16'hd09c;
        src9 <= 16'hc933;
        src10 <= 16'h1b5c;
        src11 <= 16'hb0b5;
        src12 <= 16'h1385;
        src13 <= 16'h6220;
        src14 <= 16'h7491;
        src15 <= 16'hdce8;
        src16 <= 16'ha9c3;
        src17 <= 16'h233;
        src18 <= 16'h7d17;
        src19 <= 16'h4efb;
        src20 <= 16'hde93;
        src21 <= 16'hd7d4;
        src22 <= 16'h1a6;
        src23 <= 16'h1e9;
        src24 <= 16'hd885;
        src25 <= 16'h808d;
        src26 <= 16'hf44c;
        src27 <= 16'h2a6b;
        src28 <= 16'h6af1;
        src29 <= 16'h332b;
        src30 <= 16'h6833;
        src31 <= 16'h6d87;
        src32 <= 16'h6c81;
        src33 <= 16'h2fa4;
        src34 <= 16'hb6d9;
        src35 <= 16'h5fbc;
        src36 <= 16'hca86;
        src37 <= 16'hb6b4;
        src38 <= 16'h9075;
        src39 <= 16'h5bd8;
        src40 <= 16'h5dd8;
        src41 <= 16'hab1b;
        src42 <= 16'hb704;
        src43 <= 16'hdc6b;
        src44 <= 16'hcdc1;
        src45 <= 16'h295;
        src46 <= 16'h352c;
        src47 <= 16'hbd2e;
        src48 <= 16'hb0d2;
        src49 <= 16'h5197;
        src50 <= 16'hd47;
        src51 <= 16'h9586;
        src52 <= 16'h9eef;
        src53 <= 16'hb68;
        src54 <= 16'h8089;
        src55 <= 16'h541c;
        src56 <= 16'h9891;
        src57 <= 16'hb44b;
        src58 <= 16'h1663;
        src59 <= 16'hf132;
        src60 <= 16'hcc87;
        src61 <= 16'h3915;
        src62 <= 16'h311a;
        src63 <= 16'h12ac;
        src64 <= 16'hd5;
        src65 <= 16'hedb6;
        src66 <= 16'h7564;
        src67 <= 16'h4489;
        src68 <= 16'h2455;
        src69 <= 16'he33a;
        src70 <= 16'hf55b;
        src71 <= 16'h9f39;
        src72 <= 16'h6b1;
        src73 <= 16'ha2ce;
        src74 <= 16'hccee;
        src75 <= 16'h775a;
        src76 <= 16'h5696;
        src77 <= 16'h7a04;
        src78 <= 16'h2fbd;
        src79 <= 16'h290f;
        src80 <= 16'he022;
        src81 <= 16'h81e5;
        src82 <= 16'h1af6;
        src83 <= 16'h678e;
        src84 <= 16'h9267;
        src85 <= 16'h7455;
        src86 <= 16'h9511;
        src87 <= 16'h8d71;
        src88 <= 16'h6fb4;
        src89 <= 16'h4483;
        src90 <= 16'he299;
        src91 <= 16'hb02;
        src92 <= 16'hf495;
        src93 <= 16'hbc57;
        src94 <= 16'hf20d;
        src95 <= 16'h9c06;
        src96 <= 16'he109;
        src97 <= 16'h3758;
        src98 <= 16'h5930;
        src99 <= 16'hf8a2;
        src100 <= 16'hba78;
        src101 <= 16'h209d;
        src102 <= 16'h840c;
        src103 <= 16'hd558;
        src104 <= 16'h7d08;
        src105 <= 16'h6bf7;
        src106 <= 16'h645;
        src107 <= 16'h8bba;
        src108 <= 16'hbbc0;
        src109 <= 16'h3b9d;
        src110 <= 16'h2fe4;
        src111 <= 16'hded3;
        src112 <= 16'heacb;
        src113 <= 16'h3277;
        src114 <= 16'hec3d;
        src115 <= 16'ha43;
        src116 <= 16'hf549;
        src117 <= 16'h5c6f;
        src118 <= 16'h7ccb;
        src119 <= 16'hec1e;
        src120 <= 16'h69e0;
        src121 <= 16'hcdd5;
        src122 <= 16'hb659;
        src123 <= 16'h20f4;
        src124 <= 16'h9bc5;
        src125 <= 16'he84f;
        src126 <= 16'hdc1d;
        src127 <= 16'hd809;
        src128 <= 16'h8384;
        src129 <= 16'h329b;
        src130 <= 16'h6c9d;
        src131 <= 16'h8220;
        src132 <= 16'h751b;
        src133 <= 16'h458;
        src134 <= 16'ha50f;
        src135 <= 16'h9572;
        src136 <= 16'h31e9;
        src137 <= 16'hc535;
        src138 <= 16'hbce9;
        src139 <= 16'h8d00;
        src140 <= 16'he0c3;
        src141 <= 16'h14a6;
        src142 <= 16'h150b;
        src143 <= 16'hc70a;
        src144 <= 16'h5054;
        src145 <= 16'h3b2c;
        src146 <= 16'h27ab;
        src147 <= 16'h2e3b;
        src148 <= 16'hb3d5;
        src149 <= 16'h664f;
        src150 <= 16'hb01f;
        src151 <= 16'h675e;
        src152 <= 16'hb0ff;
        src153 <= 16'hf8a3;
        src154 <= 16'h694f;
        src155 <= 16'h6e3f;
        src156 <= 16'h52f3;
        src157 <= 16'h80ec;
        src158 <= 16'h2767;
        src159 <= 16'h81c9;
        src160 <= 16'hf491;
        src161 <= 16'h8950;
        exp <= 24'h50fbeb;
        #1
        src0 <= 16'h483f;
        src1 <= 16'h3022;
        src2 <= 16'h6bc1;
        src3 <= 16'h7c81;
        src4 <= 16'h5b6b;
        src5 <= 16'ha5a3;
        src6 <= 16'h99d5;
        src7 <= 16'h759c;
        src8 <= 16'ha1bb;
        src9 <= 16'h6e12;
        src10 <= 16'h3453;
        src11 <= 16'h19d;
        src12 <= 16'h2af4;
        src13 <= 16'h87d1;
        src14 <= 16'he88d;
        src15 <= 16'hc472;
        src16 <= 16'hd91f;
        src17 <= 16'h7f4c;
        src18 <= 16'hd6c1;
        src19 <= 16'hb62d;
        src20 <= 16'h92a7;
        src21 <= 16'h34ae;
        src22 <= 16'hadab;
        src23 <= 16'h5a3;
        src24 <= 16'h2797;
        src25 <= 16'h5e85;
        src26 <= 16'h140c;
        src27 <= 16'h33cc;
        src28 <= 16'h7c8f;
        src29 <= 16'h8275;
        src30 <= 16'h86ed;
        src31 <= 16'ha7d6;
        src32 <= 16'he66e;
        src33 <= 16'h5cfa;
        src34 <= 16'h73a2;
        src35 <= 16'hae8d;
        src36 <= 16'hc0b2;
        src37 <= 16'h3a4c;
        src38 <= 16'h5be0;
        src39 <= 16'hc8fe;
        src40 <= 16'h5465;
        src41 <= 16'h97e;
        src42 <= 16'ha9f6;
        src43 <= 16'h4ab8;
        src44 <= 16'hc1f9;
        src45 <= 16'h2385;
        src46 <= 16'hb174;
        src47 <= 16'hfc09;
        src48 <= 16'h7d8b;
        src49 <= 16'ha19c;
        src50 <= 16'ha752;
        src51 <= 16'h6392;
        src52 <= 16'h4b6c;
        src53 <= 16'hc855;
        src54 <= 16'hc3e4;
        src55 <= 16'h278f;
        src56 <= 16'h5fa7;
        src57 <= 16'haa63;
        src58 <= 16'h8b0f;
        src59 <= 16'hbc5f;
        src60 <= 16'hbaf6;
        src61 <= 16'hf937;
        src62 <= 16'h971c;
        src63 <= 16'h2d94;
        src64 <= 16'h55da;
        src65 <= 16'h99a5;
        src66 <= 16'h7a6e;
        src67 <= 16'h8763;
        src68 <= 16'hcfa;
        src69 <= 16'hfea8;
        src70 <= 16'ha6d6;
        src71 <= 16'h70b7;
        src72 <= 16'h7552;
        src73 <= 16'h1e22;
        src74 <= 16'h806c;
        src75 <= 16'h7058;
        src76 <= 16'h8e2b;
        src77 <= 16'h3c06;
        src78 <= 16'h8ef9;
        src79 <= 16'hdd18;
        src80 <= 16'h87ad;
        src81 <= 16'hf6ee;
        src82 <= 16'ha678;
        src83 <= 16'h65d6;
        src84 <= 16'h252a;
        src85 <= 16'ha774;
        src86 <= 16'h5dc2;
        src87 <= 16'h7a60;
        src88 <= 16'hc7fe;
        src89 <= 16'hf796;
        src90 <= 16'ha961;
        src91 <= 16'hcfdf;
        src92 <= 16'hcb;
        src93 <= 16'h68d2;
        src94 <= 16'h2b26;
        src95 <= 16'hda0a;
        src96 <= 16'h467c;
        src97 <= 16'hb676;
        src98 <= 16'h58ab;
        src99 <= 16'h7c10;
        src100 <= 16'h918a;
        src101 <= 16'hf9a1;
        src102 <= 16'hae38;
        src103 <= 16'h86ed;
        src104 <= 16'h6336;
        src105 <= 16'hb0eb;
        src106 <= 16'h251f;
        src107 <= 16'h4c07;
        src108 <= 16'h4bec;
        src109 <= 16'hf904;
        src110 <= 16'hca5a;
        src111 <= 16'h6666;
        src112 <= 16'h9d3f;
        src113 <= 16'hc25a;
        src114 <= 16'h8874;
        src115 <= 16'h2dc2;
        src116 <= 16'h3833;
        src117 <= 16'h740a;
        src118 <= 16'h2b88;
        src119 <= 16'h323c;
        src120 <= 16'h95ee;
        src121 <= 16'h7f4d;
        src122 <= 16'hf69c;
        src123 <= 16'had04;
        src124 <= 16'h1578;
        src125 <= 16'h4865;
        src126 <= 16'h66ff;
        src127 <= 16'h9666;
        src128 <= 16'hc4c;
        src129 <= 16'h957f;
        src130 <= 16'hdb7e;
        src131 <= 16'h9639;
        src132 <= 16'h7012;
        src133 <= 16'hec8;
        src134 <= 16'h6891;
        src135 <= 16'hc01f;
        src136 <= 16'he84e;
        src137 <= 16'h3e73;
        src138 <= 16'h3f72;
        src139 <= 16'h9639;
        src140 <= 16'h7021;
        src141 <= 16'h1aaa;
        src142 <= 16'h5376;
        src143 <= 16'h7b7;
        src144 <= 16'h53c1;
        src145 <= 16'h54dd;
        src146 <= 16'h56fe;
        src147 <= 16'h44a0;
        src148 <= 16'hd01;
        src149 <= 16'hb0a9;
        src150 <= 16'h902c;
        src151 <= 16'h7618;
        src152 <= 16'h79c8;
        src153 <= 16'hed11;
        src154 <= 16'hfc5a;
        src155 <= 16'h98d4;
        src156 <= 16'h477;
        src157 <= 16'h7f44;
        src158 <= 16'h77a1;
        src159 <= 16'h5dfc;
        src160 <= 16'hcb6f;
        src161 <= 16'hfd5f;
        exp <= 24'h4ffbd8;
        #1
        src0 <= 16'h580f;
        src1 <= 16'hd5c2;
        src2 <= 16'ha7a5;
        src3 <= 16'h5880;
        src4 <= 16'hc629;
        src5 <= 16'h1444;
        src6 <= 16'hc751;
        src7 <= 16'hba02;
        src8 <= 16'h3fc7;
        src9 <= 16'h5c9e;
        src10 <= 16'ha8ae;
        src11 <= 16'hba7c;
        src12 <= 16'hf703;
        src13 <= 16'h1b13;
        src14 <= 16'hcfbb;
        src15 <= 16'h1a7e;
        src16 <= 16'h1cba;
        src17 <= 16'hcd7b;
        src18 <= 16'h98db;
        src19 <= 16'he797;
        src20 <= 16'h5c35;
        src21 <= 16'hf416;
        src22 <= 16'hcfda;
        src23 <= 16'hb553;
        src24 <= 16'h25d7;
        src25 <= 16'hcbfe;
        src26 <= 16'h8465;
        src27 <= 16'h6a12;
        src28 <= 16'h25cc;
        src29 <= 16'he474;
        src30 <= 16'hee87;
        src31 <= 16'heb07;
        src32 <= 16'h83bf;
        src33 <= 16'h13a0;
        src34 <= 16'hee9f;
        src35 <= 16'h28ca;
        src36 <= 16'h82ea;
        src37 <= 16'h9b37;
        src38 <= 16'h7e0;
        src39 <= 16'h103b;
        src40 <= 16'h5d26;
        src41 <= 16'h7299;
        src42 <= 16'h6649;
        src43 <= 16'h3d65;
        src44 <= 16'hc806;
        src45 <= 16'ha2b7;
        src46 <= 16'h2b2;
        src47 <= 16'h59bf;
        src48 <= 16'h7e24;
        src49 <= 16'h5c57;
        src50 <= 16'hdea3;
        src51 <= 16'h949d;
        src52 <= 16'hfcf2;
        src53 <= 16'h22f3;
        src54 <= 16'h1942;
        src55 <= 16'h26cb;
        src56 <= 16'hd7b0;
        src57 <= 16'h1191;
        src58 <= 16'h1c35;
        src59 <= 16'h3f7c;
        src60 <= 16'hf9be;
        src61 <= 16'hf662;
        src62 <= 16'hb110;
        src63 <= 16'h295b;
        src64 <= 16'h7ad7;
        src65 <= 16'he173;
        src66 <= 16'h6fa6;
        src67 <= 16'h1ef6;
        src68 <= 16'hd9ad;
        src69 <= 16'hc440;
        src70 <= 16'hc3c7;
        src71 <= 16'h2191;
        src72 <= 16'hf0db;
        src73 <= 16'h48d6;
        src74 <= 16'h3c11;
        src75 <= 16'h695d;
        src76 <= 16'h417c;
        src77 <= 16'hba19;
        src78 <= 16'hb2bb;
        src79 <= 16'h97cb;
        src80 <= 16'hf2fd;
        src81 <= 16'h86dc;
        src82 <= 16'h75f5;
        src83 <= 16'h264;
        src84 <= 16'h582a;
        src85 <= 16'h17bd;
        src86 <= 16'h7baf;
        src87 <= 16'h481;
        src88 <= 16'h389e;
        src89 <= 16'h4753;
        src90 <= 16'h7c27;
        src91 <= 16'h7083;
        src92 <= 16'ha806;
        src93 <= 16'h75a9;
        src94 <= 16'h7ff3;
        src95 <= 16'h6786;
        src96 <= 16'he784;
        src97 <= 16'h1396;
        src98 <= 16'hf1;
        src99 <= 16'hc3da;
        src100 <= 16'h6fe1;
        src101 <= 16'h4523;
        src102 <= 16'h6619;
        src103 <= 16'h9489;
        src104 <= 16'h9f18;
        src105 <= 16'h69c0;
        src106 <= 16'ha123;
        src107 <= 16'hc7d1;
        src108 <= 16'h88d6;
        src109 <= 16'h2347;
        src110 <= 16'h8b0b;
        src111 <= 16'h37a1;
        src112 <= 16'hb7;
        src113 <= 16'h524d;
        src114 <= 16'hecd;
        src115 <= 16'h738a;
        src116 <= 16'h254;
        src117 <= 16'hf0c8;
        src118 <= 16'h7f99;
        src119 <= 16'h5977;
        src120 <= 16'h1374;
        src121 <= 16'hafa4;
        src122 <= 16'h6a4d;
        src123 <= 16'hf76;
        src124 <= 16'h2b2e;
        src125 <= 16'hbca9;
        src126 <= 16'hfc12;
        src127 <= 16'hd094;
        src128 <= 16'h8eca;
        src129 <= 16'hdc3b;
        src130 <= 16'he7cc;
        src131 <= 16'h3edd;
        src132 <= 16'he0e5;
        src133 <= 16'h5425;
        src134 <= 16'hde46;
        src135 <= 16'hfe05;
        src136 <= 16'hfd2e;
        src137 <= 16'h615a;
        src138 <= 16'h41d0;
        src139 <= 16'hc524;
        src140 <= 16'hcc2e;
        src141 <= 16'h473d;
        src142 <= 16'hecad;
        src143 <= 16'hb635;
        src144 <= 16'h417;
        src145 <= 16'ha14a;
        src146 <= 16'h2e18;
        src147 <= 16'h7c8d;
        src148 <= 16'ha5ec;
        src149 <= 16'h6853;
        src150 <= 16'hd480;
        src151 <= 16'hb935;
        src152 <= 16'h45d0;
        src153 <= 16'h73a4;
        src154 <= 16'h45b6;
        src155 <= 16'h93da;
        src156 <= 16'ha088;
        src157 <= 16'h509d;
        src158 <= 16'h1680;
        src159 <= 16'hc1d6;
        src160 <= 16'he055;
        src161 <= 16'hc1e1;
        exp <= 24'h50da81;
        #1
        src0 <= 16'hc7e3;
        src1 <= 16'hc4dd;
        src2 <= 16'h7d8d;
        src3 <= 16'h90f6;
        src4 <= 16'hdb8d;
        src5 <= 16'h7aba;
        src6 <= 16'h5ff6;
        src7 <= 16'h6f0f;
        src8 <= 16'h780d;
        src9 <= 16'hd0c1;
        src10 <= 16'hce53;
        src11 <= 16'hf674;
        src12 <= 16'h6443;
        src13 <= 16'h5878;
        src14 <= 16'hae03;
        src15 <= 16'h2ffc;
        src16 <= 16'h3268;
        src17 <= 16'h1b7a;
        src18 <= 16'h4c5d;
        src19 <= 16'hb867;
        src20 <= 16'h836d;
        src21 <= 16'hdbc9;
        src22 <= 16'h330;
        src23 <= 16'hb570;
        src24 <= 16'h6dcf;
        src25 <= 16'hc504;
        src26 <= 16'hf72b;
        src27 <= 16'hb4;
        src28 <= 16'ha3fa;
        src29 <= 16'hf837;
        src30 <= 16'h6f3a;
        src31 <= 16'ha99;
        src32 <= 16'h3b51;
        src33 <= 16'hc143;
        src34 <= 16'h7452;
        src35 <= 16'h8661;
        src36 <= 16'h8f6d;
        src37 <= 16'h1747;
        src38 <= 16'h5d94;
        src39 <= 16'h508;
        src40 <= 16'h181;
        src41 <= 16'h1cb2;
        src42 <= 16'h5683;
        src43 <= 16'hf6d3;
        src44 <= 16'h92d0;
        src45 <= 16'h7ded;
        src46 <= 16'h49bc;
        src47 <= 16'hddc4;
        src48 <= 16'h41c7;
        src49 <= 16'hb3fc;
        src50 <= 16'hcc3f;
        src51 <= 16'h7f5f;
        src52 <= 16'h8f97;
        src53 <= 16'h342e;
        src54 <= 16'hf8d5;
        src55 <= 16'h5032;
        src56 <= 16'h4c22;
        src57 <= 16'hce8c;
        src58 <= 16'h7f37;
        src59 <= 16'h45ea;
        src60 <= 16'h84ea;
        src61 <= 16'h1297;
        src62 <= 16'hd6ee;
        src63 <= 16'h162c;
        src64 <= 16'h1855;
        src65 <= 16'had6e;
        src66 <= 16'h20c8;
        src67 <= 16'h1bff;
        src68 <= 16'h786d;
        src69 <= 16'h6fd7;
        src70 <= 16'h3f31;
        src71 <= 16'h12b5;
        src72 <= 16'h2b14;
        src73 <= 16'h106b;
        src74 <= 16'hebf4;
        src75 <= 16'hc9ee;
        src76 <= 16'hbf1a;
        src77 <= 16'h6f5a;
        src78 <= 16'h61c5;
        src79 <= 16'hb7e2;
        src80 <= 16'hd0e5;
        src81 <= 16'hf1ec;
        src82 <= 16'h4199;
        src83 <= 16'h99a2;
        src84 <= 16'h78ce;
        src85 <= 16'h4f47;
        src86 <= 16'ha15b;
        src87 <= 16'hd382;
        src88 <= 16'ha793;
        src89 <= 16'h673c;
        src90 <= 16'h18d1;
        src91 <= 16'h1fb9;
        src92 <= 16'h537f;
        src93 <= 16'h6d4;
        src94 <= 16'hbdb5;
        src95 <= 16'h98ca;
        src96 <= 16'h42d3;
        src97 <= 16'h324c;
        src98 <= 16'h1f49;
        src99 <= 16'hde0a;
        src100 <= 16'h5f19;
        src101 <= 16'hf326;
        src102 <= 16'hdca3;
        src103 <= 16'hd03d;
        src104 <= 16'h9204;
        src105 <= 16'h25a9;
        src106 <= 16'h8d09;
        src107 <= 16'h77a0;
        src108 <= 16'h5dfb;
        src109 <= 16'h89a4;
        src110 <= 16'hfff1;
        src111 <= 16'h8038;
        src112 <= 16'h5014;
        src113 <= 16'h31e0;
        src114 <= 16'h81dc;
        src115 <= 16'hd2e4;
        src116 <= 16'hcb7a;
        src117 <= 16'h2fff;
        src118 <= 16'hc99f;
        src119 <= 16'h83b3;
        src120 <= 16'h1c7a;
        src121 <= 16'haa48;
        src122 <= 16'hbe6f;
        src123 <= 16'h7206;
        src124 <= 16'h19fa;
        src125 <= 16'ha4;
        src126 <= 16'hb19d;
        src127 <= 16'h9497;
        src128 <= 16'hbb30;
        src129 <= 16'ha6da;
        src130 <= 16'h1d7e;
        src131 <= 16'h2980;
        src132 <= 16'hddbf;
        src133 <= 16'h9d0f;
        src134 <= 16'h1582;
        src135 <= 16'h3c08;
        src136 <= 16'h962d;
        src137 <= 16'h2b67;
        src138 <= 16'h9617;
        src139 <= 16'h25c4;
        src140 <= 16'hefa0;
        src141 <= 16'h68d;
        src142 <= 16'h5f4f;
        src143 <= 16'h2515;
        src144 <= 16'h9d1e;
        src145 <= 16'hf9c;
        src146 <= 16'hd0b6;
        src147 <= 16'hcc0e;
        src148 <= 16'hba2e;
        src149 <= 16'hcf13;
        src150 <= 16'h4dc9;
        src151 <= 16'h8ac0;
        src152 <= 16'h6d6c;
        src153 <= 16'h586a;
        src154 <= 16'hf7ae;
        src155 <= 16'h74c;
        src156 <= 16'h9b6a;
        src157 <= 16'h481f;
        src158 <= 16'hc12a;
        src159 <= 16'hc93;
        src160 <= 16'h101;
        src161 <= 16'hd299;
        exp <= 24'h4d23ec;
        #1
        src0 <= 16'hff12;
        src1 <= 16'hc082;
        src2 <= 16'h8022;
        src3 <= 16'h6ae9;
        src4 <= 16'h3eaf;
        src5 <= 16'h23fb;
        src6 <= 16'h2d37;
        src7 <= 16'h3dbc;
        src8 <= 16'h6af3;
        src9 <= 16'hc0;
        src10 <= 16'h64b7;
        src11 <= 16'h7dcb;
        src12 <= 16'h7fb1;
        src13 <= 16'h5bd5;
        src14 <= 16'h38a1;
        src15 <= 16'h5082;
        src16 <= 16'hb267;
        src17 <= 16'hda1f;
        src18 <= 16'h2cd4;
        src19 <= 16'he76b;
        src20 <= 16'hf85d;
        src21 <= 16'hfa63;
        src22 <= 16'h16a;
        src23 <= 16'h5669;
        src24 <= 16'h5d74;
        src25 <= 16'h87b2;
        src26 <= 16'hd899;
        src27 <= 16'ha447;
        src28 <= 16'hcb88;
        src29 <= 16'h6142;
        src30 <= 16'ha171;
        src31 <= 16'he748;
        src32 <= 16'h63a5;
        src33 <= 16'h15ac;
        src34 <= 16'h686b;
        src35 <= 16'ha7c;
        src36 <= 16'hec7d;
        src37 <= 16'h7cf9;
        src38 <= 16'h6cd4;
        src39 <= 16'hb8f5;
        src40 <= 16'h930;
        src41 <= 16'h4f56;
        src42 <= 16'he608;
        src43 <= 16'hb1a8;
        src44 <= 16'h79c9;
        src45 <= 16'hc252;
        src46 <= 16'h1229;
        src47 <= 16'he787;
        src48 <= 16'h8f2b;
        src49 <= 16'h79ec;
        src50 <= 16'hab24;
        src51 <= 16'h95b6;
        src52 <= 16'h4427;
        src53 <= 16'h690f;
        src54 <= 16'h1763;
        src55 <= 16'hfddd;
        src56 <= 16'h7ee;
        src57 <= 16'he493;
        src58 <= 16'he85a;
        src59 <= 16'h5100;
        src60 <= 16'h2bf9;
        src61 <= 16'hb27c;
        src62 <= 16'h3ec2;
        src63 <= 16'hb404;
        src64 <= 16'h35d3;
        src65 <= 16'h4c9d;
        src66 <= 16'ha5bf;
        src67 <= 16'hfe93;
        src68 <= 16'hefdc;
        src69 <= 16'h1588;
        src70 <= 16'h5696;
        src71 <= 16'hf31d;
        src72 <= 16'h8478;
        src73 <= 16'hed40;
        src74 <= 16'ha92;
        src75 <= 16'hee47;
        src76 <= 16'h85da;
        src77 <= 16'h3e6a;
        src78 <= 16'h2983;
        src79 <= 16'hc2d;
        src80 <= 16'h3272;
        src81 <= 16'hc5d3;
        src82 <= 16'h1b4d;
        src83 <= 16'h6d28;
        src84 <= 16'h2356;
        src85 <= 16'he457;
        src86 <= 16'h6abb;
        src87 <= 16'ha07a;
        src88 <= 16'haf3;
        src89 <= 16'h6bbc;
        src90 <= 16'hbac6;
        src91 <= 16'h524d;
        src92 <= 16'h7b90;
        src93 <= 16'hd49e;
        src94 <= 16'hf0e4;
        src95 <= 16'hf589;
        src96 <= 16'h19ae;
        src97 <= 16'h68e8;
        src98 <= 16'ha359;
        src99 <= 16'hd62d;
        src100 <= 16'h6c41;
        src101 <= 16'h1271;
        src102 <= 16'h7e60;
        src103 <= 16'h6e49;
        src104 <= 16'hf554;
        src105 <= 16'h675b;
        src106 <= 16'h9c36;
        src107 <= 16'hd66e;
        src108 <= 16'hf248;
        src109 <= 16'h1ef3;
        src110 <= 16'h80a7;
        src111 <= 16'hb9;
        src112 <= 16'hee19;
        src113 <= 16'h6d22;
        src114 <= 16'hb4ff;
        src115 <= 16'h4bb1;
        src116 <= 16'h66db;
        src117 <= 16'h318;
        src118 <= 16'h47a2;
        src119 <= 16'h63cf;
        src120 <= 16'h9a01;
        src121 <= 16'h5865;
        src122 <= 16'h68c5;
        src123 <= 16'h86dc;
        src124 <= 16'ha0d8;
        src125 <= 16'ha003;
        src126 <= 16'h8a6d;
        src127 <= 16'hbdd5;
        src128 <= 16'h3493;
        src129 <= 16'h5cb1;
        src130 <= 16'h49ef;
        src131 <= 16'h2bde;
        src132 <= 16'h3c80;
        src133 <= 16'h6831;
        src134 <= 16'h4b2;
        src135 <= 16'h1206;
        src136 <= 16'h5b0b;
        src137 <= 16'h59e3;
        src138 <= 16'h87a;
        src139 <= 16'h68ed;
        src140 <= 16'h973;
        src141 <= 16'h8078;
        src142 <= 16'h61fb;
        src143 <= 16'hc163;
        src144 <= 16'h84dd;
        src145 <= 16'h4356;
        src146 <= 16'hecd1;
        src147 <= 16'h6a07;
        src148 <= 16'h1525;
        src149 <= 16'hd0d7;
        src150 <= 16'hdfd9;
        src151 <= 16'h4a12;
        src152 <= 16'h9eaf;
        src153 <= 16'hf374;
        src154 <= 16'h66ab;
        src155 <= 16'hed5f;
        src156 <= 16'h3511;
        src157 <= 16'h55a0;
        src158 <= 16'h1084;
        src159 <= 16'h3a43;
        src160 <= 16'h7eb3;
        src161 <= 16'h6947;
        exp <= 24'h4d09c8;
        #1
        src0 <= 16'hca9a;
        src1 <= 16'hc3c;
        src2 <= 16'ha9b6;
        src3 <= 16'h1f6;
        src4 <= 16'h3471;
        src5 <= 16'h7e02;
        src6 <= 16'h1ecd;
        src7 <= 16'h1a48;
        src8 <= 16'hf3c8;
        src9 <= 16'hc59e;
        src10 <= 16'h7d2b;
        src11 <= 16'h5bc9;
        src12 <= 16'hed00;
        src13 <= 16'h8617;
        src14 <= 16'hf196;
        src15 <= 16'ha382;
        src16 <= 16'h470a;
        src17 <= 16'hf233;
        src18 <= 16'hdec3;
        src19 <= 16'h8410;
        src20 <= 16'h651e;
        src21 <= 16'h5b10;
        src22 <= 16'h380;
        src23 <= 16'hb38e;
        src24 <= 16'h148e;
        src25 <= 16'h6bdf;
        src26 <= 16'he407;
        src27 <= 16'hbc8b;
        src28 <= 16'h6354;
        src29 <= 16'h68bf;
        src30 <= 16'he12e;
        src31 <= 16'h9f89;
        src32 <= 16'h9560;
        src33 <= 16'h84d8;
        src34 <= 16'h9520;
        src35 <= 16'hec66;
        src36 <= 16'h53fc;
        src37 <= 16'h6807;
        src38 <= 16'h5a20;
        src39 <= 16'hc080;
        src40 <= 16'h64ef;
        src41 <= 16'ha6d3;
        src42 <= 16'h1429;
        src43 <= 16'h4fe8;
        src44 <= 16'ha255;
        src45 <= 16'ha176;
        src46 <= 16'hab9b;
        src47 <= 16'h4414;
        src48 <= 16'h4234;
        src49 <= 16'hbd13;
        src50 <= 16'h3915;
        src51 <= 16'h5f3e;
        src52 <= 16'h14a7;
        src53 <= 16'h95c4;
        src54 <= 16'h4816;
        src55 <= 16'h579e;
        src56 <= 16'hadaf;
        src57 <= 16'hff0a;
        src58 <= 16'h7969;
        src59 <= 16'h311b;
        src60 <= 16'h2649;
        src61 <= 16'h4b06;
        src62 <= 16'h2d8c;
        src63 <= 16'hbb80;
        src64 <= 16'h55cb;
        src65 <= 16'ha58e;
        src66 <= 16'h86a9;
        src67 <= 16'hd992;
        src68 <= 16'hc43e;
        src69 <= 16'h3edf;
        src70 <= 16'hfd7e;
        src71 <= 16'hfae0;
        src72 <= 16'hc38b;
        src73 <= 16'h9d92;
        src74 <= 16'he1f1;
        src75 <= 16'h35e2;
        src76 <= 16'h78a3;
        src77 <= 16'hdbef;
        src78 <= 16'he80a;
        src79 <= 16'h5d0a;
        src80 <= 16'h893b;
        src81 <= 16'hd4f8;
        src82 <= 16'h6117;
        src83 <= 16'h1a78;
        src84 <= 16'hc7cb;
        src85 <= 16'hae4a;
        src86 <= 16'hbb94;
        src87 <= 16'he2d4;
        src88 <= 16'hbc11;
        src89 <= 16'h9b3e;
        src90 <= 16'h66f3;
        src91 <= 16'he2b5;
        src92 <= 16'he5b4;
        src93 <= 16'h4795;
        src94 <= 16'h4d14;
        src95 <= 16'h8ce0;
        src96 <= 16'h8119;
        src97 <= 16'h6e75;
        src98 <= 16'h10f6;
        src99 <= 16'h77ec;
        src100 <= 16'h85f;
        src101 <= 16'h78ad;
        src102 <= 16'hc6db;
        src103 <= 16'h9f06;
        src104 <= 16'h7f93;
        src105 <= 16'h47c;
        src106 <= 16'h14d1;
        src107 <= 16'h35f8;
        src108 <= 16'hb4b3;
        src109 <= 16'hfd;
        src110 <= 16'h69e8;
        src111 <= 16'h7e0b;
        src112 <= 16'hb03a;
        src113 <= 16'h2a32;
        src114 <= 16'h42c2;
        src115 <= 16'h4659;
        src116 <= 16'h9179;
        src117 <= 16'ha1e2;
        src118 <= 16'hebe6;
        src119 <= 16'hf876;
        src120 <= 16'h9e2d;
        src121 <= 16'hf4c5;
        src122 <= 16'hb28;
        src123 <= 16'h74f7;
        src124 <= 16'h728;
        src125 <= 16'h1aae;
        src126 <= 16'hfb64;
        src127 <= 16'hc192;
        src128 <= 16'h40c;
        src129 <= 16'h89c5;
        src130 <= 16'hcfe1;
        src131 <= 16'he686;
        src132 <= 16'h57c2;
        src133 <= 16'ha186;
        src134 <= 16'hebff;
        src135 <= 16'hf4d6;
        src136 <= 16'h6829;
        src137 <= 16'hf378;
        src138 <= 16'h8e94;
        src139 <= 16'hbfd7;
        src140 <= 16'h8327;
        src141 <= 16'h6e73;
        src142 <= 16'hd3d9;
        src143 <= 16'h1b00;
        src144 <= 16'h1053;
        src145 <= 16'hf4d1;
        src146 <= 16'hf092;
        src147 <= 16'h3c8e;
        src148 <= 16'h5012;
        src149 <= 16'ha004;
        src150 <= 16'h51f1;
        src151 <= 16'hbb01;
        src152 <= 16'h1761;
        src153 <= 16'he3c6;
        src154 <= 16'hd29;
        src155 <= 16'hff9d;
        src156 <= 16'hae68;
        src157 <= 16'h98e0;
        src158 <= 16'h8a65;
        src159 <= 16'hd9eb;
        src160 <= 16'h781a;
        src161 <= 16'hf2c3;
        exp <= 24'h556234;
        #1
        src0 <= 16'h4584;
        src1 <= 16'h9512;
        src2 <= 16'h159b;
        src3 <= 16'hbbc7;
        src4 <= 16'h4003;
        src5 <= 16'h630c;
        src6 <= 16'h5767;
        src7 <= 16'h6315;
        src8 <= 16'h9948;
        src9 <= 16'h13f1;
        src10 <= 16'h77ad;
        src11 <= 16'hfd5f;
        src12 <= 16'hf962;
        src13 <= 16'h4f6c;
        src14 <= 16'h7a;
        src15 <= 16'ha471;
        src16 <= 16'h226b;
        src17 <= 16'h1c2d;
        src18 <= 16'h32fd;
        src19 <= 16'h955;
        src20 <= 16'h6f09;
        src21 <= 16'h833d;
        src22 <= 16'haa1c;
        src23 <= 16'hf338;
        src24 <= 16'h21a1;
        src25 <= 16'h94f4;
        src26 <= 16'h279;
        src27 <= 16'h5135;
        src28 <= 16'h429b;
        src29 <= 16'h6519;
        src30 <= 16'hcec2;
        src31 <= 16'h8ef;
        src32 <= 16'hdfce;
        src33 <= 16'h7dd6;
        src34 <= 16'ha400;
        src35 <= 16'h97c6;
        src36 <= 16'h632;
        src37 <= 16'h56fe;
        src38 <= 16'hcb89;
        src39 <= 16'he96d;
        src40 <= 16'h96d2;
        src41 <= 16'h115c;
        src42 <= 16'h2b7f;
        src43 <= 16'h23e7;
        src44 <= 16'h8886;
        src45 <= 16'h8a53;
        src46 <= 16'h3e3f;
        src47 <= 16'h60ae;
        src48 <= 16'h8652;
        src49 <= 16'h702b;
        src50 <= 16'h76ff;
        src51 <= 16'h4c57;
        src52 <= 16'h5703;
        src53 <= 16'h8e9a;
        src54 <= 16'hdc7b;
        src55 <= 16'h8aa1;
        src56 <= 16'hd0d0;
        src57 <= 16'hddc7;
        src58 <= 16'he91;
        src59 <= 16'ha562;
        src60 <= 16'hfa00;
        src61 <= 16'h8714;
        src62 <= 16'h441b;
        src63 <= 16'hf5c9;
        src64 <= 16'hcf35;
        src65 <= 16'hdb97;
        src66 <= 16'ha837;
        src67 <= 16'hef52;
        src68 <= 16'h5fb0;
        src69 <= 16'he4d;
        src70 <= 16'h8838;
        src71 <= 16'h5d1a;
        src72 <= 16'h7508;
        src73 <= 16'h9ad8;
        src74 <= 16'h7cdb;
        src75 <= 16'h51c3;
        src76 <= 16'h3c3d;
        src77 <= 16'hb6c;
        src78 <= 16'h897c;
        src79 <= 16'h8ac9;
        src80 <= 16'h8347;
        src81 <= 16'h3ac8;
        src82 <= 16'habd8;
        src83 <= 16'hdbf0;
        src84 <= 16'h64f4;
        src85 <= 16'hd641;
        src86 <= 16'he3c3;
        src87 <= 16'h6ff0;
        src88 <= 16'h3598;
        src89 <= 16'h4e31;
        src90 <= 16'hc0c1;
        src91 <= 16'hfed;
        src92 <= 16'he763;
        src93 <= 16'hfe3e;
        src94 <= 16'haa0b;
        src95 <= 16'ha567;
        src96 <= 16'h4feb;
        src97 <= 16'h4857;
        src98 <= 16'h2411;
        src99 <= 16'ha215;
        src100 <= 16'hecc;
        src101 <= 16'h799a;
        src102 <= 16'h9970;
        src103 <= 16'h2655;
        src104 <= 16'hb651;
        src105 <= 16'hc126;
        src106 <= 16'h34a1;
        src107 <= 16'h98b4;
        src108 <= 16'h8227;
        src109 <= 16'hb3a2;
        src110 <= 16'h8b23;
        src111 <= 16'hb41d;
        src112 <= 16'hd1df;
        src113 <= 16'h2f05;
        src114 <= 16'hf296;
        src115 <= 16'h622f;
        src116 <= 16'h7946;
        src117 <= 16'hd947;
        src118 <= 16'hda60;
        src119 <= 16'hfdf6;
        src120 <= 16'h16d1;
        src121 <= 16'h6987;
        src122 <= 16'hbc03;
        src123 <= 16'h527e;
        src124 <= 16'h15a0;
        src125 <= 16'h375d;
        src126 <= 16'hc82f;
        src127 <= 16'h2d2d;
        src128 <= 16'h8a65;
        src129 <= 16'hff4;
        src130 <= 16'hd827;
        src131 <= 16'hc863;
        src132 <= 16'hc2aa;
        src133 <= 16'h64b8;
        src134 <= 16'h6207;
        src135 <= 16'h91c1;
        src136 <= 16'h5e32;
        src137 <= 16'h86ab;
        src138 <= 16'h9b68;
        src139 <= 16'h3798;
        src140 <= 16'h3b0f;
        src141 <= 16'hbd22;
        src142 <= 16'h56d4;
        src143 <= 16'had2a;
        src144 <= 16'h4c6e;
        src145 <= 16'hfd31;
        src146 <= 16'ha078;
        src147 <= 16'h1a38;
        src148 <= 16'h2f8f;
        src149 <= 16'hf946;
        src150 <= 16'h4912;
        src151 <= 16'hac82;
        src152 <= 16'hcc40;
        src153 <= 16'hbf23;
        src154 <= 16'h23e8;
        src155 <= 16'h267c;
        src156 <= 16'heece;
        src157 <= 16'hb240;
        src158 <= 16'h7cbf;
        src159 <= 16'hbeab;
        src160 <= 16'h6c21;
        src161 <= 16'hc029;
        exp <= 24'h50127e;
        #1
        src0 <= 16'h3e17;
        src1 <= 16'h8669;
        src2 <= 16'h73ef;
        src3 <= 16'hfe22;
        src4 <= 16'hf40f;
        src5 <= 16'he63;
        src6 <= 16'h1bc1;
        src7 <= 16'hd80a;
        src8 <= 16'h7ac2;
        src9 <= 16'h5de6;
        src10 <= 16'h2e0b;
        src11 <= 16'h9007;
        src12 <= 16'h69fe;
        src13 <= 16'h1650;
        src14 <= 16'ha9ef;
        src15 <= 16'h880b;
        src16 <= 16'h3225;
        src17 <= 16'hc0a9;
        src18 <= 16'h781d;
        src19 <= 16'hcf70;
        src20 <= 16'h257;
        src21 <= 16'h91e5;
        src22 <= 16'h4038;
        src23 <= 16'hbf52;
        src24 <= 16'h102d;
        src25 <= 16'h46af;
        src26 <= 16'h601;
        src27 <= 16'hcfc8;
        src28 <= 16'hfd0a;
        src29 <= 16'h9724;
        src30 <= 16'hd1a4;
        src31 <= 16'hec20;
        src32 <= 16'h3527;
        src33 <= 16'hc6e6;
        src34 <= 16'hdc14;
        src35 <= 16'h329;
        src36 <= 16'h352c;
        src37 <= 16'he1f4;
        src38 <= 16'hab75;
        src39 <= 16'h2865;
        src40 <= 16'hee1e;
        src41 <= 16'hc90f;
        src42 <= 16'hdec6;
        src43 <= 16'hf44a;
        src44 <= 16'h5f53;
        src45 <= 16'h7bbd;
        src46 <= 16'h4935;
        src47 <= 16'h8965;
        src48 <= 16'h1011;
        src49 <= 16'ha309;
        src50 <= 16'h3c6f;
        src51 <= 16'h44d8;
        src52 <= 16'hd6d;
        src53 <= 16'h3b2a;
        src54 <= 16'h835;
        src55 <= 16'h981b;
        src56 <= 16'h63f6;
        src57 <= 16'he94d;
        src58 <= 16'h5711;
        src59 <= 16'he875;
        src60 <= 16'h8731;
        src61 <= 16'h2c94;
        src62 <= 16'h3de5;
        src63 <= 16'h55c1;
        src64 <= 16'h3efe;
        src65 <= 16'h8776;
        src66 <= 16'he520;
        src67 <= 16'h53a;
        src68 <= 16'hc683;
        src69 <= 16'hc0dc;
        src70 <= 16'h6d06;
        src71 <= 16'h64e3;
        src72 <= 16'h9c88;
        src73 <= 16'h228f;
        src74 <= 16'h12e8;
        src75 <= 16'hdea8;
        src76 <= 16'h8386;
        src77 <= 16'hcecb;
        src78 <= 16'h5d2e;
        src79 <= 16'h742c;
        src80 <= 16'h6704;
        src81 <= 16'hc463;
        src82 <= 16'h1f1b;
        src83 <= 16'hbfa3;
        src84 <= 16'h16f2;
        src85 <= 16'h29c2;
        src86 <= 16'h1f50;
        src87 <= 16'hfa1e;
        src88 <= 16'hdf74;
        src89 <= 16'hf976;
        src90 <= 16'h7265;
        src91 <= 16'he339;
        src92 <= 16'hb1e0;
        src93 <= 16'hcfec;
        src94 <= 16'hff6b;
        src95 <= 16'ha7c9;
        src96 <= 16'h7c8c;
        src97 <= 16'h625b;
        src98 <= 16'h6fce;
        src99 <= 16'hca88;
        src100 <= 16'h35c1;
        src101 <= 16'h127b;
        src102 <= 16'ha2e5;
        src103 <= 16'hf447;
        src104 <= 16'h3f08;
        src105 <= 16'hdc0c;
        src106 <= 16'hf897;
        src107 <= 16'h8028;
        src108 <= 16'h884;
        src109 <= 16'h10a9;
        src110 <= 16'ha76f;
        src111 <= 16'h5ec3;
        src112 <= 16'h3668;
        src113 <= 16'h1d33;
        src114 <= 16'hd950;
        src115 <= 16'h531b;
        src116 <= 16'hee0c;
        src117 <= 16'hb128;
        src118 <= 16'h1f08;
        src119 <= 16'h414;
        src120 <= 16'h9d5b;
        src121 <= 16'h6565;
        src122 <= 16'ha8c8;
        src123 <= 16'hbe12;
        src124 <= 16'h582b;
        src125 <= 16'h1aab;
        src126 <= 16'h727a;
        src127 <= 16'ha706;
        src128 <= 16'h41f5;
        src129 <= 16'h3fec;
        src130 <= 16'he25d;
        src131 <= 16'h9b26;
        src132 <= 16'ha80a;
        src133 <= 16'hcca4;
        src134 <= 16'h1b98;
        src135 <= 16'hab27;
        src136 <= 16'h3d70;
        src137 <= 16'ha33;
        src138 <= 16'hbb1a;
        src139 <= 16'h32a1;
        src140 <= 16'hac5b;
        src141 <= 16'h5731;
        src142 <= 16'hfed5;
        src143 <= 16'hf6a5;
        src144 <= 16'hd5fc;
        src145 <= 16'h6147;
        src146 <= 16'h88ed;
        src147 <= 16'h9177;
        src148 <= 16'hced8;
        src149 <= 16'h23b8;
        src150 <= 16'h4c6f;
        src151 <= 16'h97b9;
        src152 <= 16'h1870;
        src153 <= 16'h97f9;
        src154 <= 16'h2b55;
        src155 <= 16'h2015;
        src156 <= 16'h6ad8;
        src157 <= 16'h4b3a;
        src158 <= 16'hfa9c;
        src159 <= 16'h50c9;
        src160 <= 16'h142b;
        src161 <= 16'hc5c6;
        exp <= 24'h4f9952;
        #1
        src0 <= 16'hf119;
        src1 <= 16'h6ae2;
        src2 <= 16'hc460;
        src3 <= 16'h8831;
        src4 <= 16'h406a;
        src5 <= 16'hae7b;
        src6 <= 16'ha077;
        src7 <= 16'hb1c5;
        src8 <= 16'h55f5;
        src9 <= 16'h62d1;
        src10 <= 16'h4a69;
        src11 <= 16'h5c4;
        src12 <= 16'he481;
        src13 <= 16'h1a12;
        src14 <= 16'hdeda;
        src15 <= 16'ha427;
        src16 <= 16'hc55a;
        src17 <= 16'hcf76;
        src18 <= 16'hbb7;
        src19 <= 16'he705;
        src20 <= 16'hc79e;
        src21 <= 16'h6685;
        src22 <= 16'h33af;
        src23 <= 16'he755;
        src24 <= 16'hba03;
        src25 <= 16'hf6f7;
        src26 <= 16'h1d56;
        src27 <= 16'ha823;
        src28 <= 16'h369b;
        src29 <= 16'h653e;
        src30 <= 16'h9209;
        src31 <= 16'hd543;
        src32 <= 16'hc083;
        src33 <= 16'hd3f0;
        src34 <= 16'hbefb;
        src35 <= 16'h70d;
        src36 <= 16'h35ed;
        src37 <= 16'h2dc1;
        src38 <= 16'h9e9e;
        src39 <= 16'h60ee;
        src40 <= 16'h543d;
        src41 <= 16'h5dda;
        src42 <= 16'hba6f;
        src43 <= 16'h424a;
        src44 <= 16'h71dc;
        src45 <= 16'h43c9;
        src46 <= 16'ha756;
        src47 <= 16'h8f14;
        src48 <= 16'h1f6f;
        src49 <= 16'h2bc7;
        src50 <= 16'h8bbf;
        src51 <= 16'h220c;
        src52 <= 16'hf2ef;
        src53 <= 16'h352b;
        src54 <= 16'h79ff;
        src55 <= 16'h5b62;
        src56 <= 16'h553;
        src57 <= 16'he15e;
        src58 <= 16'hab45;
        src59 <= 16'h6731;
        src60 <= 16'hc562;
        src61 <= 16'h7fb1;
        src62 <= 16'h49a2;
        src63 <= 16'hcc83;
        src64 <= 16'h4aa4;
        src65 <= 16'hca55;
        src66 <= 16'h4efa;
        src67 <= 16'haabb;
        src68 <= 16'h4c7b;
        src69 <= 16'h82d8;
        src70 <= 16'h55d9;
        src71 <= 16'h677b;
        src72 <= 16'hdd73;
        src73 <= 16'hc8fc;
        src74 <= 16'h9fa1;
        src75 <= 16'he085;
        src76 <= 16'hcbf7;
        src77 <= 16'hd01e;
        src78 <= 16'hb4cb;
        src79 <= 16'h463b;
        src80 <= 16'h80c1;
        src81 <= 16'h37bf;
        src82 <= 16'h792c;
        src83 <= 16'h7c31;
        src84 <= 16'h8f64;
        src85 <= 16'h5784;
        src86 <= 16'h36cc;
        src87 <= 16'hbf07;
        src88 <= 16'hc3ea;
        src89 <= 16'hb57f;
        src90 <= 16'h2871;
        src91 <= 16'h5e92;
        src92 <= 16'hdcd9;
        src93 <= 16'hba8e;
        src94 <= 16'he530;
        src95 <= 16'h8258;
        src96 <= 16'h8942;
        src97 <= 16'h3200;
        src98 <= 16'hb0b1;
        src99 <= 16'h9eb5;
        src100 <= 16'hceae;
        src101 <= 16'h8f6b;
        src102 <= 16'h97a2;
        src103 <= 16'h916e;
        src104 <= 16'hf3db;
        src105 <= 16'h61e7;
        src106 <= 16'hcb47;
        src107 <= 16'h977f;
        src108 <= 16'hedd4;
        src109 <= 16'hea7c;
        src110 <= 16'hcb6d;
        src111 <= 16'hc356;
        src112 <= 16'h33a7;
        src113 <= 16'h8331;
        src114 <= 16'h94;
        src115 <= 16'ha943;
        src116 <= 16'h1268;
        src117 <= 16'h45ec;
        src118 <= 16'hcb0f;
        src119 <= 16'h4bfd;
        src120 <= 16'h9821;
        src121 <= 16'h404b;
        src122 <= 16'h39fd;
        src123 <= 16'h1d94;
        src124 <= 16'h9134;
        src125 <= 16'hd2b8;
        src126 <= 16'hb506;
        src127 <= 16'h138d;
        src128 <= 16'hb0f2;
        src129 <= 16'hc4e8;
        src130 <= 16'hca56;
        src131 <= 16'hfa35;
        src132 <= 16'hd41;
        src133 <= 16'h4e76;
        src134 <= 16'h2ce7;
        src135 <= 16'h6a5e;
        src136 <= 16'h7912;
        src137 <= 16'h4b2b;
        src138 <= 16'hf480;
        src139 <= 16'h1912;
        src140 <= 16'hea04;
        src141 <= 16'h5c25;
        src142 <= 16'h817e;
        src143 <= 16'hf213;
        src144 <= 16'hb0a4;
        src145 <= 16'h8b5a;
        src146 <= 16'h6d8d;
        src147 <= 16'hb230;
        src148 <= 16'h6f6d;
        src149 <= 16'hb35;
        src150 <= 16'hf664;
        src151 <= 16'h3911;
        src152 <= 16'h49df;
        src153 <= 16'hbba3;
        src154 <= 16'hac1;
        src155 <= 16'he0cb;
        src156 <= 16'hd877;
        src157 <= 16'h87bb;
        src158 <= 16'h728b;
        src159 <= 16'h842a;
        src160 <= 16'h1214;
        src161 <= 16'he121;
        exp <= 24'h551cc3;
        #1
        src0 <= 16'hadad;
        src1 <= 16'he0e;
        src2 <= 16'hf7b;
        src3 <= 16'h4770;
        src4 <= 16'h3d84;
        src5 <= 16'hb88e;
        src6 <= 16'h626e;
        src7 <= 16'hc8e7;
        src8 <= 16'hd305;
        src9 <= 16'h79eb;
        src10 <= 16'h749f;
        src11 <= 16'h4947;
        src12 <= 16'haf91;
        src13 <= 16'hc7f9;
        src14 <= 16'hedb0;
        src15 <= 16'h2610;
        src16 <= 16'hff19;
        src17 <= 16'h5d5;
        src18 <= 16'hffa7;
        src19 <= 16'h70a5;
        src20 <= 16'ha977;
        src21 <= 16'h6a36;
        src22 <= 16'h3cdd;
        src23 <= 16'h3f11;
        src24 <= 16'h3c35;
        src25 <= 16'hb8cf;
        src26 <= 16'h6dcc;
        src27 <= 16'hd2f0;
        src28 <= 16'h3c11;
        src29 <= 16'h3040;
        src30 <= 16'hc8cf;
        src31 <= 16'hd195;
        src32 <= 16'h1381;
        src33 <= 16'h112f;
        src34 <= 16'h47fd;
        src35 <= 16'h6be8;
        src36 <= 16'h7daf;
        src37 <= 16'h747c;
        src38 <= 16'h2065;
        src39 <= 16'hb86a;
        src40 <= 16'hb686;
        src41 <= 16'he1b3;
        src42 <= 16'h3404;
        src43 <= 16'h7ee9;
        src44 <= 16'h71cb;
        src45 <= 16'h171c;
        src46 <= 16'hc4e6;
        src47 <= 16'h4249;
        src48 <= 16'hbe4c;
        src49 <= 16'hdd95;
        src50 <= 16'h9ba0;
        src51 <= 16'ha57d;
        src52 <= 16'h522;
        src53 <= 16'hd330;
        src54 <= 16'h73f9;
        src55 <= 16'h2169;
        src56 <= 16'h2746;
        src57 <= 16'hb19d;
        src58 <= 16'h66c8;
        src59 <= 16'he14;
        src60 <= 16'h91f1;
        src61 <= 16'h5877;
        src62 <= 16'hcff9;
        src63 <= 16'h18a;
        src64 <= 16'h14a5;
        src65 <= 16'hb487;
        src66 <= 16'h622f;
        src67 <= 16'h55fa;
        src68 <= 16'hd7e0;
        src69 <= 16'hd170;
        src70 <= 16'hd32b;
        src71 <= 16'h5e08;
        src72 <= 16'hc25b;
        src73 <= 16'h5938;
        src74 <= 16'hab0f;
        src75 <= 16'hc529;
        src76 <= 16'hc56c;
        src77 <= 16'hbc9d;
        src78 <= 16'hb2b8;
        src79 <= 16'h7813;
        src80 <= 16'hcd97;
        src81 <= 16'h7208;
        src82 <= 16'hc6fc;
        src83 <= 16'h2d4b;
        src84 <= 16'h7d4e;
        src85 <= 16'h3b6d;
        src86 <= 16'hbb1b;
        src87 <= 16'h985e;
        src88 <= 16'haa82;
        src89 <= 16'hd410;
        src90 <= 16'ha44a;
        src91 <= 16'h34b7;
        src92 <= 16'h30f7;
        src93 <= 16'hf45f;
        src94 <= 16'h9af9;
        src95 <= 16'hf883;
        src96 <= 16'h8b98;
        src97 <= 16'hb833;
        src98 <= 16'h772d;
        src99 <= 16'hbcde;
        src100 <= 16'h4dd;
        src101 <= 16'h2be9;
        src102 <= 16'he15c;
        src103 <= 16'h2cec;
        src104 <= 16'h61e8;
        src105 <= 16'hbb7e;
        src106 <= 16'h6469;
        src107 <= 16'ha278;
        src108 <= 16'h4af2;
        src109 <= 16'h719f;
        src110 <= 16'h21c2;
        src111 <= 16'h22f8;
        src112 <= 16'ha65f;
        src113 <= 16'h520f;
        src114 <= 16'hce51;
        src115 <= 16'h8278;
        src116 <= 16'h93dc;
        src117 <= 16'ha0cc;
        src118 <= 16'h8b83;
        src119 <= 16'h2e4b;
        src120 <= 16'hc5d;
        src121 <= 16'hf65c;
        src122 <= 16'hd415;
        src123 <= 16'h38e0;
        src124 <= 16'h738d;
        src125 <= 16'h4eac;
        src126 <= 16'h24ff;
        src127 <= 16'ha57;
        src128 <= 16'h9e5;
        src129 <= 16'h5506;
        src130 <= 16'h1caa;
        src131 <= 16'h31a2;
        src132 <= 16'h488a;
        src133 <= 16'hd92f;
        src134 <= 16'h617f;
        src135 <= 16'h29ff;
        src136 <= 16'hc1f8;
        src137 <= 16'h12b6;
        src138 <= 16'h605e;
        src139 <= 16'h460;
        src140 <= 16'h7945;
        src141 <= 16'hcd8e;
        src142 <= 16'h65b7;
        src143 <= 16'haca2;
        src144 <= 16'h3293;
        src145 <= 16'head3;
        src146 <= 16'h1163;
        src147 <= 16'h6fd3;
        src148 <= 16'h3d1d;
        src149 <= 16'h977c;
        src150 <= 16'h586;
        src151 <= 16'h8a1e;
        src152 <= 16'he4fa;
        src153 <= 16'hc4a7;
        src154 <= 16'h943d;
        src155 <= 16'h18af;
        src156 <= 16'h7584;
        src157 <= 16'h76d1;
        src158 <= 16'h1c1a;
        src159 <= 16'h373b;
        src160 <= 16'hae63;
        src161 <= 16'h13b8;
        exp <= 24'h4c2125;
        #1
        src0 <= 16'h6598;
        src1 <= 16'h2318;
        src2 <= 16'hb4a4;
        src3 <= 16'h1a51;
        src4 <= 16'hcf6e;
        src5 <= 16'h7dfb;
        src6 <= 16'hf12c;
        src7 <= 16'h6a3b;
        src8 <= 16'h9974;
        src9 <= 16'hdf25;
        src10 <= 16'h746d;
        src11 <= 16'h3795;
        src12 <= 16'hf05c;
        src13 <= 16'h233a;
        src14 <= 16'h6883;
        src15 <= 16'h78d6;
        src16 <= 16'hda6a;
        src17 <= 16'h65f;
        src18 <= 16'he059;
        src19 <= 16'h5db3;
        src20 <= 16'hd3a3;
        src21 <= 16'h2951;
        src22 <= 16'hbd0c;
        src23 <= 16'he0a6;
        src24 <= 16'ha0cf;
        src25 <= 16'h6be9;
        src26 <= 16'h48d9;
        src27 <= 16'h9131;
        src28 <= 16'h2f67;
        src29 <= 16'h5cf;
        src30 <= 16'h8548;
        src31 <= 16'hbf70;
        src32 <= 16'h5843;
        src33 <= 16'hae8a;
        src34 <= 16'h9d76;
        src35 <= 16'h7f72;
        src36 <= 16'h99d0;
        src37 <= 16'h7831;
        src38 <= 16'hdb14;
        src39 <= 16'hef61;
        src40 <= 16'h4623;
        src41 <= 16'h1e7c;
        src42 <= 16'hc65b;
        src43 <= 16'hddbb;
        src44 <= 16'hdc83;
        src45 <= 16'h8ac3;
        src46 <= 16'hef38;
        src47 <= 16'hd521;
        src48 <= 16'hd3cd;
        src49 <= 16'he95;
        src50 <= 16'hd7c;
        src51 <= 16'h399;
        src52 <= 16'h66cc;
        src53 <= 16'hf7c0;
        src54 <= 16'hf2dd;
        src55 <= 16'h3fda;
        src56 <= 16'hcac0;
        src57 <= 16'h91fd;
        src58 <= 16'h6cb0;
        src59 <= 16'h2807;
        src60 <= 16'h4a;
        src61 <= 16'h6a82;
        src62 <= 16'h6bb9;
        src63 <= 16'hd316;
        src64 <= 16'ha102;
        src65 <= 16'h664c;
        src66 <= 16'h899b;
        src67 <= 16'h80b4;
        src68 <= 16'h5f5d;
        src69 <= 16'ha4ae;
        src70 <= 16'he49;
        src71 <= 16'ha537;
        src72 <= 16'h37e1;
        src73 <= 16'hf272;
        src74 <= 16'h396d;
        src75 <= 16'h4106;
        src76 <= 16'hbd2e;
        src77 <= 16'h74e9;
        src78 <= 16'hd778;
        src79 <= 16'hfa9d;
        src80 <= 16'h4317;
        src81 <= 16'h394;
        src82 <= 16'hd8ac;
        src83 <= 16'h4ba3;
        src84 <= 16'h3953;
        src85 <= 16'h2408;
        src86 <= 16'h1be1;
        src87 <= 16'h2729;
        src88 <= 16'h5506;
        src89 <= 16'h2b83;
        src90 <= 16'h59af;
        src91 <= 16'ha89f;
        src92 <= 16'he012;
        src93 <= 16'hda45;
        src94 <= 16'h1480;
        src95 <= 16'h6f1d;
        src96 <= 16'h4d23;
        src97 <= 16'h5f5a;
        src98 <= 16'h6769;
        src99 <= 16'hc80b;
        src100 <= 16'hc10e;
        src101 <= 16'h3cd7;
        src102 <= 16'h49ef;
        src103 <= 16'hb0c8;
        src104 <= 16'h85ff;
        src105 <= 16'h7908;
        src106 <= 16'h972e;
        src107 <= 16'h6dcc;
        src108 <= 16'ha7ba;
        src109 <= 16'hfd17;
        src110 <= 16'hc7ec;
        src111 <= 16'he0be;
        src112 <= 16'h35c7;
        src113 <= 16'hce3d;
        src114 <= 16'h619f;
        src115 <= 16'hc8be;
        src116 <= 16'h9e0a;
        src117 <= 16'h5a9;
        src118 <= 16'h2c39;
        src119 <= 16'h38b4;
        src120 <= 16'h8b4a;
        src121 <= 16'h4db4;
        src122 <= 16'h5e37;
        src123 <= 16'h96ad;
        src124 <= 16'h66cc;
        src125 <= 16'h11d9;
        src126 <= 16'h1588;
        src127 <= 16'hb431;
        src128 <= 16'h626;
        src129 <= 16'heaf8;
        src130 <= 16'hdcf8;
        src131 <= 16'hf8fe;
        src132 <= 16'h2214;
        src133 <= 16'h981b;
        src134 <= 16'h904f;
        src135 <= 16'h8de6;
        src136 <= 16'h769a;
        src137 <= 16'hdab0;
        src138 <= 16'h1602;
        src139 <= 16'ha7d5;
        src140 <= 16'ha108;
        src141 <= 16'h2d49;
        src142 <= 16'h4df0;
        src143 <= 16'hf10c;
        src144 <= 16'hc640;
        src145 <= 16'h932e;
        src146 <= 16'h268d;
        src147 <= 16'h11ea;
        src148 <= 16'h9fcd;
        src149 <= 16'h2131;
        src150 <= 16'hf7e0;
        src151 <= 16'hdf9e;
        src152 <= 16'h4ac3;
        src153 <= 16'ha73f;
        src154 <= 16'hcd95;
        src155 <= 16'hd50e;
        src156 <= 16'hc3e4;
        src157 <= 16'h84e6;
        src158 <= 16'h488d;
        src159 <= 16'h676;
        src160 <= 16'h1ae1;
        src161 <= 16'hb872;
        exp <= 24'h511a0c;
        #1
        src0 <= 16'hc003;
        src1 <= 16'h39b6;
        src2 <= 16'h6c96;
        src3 <= 16'hcf80;
        src4 <= 16'ha84e;
        src5 <= 16'he08f;
        src6 <= 16'h4552;
        src7 <= 16'he3c4;
        src8 <= 16'hb072;
        src9 <= 16'hc3f4;
        src10 <= 16'h8327;
        src11 <= 16'h3f45;
        src12 <= 16'h90ab;
        src13 <= 16'heb3c;
        src14 <= 16'h97c;
        src15 <= 16'hcfb1;
        src16 <= 16'h22cd;
        src17 <= 16'hec3e;
        src18 <= 16'h9149;
        src19 <= 16'h2915;
        src20 <= 16'hd87;
        src21 <= 16'he74c;
        src22 <= 16'h26db;
        src23 <= 16'he355;
        src24 <= 16'h792f;
        src25 <= 16'hcdcf;
        src26 <= 16'hfb3;
        src27 <= 16'h5c1;
        src28 <= 16'h84c5;
        src29 <= 16'h684d;
        src30 <= 16'h4ba7;
        src31 <= 16'hfe3d;
        src32 <= 16'h6b2a;
        src33 <= 16'h9da7;
        src34 <= 16'h563a;
        src35 <= 16'h677f;
        src36 <= 16'h722f;
        src37 <= 16'hc236;
        src38 <= 16'h5cb3;
        src39 <= 16'hc511;
        src40 <= 16'hef28;
        src41 <= 16'hb6e;
        src42 <= 16'hc102;
        src43 <= 16'hbedb;
        src44 <= 16'hb8d8;
        src45 <= 16'h7070;
        src46 <= 16'h14fd;
        src47 <= 16'h931d;
        src48 <= 16'hcfcd;
        src49 <= 16'h51e8;
        src50 <= 16'h6e74;
        src51 <= 16'h487e;
        src52 <= 16'h4133;
        src53 <= 16'h8938;
        src54 <= 16'hc8db;
        src55 <= 16'h89d4;
        src56 <= 16'h93a9;
        src57 <= 16'hd78;
        src58 <= 16'h3a15;
        src59 <= 16'hb2b5;
        src60 <= 16'h9f7c;
        src61 <= 16'hbded;
        src62 <= 16'h1405;
        src63 <= 16'hfaa7;
        src64 <= 16'he7aa;
        src65 <= 16'had56;
        src66 <= 16'hbecd;
        src67 <= 16'h858d;
        src68 <= 16'h3214;
        src69 <= 16'ha910;
        src70 <= 16'h25de;
        src71 <= 16'hfada;
        src72 <= 16'he6a5;
        src73 <= 16'h4b77;
        src74 <= 16'ha7b7;
        src75 <= 16'h8ece;
        src76 <= 16'h26a5;
        src77 <= 16'h875e;
        src78 <= 16'he007;
        src79 <= 16'h71fc;
        src80 <= 16'hc9b5;
        src81 <= 16'hdee0;
        src82 <= 16'ha51a;
        src83 <= 16'h7fc9;
        src84 <= 16'h6c0f;
        src85 <= 16'he44b;
        src86 <= 16'h53b7;
        src87 <= 16'hb47d;
        src88 <= 16'h22a0;
        src89 <= 16'h5454;
        src90 <= 16'h3cd2;
        src91 <= 16'h918b;
        src92 <= 16'h6503;
        src93 <= 16'hea3;
        src94 <= 16'h30f;
        src95 <= 16'h2221;
        src96 <= 16'hcbe1;
        src97 <= 16'h9722;
        src98 <= 16'hf465;
        src99 <= 16'hbcc5;
        src100 <= 16'hc6d8;
        src101 <= 16'h6882;
        src102 <= 16'hfd81;
        src103 <= 16'h61fd;
        src104 <= 16'h3a2b;
        src105 <= 16'h5a29;
        src106 <= 16'h35b8;
        src107 <= 16'hf9d4;
        src108 <= 16'hc915;
        src109 <= 16'hb7c9;
        src110 <= 16'h3f8b;
        src111 <= 16'hf9d3;
        src112 <= 16'had72;
        src113 <= 16'h6a73;
        src114 <= 16'h24b5;
        src115 <= 16'h427c;
        src116 <= 16'hf8da;
        src117 <= 16'h671d;
        src118 <= 16'h958d;
        src119 <= 16'hdbfa;
        src120 <= 16'h90bf;
        src121 <= 16'he524;
        src122 <= 16'h8afe;
        src123 <= 16'h1a39;
        src124 <= 16'hc32f;
        src125 <= 16'hc0fc;
        src126 <= 16'h6beb;
        src127 <= 16'ha9b7;
        src128 <= 16'h8517;
        src129 <= 16'h18a1;
        src130 <= 16'hb3d7;
        src131 <= 16'h1128;
        src132 <= 16'h8b50;
        src133 <= 16'h9f7d;
        src134 <= 16'h1d98;
        src135 <= 16'h217d;
        src136 <= 16'h874;
        src137 <= 16'h5220;
        src138 <= 16'h412b;
        src139 <= 16'h7440;
        src140 <= 16'h9b8c;
        src141 <= 16'he27c;
        src142 <= 16'h5dfe;
        src143 <= 16'h5624;
        src144 <= 16'hb413;
        src145 <= 16'h185d;
        src146 <= 16'h1f68;
        src147 <= 16'h55f5;
        src148 <= 16'h9dae;
        src149 <= 16'h26bc;
        src150 <= 16'h2c26;
        src151 <= 16'h8198;
        src152 <= 16'h45ed;
        src153 <= 16'hb092;
        src154 <= 16'h4f11;
        src155 <= 16'h3793;
        src156 <= 16'heaf9;
        src157 <= 16'h5509;
        src158 <= 16'h55e3;
        src159 <= 16'h6579;
        src160 <= 16'h6be7;
        src161 <= 16'h3758;
        exp <= 24'h516ee2;
        #1
        src0 <= 16'h5e3e;
        src1 <= 16'h1414;
        src2 <= 16'h57ef;
        src3 <= 16'h8dbd;
        src4 <= 16'hd07c;
        src5 <= 16'h7abd;
        src6 <= 16'hbc09;
        src7 <= 16'h80d4;
        src8 <= 16'h87f7;
        src9 <= 16'hea78;
        src10 <= 16'h9ea8;
        src11 <= 16'h23c8;
        src12 <= 16'hf481;
        src13 <= 16'he9c2;
        src14 <= 16'hce3e;
        src15 <= 16'hc4fc;
        src16 <= 16'h351a;
        src17 <= 16'h7b7a;
        src18 <= 16'hca12;
        src19 <= 16'hd630;
        src20 <= 16'h4f7a;
        src21 <= 16'hefd9;
        src22 <= 16'hc686;
        src23 <= 16'h3692;
        src24 <= 16'h5164;
        src25 <= 16'hd568;
        src26 <= 16'h12e7;
        src27 <= 16'he553;
        src28 <= 16'h1f60;
        src29 <= 16'hf7d3;
        src30 <= 16'h9adc;
        src31 <= 16'h139a;
        src32 <= 16'h45f2;
        src33 <= 16'he5ea;
        src34 <= 16'hc747;
        src35 <= 16'h4744;
        src36 <= 16'hebbc;
        src37 <= 16'ha8c6;
        src38 <= 16'hcf16;
        src39 <= 16'h5c2a;
        src40 <= 16'h22f1;
        src41 <= 16'h7bad;
        src42 <= 16'h89e8;
        src43 <= 16'h275a;
        src44 <= 16'h3cf;
        src45 <= 16'h2f9;
        src46 <= 16'h4b4d;
        src47 <= 16'hbd0e;
        src48 <= 16'hb15e;
        src49 <= 16'h55eb;
        src50 <= 16'h1416;
        src51 <= 16'hbfb0;
        src52 <= 16'h65e7;
        src53 <= 16'h6733;
        src54 <= 16'hdf54;
        src55 <= 16'hc9b6;
        src56 <= 16'h9427;
        src57 <= 16'h50f8;
        src58 <= 16'h9356;
        src59 <= 16'h1d50;
        src60 <= 16'hc520;
        src61 <= 16'h4317;
        src62 <= 16'h891c;
        src63 <= 16'h734c;
        src64 <= 16'he08d;
        src65 <= 16'h7f3b;
        src66 <= 16'h6251;
        src67 <= 16'h1958;
        src68 <= 16'h2c7b;
        src69 <= 16'hffae;
        src70 <= 16'hd2f8;
        src71 <= 16'hb1e8;
        src72 <= 16'hbd0a;
        src73 <= 16'h74d5;
        src74 <= 16'hbe1f;
        src75 <= 16'h23be;
        src76 <= 16'hcae9;
        src77 <= 16'h4da4;
        src78 <= 16'h98b2;
        src79 <= 16'h80c7;
        src80 <= 16'hbbb1;
        src81 <= 16'h3179;
        src82 <= 16'h1957;
        src83 <= 16'h2991;
        src84 <= 16'hca2f;
        src85 <= 16'h8dd7;
        src86 <= 16'hee6c;
        src87 <= 16'h3709;
        src88 <= 16'h52bd;
        src89 <= 16'h759a;
        src90 <= 16'h6dba;
        src91 <= 16'ha123;
        src92 <= 16'h436;
        src93 <= 16'h2144;
        src94 <= 16'h1124;
        src95 <= 16'h64f;
        src96 <= 16'hcddd;
        src97 <= 16'hf98a;
        src98 <= 16'ha81b;
        src99 <= 16'h8d7;
        src100 <= 16'ha1f;
        src101 <= 16'h5f75;
        src102 <= 16'hd43d;
        src103 <= 16'hb455;
        src104 <= 16'h77ce;
        src105 <= 16'h8d67;
        src106 <= 16'he042;
        src107 <= 16'h9d3;
        src108 <= 16'h98a9;
        src109 <= 16'h5b77;
        src110 <= 16'hda4b;
        src111 <= 16'hde42;
        src112 <= 16'hbae8;
        src113 <= 16'hbf88;
        src114 <= 16'hd24a;
        src115 <= 16'h71be;
        src116 <= 16'h66c3;
        src117 <= 16'h5a96;
        src118 <= 16'h6660;
        src119 <= 16'hfc7;
        src120 <= 16'he3a0;
        src121 <= 16'h7686;
        src122 <= 16'h40ca;
        src123 <= 16'hb9b6;
        src124 <= 16'hca40;
        src125 <= 16'h8412;
        src126 <= 16'h1eca;
        src127 <= 16'hee8b;
        src128 <= 16'hff9b;
        src129 <= 16'h3847;
        src130 <= 16'h7061;
        src131 <= 16'h54d;
        src132 <= 16'hf6cb;
        src133 <= 16'hc396;
        src134 <= 16'h251a;
        src135 <= 16'h96e6;
        src136 <= 16'h4ee8;
        src137 <= 16'h3c07;
        src138 <= 16'h5585;
        src139 <= 16'h3251;
        src140 <= 16'h14c5;
        src141 <= 16'hf2b0;
        src142 <= 16'h8ddb;
        src143 <= 16'hb0b5;
        src144 <= 16'h1c06;
        src145 <= 16'hb95e;
        src146 <= 16'hea9;
        src147 <= 16'h74cc;
        src148 <= 16'hdb12;
        src149 <= 16'h178;
        src150 <= 16'hba1;
        src151 <= 16'h83ad;
        src152 <= 16'h85b6;
        src153 <= 16'h280;
        src154 <= 16'h7e43;
        src155 <= 16'h9205;
        src156 <= 16'h48e9;
        src157 <= 16'hd0c;
        src158 <= 16'h7981;
        src159 <= 16'h885d;
        src160 <= 16'h6fac;
        src161 <= 16'h149;
        exp <= 24'h4f207a;
        #1
        src0 <= 16'hd9e4;
        src1 <= 16'h4267;
        src2 <= 16'hc46f;
        src3 <= 16'hc5b1;
        src4 <= 16'h610c;
        src5 <= 16'h32b6;
        src6 <= 16'h13ec;
        src7 <= 16'h4e94;
        src8 <= 16'h488e;
        src9 <= 16'hb97d;
        src10 <= 16'hf4da;
        src11 <= 16'h3932;
        src12 <= 16'h6e4b;
        src13 <= 16'h5e37;
        src14 <= 16'h4d8c;
        src15 <= 16'hf613;
        src16 <= 16'hcc9a;
        src17 <= 16'h5521;
        src18 <= 16'hc316;
        src19 <= 16'h7d4e;
        src20 <= 16'hdd39;
        src21 <= 16'hf5c;
        src22 <= 16'hbfcd;
        src23 <= 16'hbd58;
        src24 <= 16'hd84f;
        src25 <= 16'hb423;
        src26 <= 16'h9d0f;
        src27 <= 16'h3993;
        src28 <= 16'he638;
        src29 <= 16'hcb19;
        src30 <= 16'h4a4;
        src31 <= 16'hb15c;
        src32 <= 16'hac72;
        src33 <= 16'h853;
        src34 <= 16'h4e07;
        src35 <= 16'hd857;
        src36 <= 16'hbc67;
        src37 <= 16'hc339;
        src38 <= 16'h6e14;
        src39 <= 16'h8394;
        src40 <= 16'h9cd1;
        src41 <= 16'h4b9d;
        src42 <= 16'h79c1;
        src43 <= 16'hc6ed;
        src44 <= 16'h5888;
        src45 <= 16'hb519;
        src46 <= 16'hff8;
        src47 <= 16'hc745;
        src48 <= 16'h3af5;
        src49 <= 16'h3ab3;
        src50 <= 16'heb48;
        src51 <= 16'habc4;
        src52 <= 16'h21f0;
        src53 <= 16'hcc34;
        src54 <= 16'h103f;
        src55 <= 16'h1de5;
        src56 <= 16'h845d;
        src57 <= 16'he093;
        src58 <= 16'hb22a;
        src59 <= 16'h20d1;
        src60 <= 16'h6ca2;
        src61 <= 16'hd05e;
        src62 <= 16'h663c;
        src63 <= 16'h822a;
        src64 <= 16'h4f2;
        src65 <= 16'h8088;
        src66 <= 16'h9328;
        src67 <= 16'h2f69;
        src68 <= 16'h5ebb;
        src69 <= 16'h7802;
        src70 <= 16'h1fbe;
        src71 <= 16'hfa9e;
        src72 <= 16'h9f94;
        src73 <= 16'h4eb6;
        src74 <= 16'heb5b;
        src75 <= 16'hc4bc;
        src76 <= 16'h927a;
        src77 <= 16'hf915;
        src78 <= 16'h2432;
        src79 <= 16'h5170;
        src80 <= 16'h4f0e;
        src81 <= 16'he443;
        src82 <= 16'h72a0;
        src83 <= 16'h1c12;
        src84 <= 16'hc70d;
        src85 <= 16'h16a8;
        src86 <= 16'h9bc9;
        src87 <= 16'h339a;
        src88 <= 16'h646c;
        src89 <= 16'hb675;
        src90 <= 16'h4e7b;
        src91 <= 16'h1ccb;
        src92 <= 16'h7029;
        src93 <= 16'hc836;
        src94 <= 16'h9b08;
        src95 <= 16'h82e2;
        src96 <= 16'hb4ef;
        src97 <= 16'h6e96;
        src98 <= 16'h4bc6;
        src99 <= 16'h6522;
        src100 <= 16'hff07;
        src101 <= 16'h91d8;
        src102 <= 16'hfd99;
        src103 <= 16'h34ac;
        src104 <= 16'h2d9f;
        src105 <= 16'h88;
        src106 <= 16'haea6;
        src107 <= 16'h5b56;
        src108 <= 16'hd918;
        src109 <= 16'h1d30;
        src110 <= 16'h48c2;
        src111 <= 16'hbf2c;
        src112 <= 16'h7276;
        src113 <= 16'h1d70;
        src114 <= 16'hbb06;
        src115 <= 16'hc381;
        src116 <= 16'h2f53;
        src117 <= 16'h366d;
        src118 <= 16'hb320;
        src119 <= 16'h19f;
        src120 <= 16'hc5ef;
        src121 <= 16'haf3e;
        src122 <= 16'h21db;
        src123 <= 16'h71a7;
        src124 <= 16'h12b6;
        src125 <= 16'h897a;
        src126 <= 16'h4d89;
        src127 <= 16'h99df;
        src128 <= 16'h2b20;
        src129 <= 16'hfe1a;
        src130 <= 16'h7fa9;
        src131 <= 16'he40b;
        src132 <= 16'h9a52;
        src133 <= 16'h3ba1;
        src134 <= 16'haa07;
        src135 <= 16'ha135;
        src136 <= 16'hd0ea;
        src137 <= 16'hcc80;
        src138 <= 16'ha6ac;
        src139 <= 16'h257;
        src140 <= 16'hf234;
        src141 <= 16'hccbd;
        src142 <= 16'hb433;
        src143 <= 16'h5065;
        src144 <= 16'hb189;
        src145 <= 16'h2d4b;
        src146 <= 16'he4c6;
        src147 <= 16'hf75a;
        src148 <= 16'h3489;
        src149 <= 16'hd4ff;
        src150 <= 16'ha983;
        src151 <= 16'h7c8b;
        src152 <= 16'h345f;
        src153 <= 16'h8fab;
        src154 <= 16'h2f66;
        src155 <= 16'hb1f8;
        src156 <= 16'hc1f7;
        src157 <= 16'hb928;
        src158 <= 16'h43fb;
        src159 <= 16'haeea;
        src160 <= 16'h9c1;
        src161 <= 16'h1a49;
        exp <= 24'h51d546;
        #1
        src0 <= 16'h2b39;
        src1 <= 16'h2be;
        src2 <= 16'hb3e1;
        src3 <= 16'h699d;
        src4 <= 16'h765b;
        src5 <= 16'h8c71;
        src6 <= 16'h8ff8;
        src7 <= 16'h6f80;
        src8 <= 16'h9a4d;
        src9 <= 16'h351c;
        src10 <= 16'ha215;
        src11 <= 16'h850f;
        src12 <= 16'h5724;
        src13 <= 16'h693e;
        src14 <= 16'h48da;
        src15 <= 16'h4f96;
        src16 <= 16'h9c24;
        src17 <= 16'h1baa;
        src18 <= 16'h6b09;
        src19 <= 16'h1a4f;
        src20 <= 16'hd0c;
        src21 <= 16'hf0dc;
        src22 <= 16'ha140;
        src23 <= 16'ha0f;
        src24 <= 16'h4ade;
        src25 <= 16'h60a5;
        src26 <= 16'h593;
        src27 <= 16'hf303;
        src28 <= 16'he56e;
        src29 <= 16'h695;
        src30 <= 16'h3884;
        src31 <= 16'hcfa8;
        src32 <= 16'h67b0;
        src33 <= 16'h98fb;
        src34 <= 16'he4e0;
        src35 <= 16'ha685;
        src36 <= 16'h77e4;
        src37 <= 16'hddbf;
        src38 <= 16'h6200;
        src39 <= 16'h1e9f;
        src40 <= 16'h23de;
        src41 <= 16'h3d8b;
        src42 <= 16'h8fd2;
        src43 <= 16'h1d33;
        src44 <= 16'hfe9d;
        src45 <= 16'h68a7;
        src46 <= 16'h4648;
        src47 <= 16'h9022;
        src48 <= 16'h61a1;
        src49 <= 16'h6c36;
        src50 <= 16'hbef9;
        src51 <= 16'heac5;
        src52 <= 16'h5464;
        src53 <= 16'h9198;
        src54 <= 16'h99d;
        src55 <= 16'h26df;
        src56 <= 16'h70ff;
        src57 <= 16'h4df2;
        src58 <= 16'hd71e;
        src59 <= 16'ha677;
        src60 <= 16'he832;
        src61 <= 16'hb16b;
        src62 <= 16'h6e6a;
        src63 <= 16'h945;
        src64 <= 16'h481e;
        src65 <= 16'hedad;
        src66 <= 16'hde31;
        src67 <= 16'hb45b;
        src68 <= 16'h76d;
        src69 <= 16'he533;
        src70 <= 16'he654;
        src71 <= 16'h59e9;
        src72 <= 16'h148d;
        src73 <= 16'hedf5;
        src74 <= 16'he161;
        src75 <= 16'he612;
        src76 <= 16'heb9b;
        src77 <= 16'hf99f;
        src78 <= 16'hd7fe;
        src79 <= 16'h9d5c;
        src80 <= 16'hc9e7;
        src81 <= 16'hc664;
        src82 <= 16'hade1;
        src83 <= 16'h9754;
        src84 <= 16'h7c1;
        src85 <= 16'h81c1;
        src86 <= 16'had9b;
        src87 <= 16'hbb97;
        src88 <= 16'hf1bc;
        src89 <= 16'h94e2;
        src90 <= 16'h4d0a;
        src91 <= 16'h5c24;
        src92 <= 16'h39f4;
        src93 <= 16'hd44e;
        src94 <= 16'h36ab;
        src95 <= 16'he953;
        src96 <= 16'h8fca;
        src97 <= 16'hf488;
        src98 <= 16'h2fe9;
        src99 <= 16'h711c;
        src100 <= 16'h77ba;
        src101 <= 16'hd16b;
        src102 <= 16'h93e1;
        src103 <= 16'ha7ca;
        src104 <= 16'ha111;
        src105 <= 16'h964d;
        src106 <= 16'h4b0b;
        src107 <= 16'h4736;
        src108 <= 16'ha482;
        src109 <= 16'hbfd8;
        src110 <= 16'h8e3;
        src111 <= 16'h8320;
        src112 <= 16'h3f4;
        src113 <= 16'h8758;
        src114 <= 16'hea1d;
        src115 <= 16'h2f20;
        src116 <= 16'h5c65;
        src117 <= 16'hfaae;
        src118 <= 16'h8523;
        src119 <= 16'h57f;
        src120 <= 16'hb9d3;
        src121 <= 16'h79a7;
        src122 <= 16'h428c;
        src123 <= 16'hec31;
        src124 <= 16'h7ca3;
        src125 <= 16'h50fa;
        src126 <= 16'h3320;
        src127 <= 16'hb94f;
        src128 <= 16'h99c9;
        src129 <= 16'h74a3;
        src130 <= 16'h137;
        src131 <= 16'h1074;
        src132 <= 16'h6d6b;
        src133 <= 16'hefe0;
        src134 <= 16'hdf7b;
        src135 <= 16'h6276;
        src136 <= 16'h996a;
        src137 <= 16'h798a;
        src138 <= 16'h321f;
        src139 <= 16'hb559;
        src140 <= 16'h4f7a;
        src141 <= 16'h3f77;
        src142 <= 16'he93e;
        src143 <= 16'ha31d;
        src144 <= 16'haaa3;
        src145 <= 16'h706e;
        src146 <= 16'h26ed;
        src147 <= 16'hfc92;
        src148 <= 16'h51ea;
        src149 <= 16'hf51d;
        src150 <= 16'hddfe;
        src151 <= 16'h8096;
        src152 <= 16'h390a;
        src153 <= 16'hb86e;
        src154 <= 16'h1964;
        src155 <= 16'h5004;
        src156 <= 16'h88f5;
        src157 <= 16'h294c;
        src158 <= 16'h4fb4;
        src159 <= 16'h6646;
        src160 <= 16'ha91d;
        src161 <= 16'hb4b6;
        exp <= 24'h51c6cf;
        #1
        src0 <= 16'he1a2;
        src1 <= 16'h89bf;
        src2 <= 16'hedb5;
        src3 <= 16'h528b;
        src4 <= 16'hf7b4;
        src5 <= 16'h6e0a;
        src6 <= 16'h31ec;
        src7 <= 16'h4af;
        src8 <= 16'h9584;
        src9 <= 16'h610c;
        src10 <= 16'h98d7;
        src11 <= 16'hcdc0;
        src12 <= 16'h561e;
        src13 <= 16'h5c5a;
        src14 <= 16'heb52;
        src15 <= 16'h85af;
        src16 <= 16'he538;
        src17 <= 16'he93b;
        src18 <= 16'h4b44;
        src19 <= 16'ha0f1;
        src20 <= 16'h87f2;
        src21 <= 16'hec65;
        src22 <= 16'h967f;
        src23 <= 16'h90aa;
        src24 <= 16'h583c;
        src25 <= 16'h3ff3;
        src26 <= 16'hf30a;
        src27 <= 16'h5628;
        src28 <= 16'hc3a9;
        src29 <= 16'h9352;
        src30 <= 16'ha4b5;
        src31 <= 16'h2157;
        src32 <= 16'hfba4;
        src33 <= 16'hfd0;
        src34 <= 16'hfbb0;
        src35 <= 16'heb1e;
        src36 <= 16'h9e9f;
        src37 <= 16'h43fe;
        src38 <= 16'heb62;
        src39 <= 16'h1ceb;
        src40 <= 16'hc2a8;
        src41 <= 16'h3be9;
        src42 <= 16'he24;
        src43 <= 16'hb437;
        src44 <= 16'h82a2;
        src45 <= 16'hd316;
        src46 <= 16'h223c;
        src47 <= 16'h562f;
        src48 <= 16'hfae8;
        src49 <= 16'ha77d;
        src50 <= 16'h69ee;
        src51 <= 16'h6440;
        src52 <= 16'h60ad;
        src53 <= 16'h404d;
        src54 <= 16'hb2ee;
        src55 <= 16'h7350;
        src56 <= 16'hf3f4;
        src57 <= 16'hc58a;
        src58 <= 16'h79df;
        src59 <= 16'h6ae1;
        src60 <= 16'ha19e;
        src61 <= 16'h848;
        src62 <= 16'hde78;
        src63 <= 16'h2bde;
        src64 <= 16'h98d6;
        src65 <= 16'h5937;
        src66 <= 16'h1cd2;
        src67 <= 16'h43bf;
        src68 <= 16'he81a;
        src69 <= 16'hb7f6;
        src70 <= 16'hf267;
        src71 <= 16'h4451;
        src72 <= 16'h2b6e;
        src73 <= 16'h6416;
        src74 <= 16'h85ea;
        src75 <= 16'hdd37;
        src76 <= 16'hbc1a;
        src77 <= 16'h7e4f;
        src78 <= 16'h42f6;
        src79 <= 16'h6859;
        src80 <= 16'he58c;
        src81 <= 16'h7474;
        src82 <= 16'hee1e;
        src83 <= 16'hdcf6;
        src84 <= 16'h6b1f;
        src85 <= 16'h67ff;
        src86 <= 16'h2889;
        src87 <= 16'h10bb;
        src88 <= 16'h3739;
        src89 <= 16'hbab0;
        src90 <= 16'h364d;
        src91 <= 16'hdf76;
        src92 <= 16'hf955;
        src93 <= 16'hfb3d;
        src94 <= 16'h3f71;
        src95 <= 16'h9879;
        src96 <= 16'h2d20;
        src97 <= 16'h104f;
        src98 <= 16'h4084;
        src99 <= 16'he379;
        src100 <= 16'h34f6;
        src101 <= 16'habf8;
        src102 <= 16'h867f;
        src103 <= 16'ha631;
        src104 <= 16'h883c;
        src105 <= 16'hd778;
        src106 <= 16'h64a6;
        src107 <= 16'hb3c7;
        src108 <= 16'h82a0;
        src109 <= 16'ha7f4;
        src110 <= 16'h82c7;
        src111 <= 16'had03;
        src112 <= 16'haa41;
        src113 <= 16'hdbaa;
        src114 <= 16'h35d;
        src115 <= 16'h27ee;
        src116 <= 16'h7629;
        src117 <= 16'hd48e;
        src118 <= 16'h9076;
        src119 <= 16'he99b;
        src120 <= 16'hf1e0;
        src121 <= 16'he46d;
        src122 <= 16'h1c05;
        src123 <= 16'hc60c;
        src124 <= 16'hcf65;
        src125 <= 16'h4d4d;
        src126 <= 16'ha6bf;
        src127 <= 16'hb52c;
        src128 <= 16'he6d5;
        src129 <= 16'h35af;
        src130 <= 16'h7f5d;
        src131 <= 16'hf5bf;
        src132 <= 16'hd506;
        src133 <= 16'hd5ba;
        src134 <= 16'h1598;
        src135 <= 16'hcda3;
        src136 <= 16'hca9;
        src137 <= 16'h6cac;
        src138 <= 16'h8340;
        src139 <= 16'hf16d;
        src140 <= 16'hc936;
        src141 <= 16'hb484;
        src142 <= 16'hd567;
        src143 <= 16'h457e;
        src144 <= 16'haac3;
        src145 <= 16'h74db;
        src146 <= 16'haf4c;
        src147 <= 16'hb064;
        src148 <= 16'h4386;
        src149 <= 16'hc6e4;
        src150 <= 16'h82dd;
        src151 <= 16'hba96;
        src152 <= 16'hae79;
        src153 <= 16'h1c9e;
        src154 <= 16'h8717;
        src155 <= 16'h5a08;
        src156 <= 16'hdea2;
        src157 <= 16'he125;
        src158 <= 16'h854d;
        src159 <= 16'h56b8;
        src160 <= 16'h574c;
        src161 <= 16'hce92;
        exp <= 24'h59ded4;
        #1
        src0 <= 16'h77b;
        src1 <= 16'h6dbd;
        src2 <= 16'h7a7f;
        src3 <= 16'h8cdf;
        src4 <= 16'hafc7;
        src5 <= 16'h4c51;
        src6 <= 16'h6598;
        src7 <= 16'h1d86;
        src8 <= 16'h12d6;
        src9 <= 16'h3b66;
        src10 <= 16'haf0;
        src11 <= 16'h59bc;
        src12 <= 16'hb4b4;
        src13 <= 16'hd2aa;
        src14 <= 16'hd1df;
        src15 <= 16'h87a1;
        src16 <= 16'h539c;
        src17 <= 16'h5d5c;
        src18 <= 16'hfbfc;
        src19 <= 16'h4c1e;
        src20 <= 16'hda30;
        src21 <= 16'h1183;
        src22 <= 16'ha4e7;
        src23 <= 16'h81c;
        src24 <= 16'hacf5;
        src25 <= 16'h240d;
        src26 <= 16'hcf1c;
        src27 <= 16'h1eb5;
        src28 <= 16'h3fe2;
        src29 <= 16'hfe0e;
        src30 <= 16'h76c6;
        src31 <= 16'h25b3;
        src32 <= 16'h77b6;
        src33 <= 16'h585e;
        src34 <= 16'ha8ed;
        src35 <= 16'hf17a;
        src36 <= 16'he55e;
        src37 <= 16'h857f;
        src38 <= 16'h318f;
        src39 <= 16'hb45;
        src40 <= 16'h4c6;
        src41 <= 16'h71b7;
        src42 <= 16'h294b;
        src43 <= 16'h7987;
        src44 <= 16'h7b8d;
        src45 <= 16'hba52;
        src46 <= 16'h6e7a;
        src47 <= 16'hcb66;
        src48 <= 16'h2a66;
        src49 <= 16'h1ac8;
        src50 <= 16'hcb2d;
        src51 <= 16'h89c3;
        src52 <= 16'hcaf2;
        src53 <= 16'h4521;
        src54 <= 16'h7162;
        src55 <= 16'he336;
        src56 <= 16'h96a6;
        src57 <= 16'h942f;
        src58 <= 16'hd790;
        src59 <= 16'h49d8;
        src60 <= 16'h6453;
        src61 <= 16'h4eec;
        src62 <= 16'h7689;
        src63 <= 16'h8be;
        src64 <= 16'haad1;
        src65 <= 16'h71b5;
        src66 <= 16'h5037;
        src67 <= 16'hd845;
        src68 <= 16'hac07;
        src69 <= 16'hb9a7;
        src70 <= 16'hbe0a;
        src71 <= 16'hbc9a;
        src72 <= 16'h986a;
        src73 <= 16'hd817;
        src74 <= 16'h3f66;
        src75 <= 16'ha063;
        src76 <= 16'h157d;
        src77 <= 16'hf78b;
        src78 <= 16'h908d;
        src79 <= 16'h9eee;
        src80 <= 16'hb787;
        src81 <= 16'hc490;
        src82 <= 16'h2753;
        src83 <= 16'h1c03;
        src84 <= 16'h5f03;
        src85 <= 16'h5e8f;
        src86 <= 16'h333;
        src87 <= 16'h1167;
        src88 <= 16'h2fe4;
        src89 <= 16'h55bb;
        src90 <= 16'h7f32;
        src91 <= 16'hbd1c;
        src92 <= 16'h85e;
        src93 <= 16'h778e;
        src94 <= 16'hdc89;
        src95 <= 16'h4f2c;
        src96 <= 16'h21a;
        src97 <= 16'ha215;
        src98 <= 16'h6e60;
        src99 <= 16'h34b6;
        src100 <= 16'h8ef0;
        src101 <= 16'hfe33;
        src102 <= 16'hf64;
        src103 <= 16'h9b72;
        src104 <= 16'h7ffe;
        src105 <= 16'hb7cc;
        src106 <= 16'h83b4;
        src107 <= 16'h1c15;
        src108 <= 16'h70ff;
        src109 <= 16'h2fab;
        src110 <= 16'hc89;
        src111 <= 16'hf4df;
        src112 <= 16'h3288;
        src113 <= 16'hba91;
        src114 <= 16'h5a46;
        src115 <= 16'h54f7;
        src116 <= 16'hb7f6;
        src117 <= 16'he2cb;
        src118 <= 16'hd3fb;
        src119 <= 16'h4c2b;
        src120 <= 16'h8c04;
        src121 <= 16'h84f4;
        src122 <= 16'ha1e8;
        src123 <= 16'h54dd;
        src124 <= 16'hd817;
        src125 <= 16'hd734;
        src126 <= 16'h6788;
        src127 <= 16'h610d;
        src128 <= 16'hcc6;
        src129 <= 16'h750e;
        src130 <= 16'hbf6;
        src131 <= 16'h6f59;
        src132 <= 16'h48b0;
        src133 <= 16'hba41;
        src134 <= 16'h8799;
        src135 <= 16'h98f9;
        src136 <= 16'h4012;
        src137 <= 16'h924f;
        src138 <= 16'hd603;
        src139 <= 16'heb65;
        src140 <= 16'hc88f;
        src141 <= 16'h1013;
        src142 <= 16'h4828;
        src143 <= 16'h37f;
        src144 <= 16'hf23c;
        src145 <= 16'h9499;
        src146 <= 16'h4f4f;
        src147 <= 16'h1340;
        src148 <= 16'ha1a2;
        src149 <= 16'heb5a;
        src150 <= 16'h8183;
        src151 <= 16'hb2d8;
        src152 <= 16'h1c56;
        src153 <= 16'h60d7;
        src154 <= 16'h57ff;
        src155 <= 16'he377;
        src156 <= 16'h8cc6;
        src157 <= 16'h6c9f;
        src158 <= 16'h51ab;
        src159 <= 16'hfd8e;
        src160 <= 16'hd466;
        src161 <= 16'hf204;
        exp <= 24'h4d9f7f;
        #1
        src0 <= 16'hf34;
        src1 <= 16'h8df4;
        src2 <= 16'h583e;
        src3 <= 16'ha165;
        src4 <= 16'hd4c9;
        src5 <= 16'h7a84;
        src6 <= 16'h30e2;
        src7 <= 16'hbbb;
        src8 <= 16'hc695;
        src9 <= 16'h359b;
        src10 <= 16'hd952;
        src11 <= 16'hc91d;
        src12 <= 16'hd922;
        src13 <= 16'hec04;
        src14 <= 16'hca36;
        src15 <= 16'h3a61;
        src16 <= 16'hae73;
        src17 <= 16'h669f;
        src18 <= 16'h70ce;
        src19 <= 16'h8871;
        src20 <= 16'h33e7;
        src21 <= 16'hb414;
        src22 <= 16'h920d;
        src23 <= 16'h7fcd;
        src24 <= 16'h6a2f;
        src25 <= 16'hbf8b;
        src26 <= 16'h3be4;
        src27 <= 16'hddfb;
        src28 <= 16'haf45;
        src29 <= 16'hd8f;
        src30 <= 16'h6354;
        src31 <= 16'haead;
        src32 <= 16'h7f60;
        src33 <= 16'h62d5;
        src34 <= 16'habb6;
        src35 <= 16'hc88f;
        src36 <= 16'h9449;
        src37 <= 16'hd7b9;
        src38 <= 16'h950f;
        src39 <= 16'h7689;
        src40 <= 16'h45c5;
        src41 <= 16'h500a;
        src42 <= 16'hdee8;
        src43 <= 16'he42;
        src44 <= 16'h6b8c;
        src45 <= 16'hc5fa;
        src46 <= 16'h4e0d;
        src47 <= 16'hd373;
        src48 <= 16'hc5d0;
        src49 <= 16'h30e6;
        src50 <= 16'hff2a;
        src51 <= 16'h679f;
        src52 <= 16'hb91f;
        src53 <= 16'h5c89;
        src54 <= 16'hb044;
        src55 <= 16'h38dd;
        src56 <= 16'h5d1b;
        src57 <= 16'h5e05;
        src58 <= 16'h2176;
        src59 <= 16'h6ae2;
        src60 <= 16'h2937;
        src61 <= 16'h77bd;
        src62 <= 16'h3b1;
        src63 <= 16'he9bf;
        src64 <= 16'h2045;
        src65 <= 16'h2f5b;
        src66 <= 16'h36ac;
        src67 <= 16'h430e;
        src68 <= 16'h415c;
        src69 <= 16'h6b66;
        src70 <= 16'he6a4;
        src71 <= 16'he5e0;
        src72 <= 16'h8c57;
        src73 <= 16'h93df;
        src74 <= 16'h5a19;
        src75 <= 16'h8a47;
        src76 <= 16'h6ed6;
        src77 <= 16'hfe29;
        src78 <= 16'h8822;
        src79 <= 16'h74aa;
        src80 <= 16'h7871;
        src81 <= 16'h11da;
        src82 <= 16'hd709;
        src83 <= 16'h5189;
        src84 <= 16'h18cd;
        src85 <= 16'h8832;
        src86 <= 16'haa5f;
        src87 <= 16'he68;
        src88 <= 16'h76b6;
        src89 <= 16'hd8af;
        src90 <= 16'hd2a9;
        src91 <= 16'h1eb1;
        src92 <= 16'h927f;
        src93 <= 16'hb4ab;
        src94 <= 16'h4c51;
        src95 <= 16'h69da;
        src96 <= 16'h7aa9;
        src97 <= 16'hcc59;
        src98 <= 16'he182;
        src99 <= 16'hf86e;
        src100 <= 16'h4b78;
        src101 <= 16'h10c2;
        src102 <= 16'ha663;
        src103 <= 16'h4ee3;
        src104 <= 16'h124c;
        src105 <= 16'h779d;
        src106 <= 16'h2eac;
        src107 <= 16'hfa9e;
        src108 <= 16'hbd0d;
        src109 <= 16'h41ad;
        src110 <= 16'hd15f;
        src111 <= 16'h9f7d;
        src112 <= 16'h85fe;
        src113 <= 16'h539c;
        src114 <= 16'h3dfe;
        src115 <= 16'ha0f9;
        src116 <= 16'h984f;
        src117 <= 16'h2633;
        src118 <= 16'h43d2;
        src119 <= 16'h24ce;
        src120 <= 16'hd4e9;
        src121 <= 16'h7bec;
        src122 <= 16'he9bc;
        src123 <= 16'h6758;
        src124 <= 16'h8c59;
        src125 <= 16'h2c2c;
        src126 <= 16'hd000;
        src127 <= 16'h35d5;
        src128 <= 16'h8901;
        src129 <= 16'hbe90;
        src130 <= 16'h5b8e;
        src131 <= 16'hde7a;
        src132 <= 16'hf3c4;
        src133 <= 16'h9eb8;
        src134 <= 16'h5dbc;
        src135 <= 16'hf586;
        src136 <= 16'h77ba;
        src137 <= 16'h3487;
        src138 <= 16'hfdaa;
        src139 <= 16'h1382;
        src140 <= 16'hd491;
        src141 <= 16'hac2;
        src142 <= 16'h87a3;
        src143 <= 16'h8801;
        src144 <= 16'hb0fb;
        src145 <= 16'h2461;
        src146 <= 16'h963a;
        src147 <= 16'h18f6;
        src148 <= 16'hea9f;
        src149 <= 16'h72f3;
        src150 <= 16'h488b;
        src151 <= 16'heb17;
        src152 <= 16'h879a;
        src153 <= 16'hf76a;
        src154 <= 16'hd96d;
        src155 <= 16'hf62e;
        src156 <= 16'h19cc;
        src157 <= 16'hfba2;
        src158 <= 16'hc9ae;
        src159 <= 16'hc08;
        src160 <= 16'hb847;
        src161 <= 16'h9ff8;
        exp <= 24'h530842;
        #1
        src0 <= 16'h7dad;
        src1 <= 16'h1add;
        src2 <= 16'h26cb;
        src3 <= 16'hf161;
        src4 <= 16'hc4ab;
        src5 <= 16'h92f;
        src6 <= 16'h8a04;
        src7 <= 16'h18e8;
        src8 <= 16'h3987;
        src9 <= 16'hdb2e;
        src10 <= 16'h3338;
        src11 <= 16'h1680;
        src12 <= 16'h1d3b;
        src13 <= 16'h5e99;
        src14 <= 16'h84c6;
        src15 <= 16'he3d7;
        src16 <= 16'hd161;
        src17 <= 16'h95b;
        src18 <= 16'h766b;
        src19 <= 16'hb95;
        src20 <= 16'h3deb;
        src21 <= 16'hb349;
        src22 <= 16'h86d0;
        src23 <= 16'h3283;
        src24 <= 16'h64a4;
        src25 <= 16'h139b;
        src26 <= 16'h6e34;
        src27 <= 16'h1eee;
        src28 <= 16'hb72a;
        src29 <= 16'hf109;
        src30 <= 16'hbfb0;
        src31 <= 16'he9cf;
        src32 <= 16'h12cb;
        src33 <= 16'h9593;
        src34 <= 16'h6a6c;
        src35 <= 16'h3d1;
        src36 <= 16'h908b;
        src37 <= 16'h6d87;
        src38 <= 16'h8529;
        src39 <= 16'h40b2;
        src40 <= 16'h6bb0;
        src41 <= 16'hf5ea;
        src42 <= 16'h46fd;
        src43 <= 16'h6a27;
        src44 <= 16'h1aa1;
        src45 <= 16'hc58a;
        src46 <= 16'he5bc;
        src47 <= 16'hcd86;
        src48 <= 16'hb393;
        src49 <= 16'h1f21;
        src50 <= 16'h7cbd;
        src51 <= 16'hde5b;
        src52 <= 16'h81ac;
        src53 <= 16'h9e93;
        src54 <= 16'ha9cb;
        src55 <= 16'hfd21;
        src56 <= 16'h3e87;
        src57 <= 16'hb0a5;
        src58 <= 16'h2fd0;
        src59 <= 16'hc91;
        src60 <= 16'he629;
        src61 <= 16'ha6aa;
        src62 <= 16'h1373;
        src63 <= 16'hf230;
        src64 <= 16'h23eb;
        src65 <= 16'h8306;
        src66 <= 16'h288;
        src67 <= 16'h62b0;
        src68 <= 16'h4198;
        src69 <= 16'hc83c;
        src70 <= 16'h5d6f;
        src71 <= 16'h3da6;
        src72 <= 16'hbae9;
        src73 <= 16'h948;
        src74 <= 16'hf411;
        src75 <= 16'h2708;
        src76 <= 16'h9f2c;
        src77 <= 16'hb426;
        src78 <= 16'ha527;
        src79 <= 16'h3023;
        src80 <= 16'h1de7;
        src81 <= 16'h7a31;
        src82 <= 16'h27ce;
        src83 <= 16'hb60f;
        src84 <= 16'ha323;
        src85 <= 16'hbf3c;
        src86 <= 16'h2a12;
        src87 <= 16'ha0e0;
        src88 <= 16'h7cfb;
        src89 <= 16'h7851;
        src90 <= 16'h24ed;
        src91 <= 16'hb20;
        src92 <= 16'hdfd;
        src93 <= 16'h8adf;
        src94 <= 16'h4367;
        src95 <= 16'ha1d;
        src96 <= 16'h8b2;
        src97 <= 16'h237f;
        src98 <= 16'h1824;
        src99 <= 16'h64ad;
        src100 <= 16'hadce;
        src101 <= 16'h56ab;
        src102 <= 16'h112b;
        src103 <= 16'hd17b;
        src104 <= 16'h6ce5;
        src105 <= 16'h66c0;
        src106 <= 16'h7e8f;
        src107 <= 16'hbe2d;
        src108 <= 16'h3d86;
        src109 <= 16'h2ded;
        src110 <= 16'hac44;
        src111 <= 16'h7b7e;
        src112 <= 16'ha7b5;
        src113 <= 16'h1b5f;
        src114 <= 16'h4e45;
        src115 <= 16'h3469;
        src116 <= 16'h443a;
        src117 <= 16'h1ae2;
        src118 <= 16'h66d6;
        src119 <= 16'h9256;
        src120 <= 16'ha65b;
        src121 <= 16'hf6d1;
        src122 <= 16'hb7db;
        src123 <= 16'h8fd1;
        src124 <= 16'h4704;
        src125 <= 16'h2c3a;
        src126 <= 16'h356d;
        src127 <= 16'h2c70;
        src128 <= 16'hda85;
        src129 <= 16'hb30f;
        src130 <= 16'h9327;
        src131 <= 16'h59e;
        src132 <= 16'hcb8a;
        src133 <= 16'h6f76;
        src134 <= 16'hcb5c;
        src135 <= 16'hfee5;
        src136 <= 16'h4db2;
        src137 <= 16'h7503;
        src138 <= 16'h38d3;
        src139 <= 16'h8ab;
        src140 <= 16'hce76;
        src141 <= 16'hde00;
        src142 <= 16'hb71d;
        src143 <= 16'hb4a7;
        src144 <= 16'hb5f0;
        src145 <= 16'hc9fa;
        src146 <= 16'h7fa0;
        src147 <= 16'h4500;
        src148 <= 16'he81e;
        src149 <= 16'h6e69;
        src150 <= 16'hb252;
        src151 <= 16'h7c4d;
        src152 <= 16'h809a;
        src153 <= 16'hc38f;
        src154 <= 16'h109c;
        src155 <= 16'h971f;
        src156 <= 16'hce8c;
        src157 <= 16'h2961;
        src158 <= 16'h791a;
        src159 <= 16'hf426;
        src160 <= 16'he01d;
        src161 <= 16'hffdd;
        exp <= 24'h4b2cca;
        #1
        src0 <= 16'h97f;
        src1 <= 16'h8c65;
        src2 <= 16'hb1c7;
        src3 <= 16'he97a;
        src4 <= 16'h735f;
        src5 <= 16'he709;
        src6 <= 16'hfa62;
        src7 <= 16'h92fd;
        src8 <= 16'h9054;
        src9 <= 16'h172a;
        src10 <= 16'hd9e5;
        src11 <= 16'h9348;
        src12 <= 16'h4040;
        src13 <= 16'h3735;
        src14 <= 16'haac3;
        src15 <= 16'h9aef;
        src16 <= 16'h29e3;
        src17 <= 16'h3a2b;
        src18 <= 16'he0e8;
        src19 <= 16'h1602;
        src20 <= 16'ha0b4;
        src21 <= 16'h790e;
        src22 <= 16'hf7df;
        src23 <= 16'h8ade;
        src24 <= 16'he9b8;
        src25 <= 16'hdd33;
        src26 <= 16'hc13c;
        src27 <= 16'h569;
        src28 <= 16'he520;
        src29 <= 16'hdc17;
        src30 <= 16'h3c3d;
        src31 <= 16'hd71d;
        src32 <= 16'hd6ed;
        src33 <= 16'h4d46;
        src34 <= 16'h4b2a;
        src35 <= 16'h7ca7;
        src36 <= 16'h8f54;
        src37 <= 16'h8abe;
        src38 <= 16'h94ab;
        src39 <= 16'h6541;
        src40 <= 16'hd17b;
        src41 <= 16'h6b09;
        src42 <= 16'hefe8;
        src43 <= 16'h6076;
        src44 <= 16'hc246;
        src45 <= 16'h71d3;
        src46 <= 16'h53d4;
        src47 <= 16'h66;
        src48 <= 16'hbc41;
        src49 <= 16'ha3f0;
        src50 <= 16'h4258;
        src51 <= 16'h47e;
        src52 <= 16'h46e6;
        src53 <= 16'h962;
        src54 <= 16'h9587;
        src55 <= 16'h8104;
        src56 <= 16'hf558;
        src57 <= 16'hac5f;
        src58 <= 16'h1840;
        src59 <= 16'h2974;
        src60 <= 16'hd148;
        src61 <= 16'h1434;
        src62 <= 16'h2fb0;
        src63 <= 16'h9208;
        src64 <= 16'h553d;
        src65 <= 16'hdfb;
        src66 <= 16'hd436;
        src67 <= 16'hb03e;
        src68 <= 16'h7a9e;
        src69 <= 16'h2568;
        src70 <= 16'hb5d4;
        src71 <= 16'h539a;
        src72 <= 16'h4115;
        src73 <= 16'h6031;
        src74 <= 16'h2c6e;
        src75 <= 16'h4cfe;
        src76 <= 16'hf13c;
        src77 <= 16'h4e02;
        src78 <= 16'heed8;
        src79 <= 16'h7b82;
        src80 <= 16'h6b74;
        src81 <= 16'h775a;
        src82 <= 16'hf4fd;
        src83 <= 16'h94aa;
        src84 <= 16'hf57a;
        src85 <= 16'hcdcb;
        src86 <= 16'hbaf0;
        src87 <= 16'hbf5f;
        src88 <= 16'h3937;
        src89 <= 16'h7e26;
        src90 <= 16'hbc37;
        src91 <= 16'h9686;
        src92 <= 16'hac91;
        src93 <= 16'h89cd;
        src94 <= 16'h6e86;
        src95 <= 16'he6d0;
        src96 <= 16'h8b63;
        src97 <= 16'h370c;
        src98 <= 16'hb8c4;
        src99 <= 16'ha8e2;
        src100 <= 16'hca4c;
        src101 <= 16'h2618;
        src102 <= 16'h28c0;
        src103 <= 16'h8f0a;
        src104 <= 16'h7be5;
        src105 <= 16'h35da;
        src106 <= 16'h6675;
        src107 <= 16'h2f7c;
        src108 <= 16'hf9d2;
        src109 <= 16'h5e89;
        src110 <= 16'h9a82;
        src111 <= 16'hdc68;
        src112 <= 16'h3088;
        src113 <= 16'hc5bf;
        src114 <= 16'hbc75;
        src115 <= 16'hd9ac;
        src116 <= 16'ha34b;
        src117 <= 16'h160b;
        src118 <= 16'ha65b;
        src119 <= 16'h1dc7;
        src120 <= 16'hbbb9;
        src121 <= 16'h723e;
        src122 <= 16'h628c;
        src123 <= 16'hcfba;
        src124 <= 16'hfc15;
        src125 <= 16'h7109;
        src126 <= 16'hcf3;
        src127 <= 16'hfe92;
        src128 <= 16'h330b;
        src129 <= 16'h3271;
        src130 <= 16'h973c;
        src131 <= 16'hc3f2;
        src132 <= 16'hf412;
        src133 <= 16'hc708;
        src134 <= 16'h7db1;
        src135 <= 16'h7908;
        src136 <= 16'h3bf0;
        src137 <= 16'h14ec;
        src138 <= 16'h36b0;
        src139 <= 16'h280c;
        src140 <= 16'h1834;
        src141 <= 16'h41eb;
        src142 <= 16'h288b;
        src143 <= 16'hccc7;
        src144 <= 16'hbe46;
        src145 <= 16'h3452;
        src146 <= 16'hb07b;
        src147 <= 16'hf360;
        src148 <= 16'haaaa;
        src149 <= 16'hb01c;
        src150 <= 16'hf5ff;
        src151 <= 16'hbe95;
        src152 <= 16'h83ef;
        src153 <= 16'h54b6;
        src154 <= 16'hb5c1;
        src155 <= 16'hedf5;
        src156 <= 16'he1b;
        src157 <= 16'hb3c;
        src158 <= 16'h3c63;
        src159 <= 16'h4dfa;
        src160 <= 16'h808f;
        src161 <= 16'hc826;
        exp <= 24'h53cd56;
        #1
        src0 <= 16'hb9d9;
        src1 <= 16'hc074;
        src2 <= 16'h88c3;
        src3 <= 16'h86c9;
        src4 <= 16'hff72;
        src5 <= 16'h2263;
        src6 <= 16'h3725;
        src7 <= 16'hdc0d;
        src8 <= 16'ha4e6;
        src9 <= 16'hb09d;
        src10 <= 16'he7f5;
        src11 <= 16'h68f6;
        src12 <= 16'h170b;
        src13 <= 16'hd6c7;
        src14 <= 16'hf97;
        src15 <= 16'h5180;
        src16 <= 16'h5d24;
        src17 <= 16'h6c0b;
        src18 <= 16'ha604;
        src19 <= 16'h7092;
        src20 <= 16'h2b35;
        src21 <= 16'h52c5;
        src22 <= 16'hb876;
        src23 <= 16'ha309;
        src24 <= 16'h4998;
        src25 <= 16'h2684;
        src26 <= 16'h670c;
        src27 <= 16'hf9dc;
        src28 <= 16'hd28a;
        src29 <= 16'h9749;
        src30 <= 16'h5bb;
        src31 <= 16'h5e93;
        src32 <= 16'h53a2;
        src33 <= 16'h6e10;
        src34 <= 16'h15c4;
        src35 <= 16'he142;
        src36 <= 16'h3569;
        src37 <= 16'h39a1;
        src38 <= 16'h182;
        src39 <= 16'h2efb;
        src40 <= 16'h379;
        src41 <= 16'h7465;
        src42 <= 16'h6882;
        src43 <= 16'hb4c6;
        src44 <= 16'h7839;
        src45 <= 16'he985;
        src46 <= 16'h8cd0;
        src47 <= 16'hb2e2;
        src48 <= 16'h6b1b;
        src49 <= 16'h9519;
        src50 <= 16'hb85d;
        src51 <= 16'hf009;
        src52 <= 16'h3e45;
        src53 <= 16'h43fd;
        src54 <= 16'h10b7;
        src55 <= 16'hfdae;
        src56 <= 16'hc9d1;
        src57 <= 16'ha3df;
        src58 <= 16'hfc2;
        src59 <= 16'h7d83;
        src60 <= 16'hb755;
        src61 <= 16'hd820;
        src62 <= 16'hafa0;
        src63 <= 16'h7f7;
        src64 <= 16'h868c;
        src65 <= 16'h9a3b;
        src66 <= 16'h902b;
        src67 <= 16'h20c0;
        src68 <= 16'h7b32;
        src69 <= 16'he9fb;
        src70 <= 16'h5f44;
        src71 <= 16'h6e1f;
        src72 <= 16'h34ca;
        src73 <= 16'h9ffc;
        src74 <= 16'h5b4e;
        src75 <= 16'ha196;
        src76 <= 16'h6f2d;
        src77 <= 16'he8c7;
        src78 <= 16'h3259;
        src79 <= 16'h1c2d;
        src80 <= 16'h8562;
        src81 <= 16'he1ad;
        src82 <= 16'hc096;
        src83 <= 16'he998;
        src84 <= 16'hbcb7;
        src85 <= 16'hbf02;
        src86 <= 16'h1e68;
        src87 <= 16'hddff;
        src88 <= 16'h2956;
        src89 <= 16'hcb05;
        src90 <= 16'h9d55;
        src91 <= 16'h344a;
        src92 <= 16'h901c;
        src93 <= 16'h3bc7;
        src94 <= 16'h217e;
        src95 <= 16'haaa2;
        src96 <= 16'h70b0;
        src97 <= 16'h3310;
        src98 <= 16'h3f01;
        src99 <= 16'hc48b;
        src100 <= 16'h8d0;
        src101 <= 16'h9846;
        src102 <= 16'h7ba4;
        src103 <= 16'h3c4d;
        src104 <= 16'h4c74;
        src105 <= 16'h90da;
        src106 <= 16'hd0b7;
        src107 <= 16'hc1ea;
        src108 <= 16'h25ed;
        src109 <= 16'hdef6;
        src110 <= 16'h1d77;
        src111 <= 16'h1f4c;
        src112 <= 16'ha314;
        src113 <= 16'h7e7b;
        src114 <= 16'h56b1;
        src115 <= 16'h8de7;
        src116 <= 16'h485f;
        src117 <= 16'h2300;
        src118 <= 16'h17eb;
        src119 <= 16'hd46;
        src120 <= 16'he2cf;
        src121 <= 16'h1826;
        src122 <= 16'h7853;
        src123 <= 16'h797d;
        src124 <= 16'hbf45;
        src125 <= 16'h58ea;
        src126 <= 16'hfe52;
        src127 <= 16'hfaaa;
        src128 <= 16'hd95;
        src129 <= 16'h9661;
        src130 <= 16'h9f98;
        src131 <= 16'hce32;
        src132 <= 16'h4a7a;
        src133 <= 16'h9a01;
        src134 <= 16'h5567;
        src135 <= 16'h997b;
        src136 <= 16'he4cf;
        src137 <= 16'he630;
        src138 <= 16'h4339;
        src139 <= 16'h6926;
        src140 <= 16'ha361;
        src141 <= 16'h2444;
        src142 <= 16'h202;
        src143 <= 16'he17c;
        src144 <= 16'h6961;
        src145 <= 16'hd55;
        src146 <= 16'h15a2;
        src147 <= 16'h20e1;
        src148 <= 16'hba33;
        src149 <= 16'h2ce0;
        src150 <= 16'h9dbe;
        src151 <= 16'hf44e;
        src152 <= 16'hab43;
        src153 <= 16'h5e60;
        src154 <= 16'h1a2b;
        src155 <= 16'h6b24;
        src156 <= 16'h64d7;
        src157 <= 16'h7df0;
        src158 <= 16'h5a65;
        src159 <= 16'hab1d;
        src160 <= 16'h43b1;
        src161 <= 16'hae7f;
        exp <= 24'h4d5861;
        #1
        src0 <= 16'hbec0;
        src1 <= 16'h1f64;
        src2 <= 16'h9b1d;
        src3 <= 16'h20ec;
        src4 <= 16'h5304;
        src5 <= 16'hb906;
        src6 <= 16'h97e0;
        src7 <= 16'hb14c;
        src8 <= 16'hfc01;
        src9 <= 16'hd284;
        src10 <= 16'h85e1;
        src11 <= 16'hebb;
        src12 <= 16'h3576;
        src13 <= 16'h75e1;
        src14 <= 16'hce1c;
        src15 <= 16'ha545;
        src16 <= 16'heaf5;
        src17 <= 16'h816b;
        src18 <= 16'hb0ad;
        src19 <= 16'h9b2f;
        src20 <= 16'hbe08;
        src21 <= 16'hbcd7;
        src22 <= 16'h1c6d;
        src23 <= 16'hb515;
        src24 <= 16'h9538;
        src25 <= 16'h4813;
        src26 <= 16'h6a2b;
        src27 <= 16'hd0f;
        src28 <= 16'h7f53;
        src29 <= 16'hadf6;
        src30 <= 16'hedba;
        src31 <= 16'h3f18;
        src32 <= 16'h305e;
        src33 <= 16'h1928;
        src34 <= 16'h4bf9;
        src35 <= 16'hf274;
        src36 <= 16'h1d7d;
        src37 <= 16'hcdb2;
        src38 <= 16'h90f5;
        src39 <= 16'h708b;
        src40 <= 16'haa07;
        src41 <= 16'h6188;
        src42 <= 16'h1fa;
        src43 <= 16'h4146;
        src44 <= 16'h9127;
        src45 <= 16'h1827;
        src46 <= 16'h13e5;
        src47 <= 16'h28b8;
        src48 <= 16'h7e6c;
        src49 <= 16'he34c;
        src50 <= 16'h23ad;
        src51 <= 16'hd2ad;
        src52 <= 16'h4cd5;
        src53 <= 16'ha358;
        src54 <= 16'ha40;
        src55 <= 16'hcf7e;
        src56 <= 16'h3f48;
        src57 <= 16'hc06a;
        src58 <= 16'h1209;
        src59 <= 16'hf62a;
        src60 <= 16'h6789;
        src61 <= 16'h8a02;
        src62 <= 16'h23bb;
        src63 <= 16'h1c27;
        src64 <= 16'hd539;
        src65 <= 16'hb9d3;
        src66 <= 16'h760c;
        src67 <= 16'h242e;
        src68 <= 16'h382f;
        src69 <= 16'h9f88;
        src70 <= 16'h2048;
        src71 <= 16'h8a2c;
        src72 <= 16'hc3d1;
        src73 <= 16'hb674;
        src74 <= 16'h4d5b;
        src75 <= 16'hbf08;
        src76 <= 16'h85f;
        src77 <= 16'hf578;
        src78 <= 16'h198a;
        src79 <= 16'hda86;
        src80 <= 16'h8bcb;
        src81 <= 16'h4eca;
        src82 <= 16'hb469;
        src83 <= 16'hbbdd;
        src84 <= 16'h4ebd;
        src85 <= 16'h804f;
        src86 <= 16'hecc8;
        src87 <= 16'h8c62;
        src88 <= 16'h76f;
        src89 <= 16'h49ae;
        src90 <= 16'h4811;
        src91 <= 16'hcbf1;
        src92 <= 16'hf8fc;
        src93 <= 16'heb73;
        src94 <= 16'hd8c2;
        src95 <= 16'h3933;
        src96 <= 16'h5f81;
        src97 <= 16'hb330;
        src98 <= 16'hddfc;
        src99 <= 16'h7bbf;
        src100 <= 16'h90da;
        src101 <= 16'h54e2;
        src102 <= 16'h22a9;
        src103 <= 16'h284a;
        src104 <= 16'hf063;
        src105 <= 16'h8252;
        src106 <= 16'h1f18;
        src107 <= 16'h5d70;
        src108 <= 16'hea93;
        src109 <= 16'h9a40;
        src110 <= 16'h6d74;
        src111 <= 16'h878;
        src112 <= 16'hffa3;
        src113 <= 16'h9259;
        src114 <= 16'h7928;
        src115 <= 16'h6008;
        src116 <= 16'h4562;
        src117 <= 16'h74ab;
        src118 <= 16'haf6c;
        src119 <= 16'h1de5;
        src120 <= 16'he73d;
        src121 <= 16'h410c;
        src122 <= 16'h6c84;
        src123 <= 16'h2b88;
        src124 <= 16'hd17;
        src125 <= 16'h1473;
        src126 <= 16'h48aa;
        src127 <= 16'h3566;
        src128 <= 16'hf75d;
        src129 <= 16'hdbde;
        src130 <= 16'hc625;
        src131 <= 16'hbad9;
        src132 <= 16'h4637;
        src133 <= 16'hbee2;
        src134 <= 16'h6fab;
        src135 <= 16'h2271;
        src136 <= 16'h22e0;
        src137 <= 16'hb3c3;
        src138 <= 16'h9bf9;
        src139 <= 16'h8347;
        src140 <= 16'hf83;
        src141 <= 16'hd3f3;
        src142 <= 16'hca7;
        src143 <= 16'hed99;
        src144 <= 16'h9a48;
        src145 <= 16'h45b6;
        src146 <= 16'hfebf;
        src147 <= 16'hfa68;
        src148 <= 16'hbbf0;
        src149 <= 16'h6177;
        src150 <= 16'h3035;
        src151 <= 16'hbe3f;
        src152 <= 16'hdf8a;
        src153 <= 16'h1afb;
        src154 <= 16'h879c;
        src155 <= 16'h782b;
        src156 <= 16'h5be1;
        src157 <= 16'h6858;
        src158 <= 16'h2544;
        src159 <= 16'h6651;
        src160 <= 16'h9e95;
        src161 <= 16'h1ec5;
        exp <= 24'h4ec0c3;
        #1
        src0 <= 16'h8bf6;
        src1 <= 16'h9ac0;
        src2 <= 16'h1ae4;
        src3 <= 16'h8860;
        src4 <= 16'hc68;
        src5 <= 16'haa61;
        src6 <= 16'hcd9c;
        src7 <= 16'hd47d;
        src8 <= 16'h2afc;
        src9 <= 16'hd33f;
        src10 <= 16'h214;
        src11 <= 16'h6f39;
        src12 <= 16'h42a9;
        src13 <= 16'h13ba;
        src14 <= 16'h15d9;
        src15 <= 16'h60b2;
        src16 <= 16'h6c4c;
        src17 <= 16'h68ef;
        src18 <= 16'hc809;
        src19 <= 16'ha360;
        src20 <= 16'h52d7;
        src21 <= 16'hb26b;
        src22 <= 16'he77b;
        src23 <= 16'h1a;
        src24 <= 16'he5e9;
        src25 <= 16'h9358;
        src26 <= 16'h5613;
        src27 <= 16'h6a06;
        src28 <= 16'had86;
        src29 <= 16'h382b;
        src30 <= 16'h53c4;
        src31 <= 16'h235c;
        src32 <= 16'h512f;
        src33 <= 16'h4774;
        src34 <= 16'h8c72;
        src35 <= 16'hda5f;
        src36 <= 16'h5b66;
        src37 <= 16'hda7d;
        src38 <= 16'hcc19;
        src39 <= 16'h3f6d;
        src40 <= 16'hd083;
        src41 <= 16'h97a;
        src42 <= 16'h4c34;
        src43 <= 16'h1b2b;
        src44 <= 16'h6059;
        src45 <= 16'hf8fe;
        src46 <= 16'h913b;
        src47 <= 16'h2cd6;
        src48 <= 16'h8b82;
        src49 <= 16'h3efd;
        src50 <= 16'hf716;
        src51 <= 16'h168b;
        src52 <= 16'h28d3;
        src53 <= 16'h9ecb;
        src54 <= 16'h357b;
        src55 <= 16'h40b8;
        src56 <= 16'h53b5;
        src57 <= 16'h3fd2;
        src58 <= 16'hb5aa;
        src59 <= 16'h3ed7;
        src60 <= 16'hdc10;
        src61 <= 16'h496f;
        src62 <= 16'hb2b0;
        src63 <= 16'h7fa1;
        src64 <= 16'hc8d5;
        src65 <= 16'h5997;
        src66 <= 16'ha187;
        src67 <= 16'h42d9;
        src68 <= 16'hccd3;
        src69 <= 16'hb459;
        src70 <= 16'he82;
        src71 <= 16'hdb96;
        src72 <= 16'h5302;
        src73 <= 16'h449f;
        src74 <= 16'h2982;
        src75 <= 16'h556c;
        src76 <= 16'h28e9;
        src77 <= 16'h782d;
        src78 <= 16'h7fe4;
        src79 <= 16'h6ebd;
        src80 <= 16'h90c9;
        src81 <= 16'he928;
        src82 <= 16'h1efb;
        src83 <= 16'h2096;
        src84 <= 16'h1839;
        src85 <= 16'h1bfb;
        src86 <= 16'haf11;
        src87 <= 16'h8ce2;
        src88 <= 16'h707f;
        src89 <= 16'he37f;
        src90 <= 16'h9471;
        src91 <= 16'h1ce7;
        src92 <= 16'h8cf4;
        src93 <= 16'he122;
        src94 <= 16'h71d9;
        src95 <= 16'h8ba9;
        src96 <= 16'hf39b;
        src97 <= 16'h4674;
        src98 <= 16'h6f6f;
        src99 <= 16'hd19a;
        src100 <= 16'hbfed;
        src101 <= 16'hee4;
        src102 <= 16'h19ac;
        src103 <= 16'h7cbf;
        src104 <= 16'h3991;
        src105 <= 16'h99bd;
        src106 <= 16'hc3b3;
        src107 <= 16'h2a6c;
        src108 <= 16'h4bb5;
        src109 <= 16'h48a7;
        src110 <= 16'hda58;
        src111 <= 16'h9147;
        src112 <= 16'hd433;
        src113 <= 16'hff6a;
        src114 <= 16'h85f4;
        src115 <= 16'hfae1;
        src116 <= 16'hba1e;
        src117 <= 16'h2180;
        src118 <= 16'h38bf;
        src119 <= 16'h4ba6;
        src120 <= 16'hcfb9;
        src121 <= 16'hf958;
        src122 <= 16'h5905;
        src123 <= 16'hc72e;
        src124 <= 16'h4661;
        src125 <= 16'hf324;
        src126 <= 16'hd55c;
        src127 <= 16'h8544;
        src128 <= 16'hdce6;
        src129 <= 16'hf5d;
        src130 <= 16'h5b6d;
        src131 <= 16'h26a8;
        src132 <= 16'h7549;
        src133 <= 16'h66bd;
        src134 <= 16'h343;
        src135 <= 16'h524b;
        src136 <= 16'hee8c;
        src137 <= 16'h6d3c;
        src138 <= 16'h438a;
        src139 <= 16'h704c;
        src140 <= 16'hc773;
        src141 <= 16'h90bd;
        src142 <= 16'h8ec1;
        src143 <= 16'h22ed;
        src144 <= 16'h2c9e;
        src145 <= 16'h18f4;
        src146 <= 16'ha08b;
        src147 <= 16'hbbf;
        src148 <= 16'h385e;
        src149 <= 16'h51ae;
        src150 <= 16'ha6c2;
        src151 <= 16'h1c4c;
        src152 <= 16'h606b;
        src153 <= 16'hf861;
        src154 <= 16'hb8ab;
        src155 <= 16'h828;
        src156 <= 16'h4b99;
        src157 <= 16'h4f3;
        src158 <= 16'hfc73;
        src159 <= 16'h90e0;
        src160 <= 16'hf5ae;
        src161 <= 16'hc223;
        exp <= 24'h4be096;
        #1
        src0 <= 16'he687;
        src1 <= 16'h4f1f;
        src2 <= 16'h289d;
        src3 <= 16'h2a60;
        src4 <= 16'h8aaf;
        src5 <= 16'h4b6;
        src6 <= 16'h2c6;
        src7 <= 16'hc33a;
        src8 <= 16'ha26b;
        src9 <= 16'hec84;
        src10 <= 16'hc2e;
        src11 <= 16'hcb91;
        src12 <= 16'h9e3c;
        src13 <= 16'h2ee0;
        src14 <= 16'hb1d3;
        src15 <= 16'h8478;
        src16 <= 16'h1cec;
        src17 <= 16'h64c2;
        src18 <= 16'h2789;
        src19 <= 16'h34a8;
        src20 <= 16'h2c90;
        src21 <= 16'h4c0a;
        src22 <= 16'hc4a2;
        src23 <= 16'he640;
        src24 <= 16'h23b3;
        src25 <= 16'h5f9f;
        src26 <= 16'h4bdf;
        src27 <= 16'h583f;
        src28 <= 16'h7ec3;
        src29 <= 16'ha0dc;
        src30 <= 16'hdf5c;
        src31 <= 16'hcf5f;
        src32 <= 16'h998;
        src33 <= 16'h67dc;
        src34 <= 16'heaea;
        src35 <= 16'h2707;
        src36 <= 16'h21a4;
        src37 <= 16'h2142;
        src38 <= 16'h4a40;
        src39 <= 16'h40e;
        src40 <= 16'h87c1;
        src41 <= 16'hb21e;
        src42 <= 16'hbe68;
        src43 <= 16'hb047;
        src44 <= 16'hc907;
        src45 <= 16'h97b0;
        src46 <= 16'hf9b7;
        src47 <= 16'h35cc;
        src48 <= 16'h6e37;
        src49 <= 16'hd31f;
        src50 <= 16'hee26;
        src51 <= 16'hbbfc;
        src52 <= 16'h7e16;
        src53 <= 16'hcdfd;
        src54 <= 16'hdbe3;
        src55 <= 16'h72c1;
        src56 <= 16'h6e0c;
        src57 <= 16'he499;
        src58 <= 16'hdfe8;
        src59 <= 16'h5b3b;
        src60 <= 16'h3e74;
        src61 <= 16'hc2d0;
        src62 <= 16'hd95f;
        src63 <= 16'h254d;
        src64 <= 16'h115b;
        src65 <= 16'h7e78;
        src66 <= 16'hb7c2;
        src67 <= 16'h5848;
        src68 <= 16'hd1a5;
        src69 <= 16'h5d78;
        src70 <= 16'h8afc;
        src71 <= 16'h4498;
        src72 <= 16'h54a7;
        src73 <= 16'h37b1;
        src74 <= 16'hf619;
        src75 <= 16'h57fe;
        src76 <= 16'hc93;
        src77 <= 16'h945d;
        src78 <= 16'heaee;
        src79 <= 16'hca72;
        src80 <= 16'h6678;
        src81 <= 16'hab95;
        src82 <= 16'hedf7;
        src83 <= 16'h1641;
        src84 <= 16'h6637;
        src85 <= 16'hf206;
        src86 <= 16'hd6a4;
        src87 <= 16'hfa2d;
        src88 <= 16'h8f42;
        src89 <= 16'h1ff2;
        src90 <= 16'h3d8;
        src91 <= 16'h3f26;
        src92 <= 16'h2e10;
        src93 <= 16'h3915;
        src94 <= 16'ha1af;
        src95 <= 16'h2e20;
        src96 <= 16'hb37f;
        src97 <= 16'h9237;
        src98 <= 16'hf6cc;
        src99 <= 16'hbcd6;
        src100 <= 16'h6983;
        src101 <= 16'h31fe;
        src102 <= 16'he27a;
        src103 <= 16'h2348;
        src104 <= 16'h6126;
        src105 <= 16'h1b8b;
        src106 <= 16'hfdbb;
        src107 <= 16'h9da4;
        src108 <= 16'h7b5a;
        src109 <= 16'h4094;
        src110 <= 16'he371;
        src111 <= 16'hc3bb;
        src112 <= 16'ha8a0;
        src113 <= 16'h3e9a;
        src114 <= 16'h6d05;
        src115 <= 16'hbceb;
        src116 <= 16'h735f;
        src117 <= 16'h90ac;
        src118 <= 16'he71c;
        src119 <= 16'h5f4c;
        src120 <= 16'h8f2b;
        src121 <= 16'h791b;
        src122 <= 16'ha795;
        src123 <= 16'h1d63;
        src124 <= 16'h88de;
        src125 <= 16'hc327;
        src126 <= 16'hdfd9;
        src127 <= 16'h23c1;
        src128 <= 16'h4e6d;
        src129 <= 16'ha3f0;
        src130 <= 16'hed88;
        src131 <= 16'hb03;
        src132 <= 16'h25d4;
        src133 <= 16'h3117;
        src134 <= 16'h9108;
        src135 <= 16'hfe86;
        src136 <= 16'h11a4;
        src137 <= 16'h618;
        src138 <= 16'h70e;
        src139 <= 16'hbe4f;
        src140 <= 16'h8907;
        src141 <= 16'h3c0;
        src142 <= 16'hfe46;
        src143 <= 16'hb6c0;
        src144 <= 16'h2ac8;
        src145 <= 16'h7c07;
        src146 <= 16'hc035;
        src147 <= 16'h61e4;
        src148 <= 16'h4cbc;
        src149 <= 16'hf97f;
        src150 <= 16'h1dcd;
        src151 <= 16'h63a6;
        src152 <= 16'hcf29;
        src153 <= 16'hcbde;
        src154 <= 16'h1b23;
        src155 <= 16'hcfe;
        src156 <= 16'h6e8e;
        src157 <= 16'h3b3d;
        src158 <= 16'h9fc0;
        src159 <= 16'hff21;
        src160 <= 16'hd4c5;
        src161 <= 16'h87d2;
        exp <= 24'h504fd7;
        #1
        src0 <= 16'hd666;
        src1 <= 16'ha79e;
        src2 <= 16'h77d;
        src3 <= 16'hf86a;
        src4 <= 16'h9192;
        src5 <= 16'h7c37;
        src6 <= 16'h4d5e;
        src7 <= 16'h90cd;
        src8 <= 16'he86c;
        src9 <= 16'h62d8;
        src10 <= 16'hb278;
        src11 <= 16'h6531;
        src12 <= 16'h3b39;
        src13 <= 16'hb8ab;
        src14 <= 16'h720a;
        src15 <= 16'h18d8;
        src16 <= 16'habbf;
        src17 <= 16'h571d;
        src18 <= 16'h1c03;
        src19 <= 16'h558d;
        src20 <= 16'h348c;
        src21 <= 16'h3aa1;
        src22 <= 16'hcdaf;
        src23 <= 16'h3d72;
        src24 <= 16'h42c2;
        src25 <= 16'hdf55;
        src26 <= 16'h7d1;
        src27 <= 16'hd062;
        src28 <= 16'h8c93;
        src29 <= 16'h3d38;
        src30 <= 16'h59a0;
        src31 <= 16'h27ec;
        src32 <= 16'he2df;
        src33 <= 16'h738c;
        src34 <= 16'hed8f;
        src35 <= 16'he816;
        src36 <= 16'h6cde;
        src37 <= 16'hecec;
        src38 <= 16'hfbf6;
        src39 <= 16'h9f0c;
        src40 <= 16'h46f5;
        src41 <= 16'h5477;
        src42 <= 16'h23b1;
        src43 <= 16'haa25;
        src44 <= 16'h78e3;
        src45 <= 16'h6c1;
        src46 <= 16'h8782;
        src47 <= 16'he51c;
        src48 <= 16'h2058;
        src49 <= 16'hf520;
        src50 <= 16'h1873;
        src51 <= 16'hcc70;
        src52 <= 16'hbe2a;
        src53 <= 16'ha2e7;
        src54 <= 16'h99af;
        src55 <= 16'h1f4b;
        src56 <= 16'hb0e9;
        src57 <= 16'h6e37;
        src58 <= 16'h2f06;
        src59 <= 16'had9c;
        src60 <= 16'hec5;
        src61 <= 16'h9552;
        src62 <= 16'hebdd;
        src63 <= 16'h5588;
        src64 <= 16'h642;
        src65 <= 16'h3c1a;
        src66 <= 16'hf15b;
        src67 <= 16'h59db;
        src68 <= 16'h8610;
        src69 <= 16'h78b3;
        src70 <= 16'h2208;
        src71 <= 16'hefeb;
        src72 <= 16'h530b;
        src73 <= 16'h8d2c;
        src74 <= 16'hc5cf;
        src75 <= 16'h7837;
        src76 <= 16'hee75;
        src77 <= 16'hf948;
        src78 <= 16'h67cc;
        src79 <= 16'he755;
        src80 <= 16'h810a;
        src81 <= 16'ha55c;
        src82 <= 16'hfec6;
        src83 <= 16'h5761;
        src84 <= 16'h1b44;
        src85 <= 16'heac4;
        src86 <= 16'hc649;
        src87 <= 16'hb9e7;
        src88 <= 16'h2494;
        src89 <= 16'h1fc3;
        src90 <= 16'h343c;
        src91 <= 16'ha4a2;
        src92 <= 16'h547f;
        src93 <= 16'hed6b;
        src94 <= 16'hf1a2;
        src95 <= 16'h6f08;
        src96 <= 16'h8a5e;
        src97 <= 16'he508;
        src98 <= 16'h2854;
        src99 <= 16'h4b3d;
        src100 <= 16'hc061;
        src101 <= 16'h8b4;
        src102 <= 16'hbd17;
        src103 <= 16'hc74c;
        src104 <= 16'h1083;
        src105 <= 16'hb9f9;
        src106 <= 16'h787e;
        src107 <= 16'ha68d;
        src108 <= 16'h4801;
        src109 <= 16'h31f6;
        src110 <= 16'h1f0f;
        src111 <= 16'hb7c;
        src112 <= 16'hcf23;
        src113 <= 16'hcb36;
        src114 <= 16'h2ee3;
        src115 <= 16'h89d;
        src116 <= 16'h69ff;
        src117 <= 16'h5c8d;
        src118 <= 16'h730e;
        src119 <= 16'ha64b;
        src120 <= 16'hdf68;
        src121 <= 16'h18c8;
        src122 <= 16'h6960;
        src123 <= 16'h2fa5;
        src124 <= 16'h90ef;
        src125 <= 16'h458d;
        src126 <= 16'h4613;
        src127 <= 16'h331d;
        src128 <= 16'h6f5b;
        src129 <= 16'hbe2d;
        src130 <= 16'h923b;
        src131 <= 16'h41d2;
        src132 <= 16'h6846;
        src133 <= 16'h3ab0;
        src134 <= 16'hbefc;
        src135 <= 16'hd6fb;
        src136 <= 16'h97a1;
        src137 <= 16'h68fc;
        src138 <= 16'h5036;
        src139 <= 16'h9016;
        src140 <= 16'h782c;
        src141 <= 16'h52e2;
        src142 <= 16'hd3aa;
        src143 <= 16'h481f;
        src144 <= 16'hf417;
        src145 <= 16'h8d52;
        src146 <= 16'h8d0d;
        src147 <= 16'he895;
        src148 <= 16'h321f;
        src149 <= 16'hd865;
        src150 <= 16'h9b0f;
        src151 <= 16'hcb79;
        src152 <= 16'h1832;
        src153 <= 16'hfc94;
        src154 <= 16'hfb19;
        src155 <= 16'h276a;
        src156 <= 16'h4222;
        src157 <= 16'h4f33;
        src158 <= 16'h5a5c;
        src159 <= 16'h3559;
        src160 <= 16'h53d;
        src161 <= 16'h2aa2;
        exp <= 24'h4fe584;
        #1
        src0 <= 16'h2d41;
        src1 <= 16'hf205;
        src2 <= 16'hd833;
        src3 <= 16'h3dae;
        src4 <= 16'h7c91;
        src5 <= 16'h55db;
        src6 <= 16'h9766;
        src7 <= 16'h6e76;
        src8 <= 16'hc4eb;
        src9 <= 16'hd3ea;
        src10 <= 16'heb64;
        src11 <= 16'hfa46;
        src12 <= 16'h252e;
        src13 <= 16'h3790;
        src14 <= 16'h4aa0;
        src15 <= 16'h761d;
        src16 <= 16'h3d5f;
        src17 <= 16'hbbb2;
        src18 <= 16'hd4a;
        src19 <= 16'h1737;
        src20 <= 16'h9734;
        src21 <= 16'ha175;
        src22 <= 16'h212b;
        src23 <= 16'h55ae;
        src24 <= 16'h75ff;
        src25 <= 16'h999e;
        src26 <= 16'h2e90;
        src27 <= 16'h10f9;
        src28 <= 16'hf1c9;
        src29 <= 16'h2857;
        src30 <= 16'he09f;
        src31 <= 16'hf63a;
        src32 <= 16'h6749;
        src33 <= 16'hd9;
        src34 <= 16'h2426;
        src35 <= 16'h727f;
        src36 <= 16'h8195;
        src37 <= 16'h8d7d;
        src38 <= 16'hb9bf;
        src39 <= 16'h6bd5;
        src40 <= 16'ha282;
        src41 <= 16'h90b0;
        src42 <= 16'h8d9a;
        src43 <= 16'hb72c;
        src44 <= 16'h62ba;
        src45 <= 16'h64d3;
        src46 <= 16'hc559;
        src47 <= 16'hbb79;
        src48 <= 16'h7b2d;
        src49 <= 16'h9d00;
        src50 <= 16'hce66;
        src51 <= 16'h80b1;
        src52 <= 16'hc1a;
        src53 <= 16'he754;
        src54 <= 16'he768;
        src55 <= 16'hf156;
        src56 <= 16'hb69c;
        src57 <= 16'h7db1;
        src58 <= 16'h8dda;
        src59 <= 16'h695f;
        src60 <= 16'h1758;
        src61 <= 16'ha13c;
        src62 <= 16'h22aa;
        src63 <= 16'hd4f6;
        src64 <= 16'hc9a6;
        src65 <= 16'hfc49;
        src66 <= 16'ha46d;
        src67 <= 16'h5e94;
        src68 <= 16'h2046;
        src69 <= 16'h2de;
        src70 <= 16'h868e;
        src71 <= 16'hc1d1;
        src72 <= 16'h6f25;
        src73 <= 16'h2669;
        src74 <= 16'ha0d0;
        src75 <= 16'h1590;
        src76 <= 16'hcc3e;
        src77 <= 16'he909;
        src78 <= 16'h56e5;
        src79 <= 16'h4c5a;
        src80 <= 16'h6f4d;
        src81 <= 16'hc081;
        src82 <= 16'h76e9;
        src83 <= 16'hf19d;
        src84 <= 16'h3147;
        src85 <= 16'h57ab;
        src86 <= 16'h3ac6;
        src87 <= 16'h9baf;
        src88 <= 16'h9a4a;
        src89 <= 16'h14f7;
        src90 <= 16'hf4d0;
        src91 <= 16'h580d;
        src92 <= 16'h911a;
        src93 <= 16'h1eb5;
        src94 <= 16'hdea9;
        src95 <= 16'h806f;
        src96 <= 16'hd948;
        src97 <= 16'hbc5d;
        src98 <= 16'h8976;
        src99 <= 16'h6037;
        src100 <= 16'h6d2f;
        src101 <= 16'h116b;
        src102 <= 16'h7553;
        src103 <= 16'hd44c;
        src104 <= 16'hcdd4;
        src105 <= 16'h1531;
        src106 <= 16'ha048;
        src107 <= 16'h334a;
        src108 <= 16'h99c9;
        src109 <= 16'h43d4;
        src110 <= 16'hff82;
        src111 <= 16'h3d7b;
        src112 <= 16'h7996;
        src113 <= 16'h189c;
        src114 <= 16'hf2a0;
        src115 <= 16'hfce5;
        src116 <= 16'hadfd;
        src117 <= 16'h6fe7;
        src118 <= 16'h39da;
        src119 <= 16'h429;
        src120 <= 16'hfa37;
        src121 <= 16'h7c3c;
        src122 <= 16'h5c87;
        src123 <= 16'h8ade;
        src124 <= 16'h5dfb;
        src125 <= 16'h4e6c;
        src126 <= 16'h711;
        src127 <= 16'h103e;
        src128 <= 16'hbec9;
        src129 <= 16'h445f;
        src130 <= 16'h3aab;
        src131 <= 16'hf295;
        src132 <= 16'h6d45;
        src133 <= 16'he48;
        src134 <= 16'h7cb3;
        src135 <= 16'h7ead;
        src136 <= 16'he06c;
        src137 <= 16'h75f;
        src138 <= 16'h4d2d;
        src139 <= 16'hfdee;
        src140 <= 16'h41df;
        src141 <= 16'h9ad3;
        src142 <= 16'h9f9e;
        src143 <= 16'h4268;
        src144 <= 16'ha411;
        src145 <= 16'hb823;
        src146 <= 16'h4cd1;
        src147 <= 16'haf2;
        src148 <= 16'hfc70;
        src149 <= 16'hdfff;
        src150 <= 16'he93b;
        src151 <= 16'h8155;
        src152 <= 16'h5fdb;
        src153 <= 16'hbc50;
        src154 <= 16'hfe8b;
        src155 <= 16'heb6f;
        src156 <= 16'h3418;
        src157 <= 16'h189d;
        src158 <= 16'h6b3d;
        src159 <= 16'h47d;
        src160 <= 16'h7998;
        src161 <= 16'he54a;
        exp <= 24'h516278;
        #1
        src0 <= 16'hdb0d;
        src1 <= 16'h4336;
        src2 <= 16'h2df8;
        src3 <= 16'hdc8b;
        src4 <= 16'hf877;
        src5 <= 16'h5f00;
        src6 <= 16'h88a6;
        src7 <= 16'ha7f5;
        src8 <= 16'h167;
        src9 <= 16'h4481;
        src10 <= 16'h371c;
        src11 <= 16'h11df;
        src12 <= 16'h602c;
        src13 <= 16'h921b;
        src14 <= 16'hbee0;
        src15 <= 16'hcb2;
        src16 <= 16'hc4ac;
        src17 <= 16'ha184;
        src18 <= 16'hbc2;
        src19 <= 16'h1c6d;
        src20 <= 16'h138f;
        src21 <= 16'hac08;
        src22 <= 16'h5ceb;
        src23 <= 16'ha521;
        src24 <= 16'h8921;
        src25 <= 16'h5c6;
        src26 <= 16'h75d8;
        src27 <= 16'h6be;
        src28 <= 16'hab1;
        src29 <= 16'h2085;
        src30 <= 16'h525d;
        src31 <= 16'hf08b;
        src32 <= 16'hbe44;
        src33 <= 16'h33b9;
        src34 <= 16'h20a7;
        src35 <= 16'had70;
        src36 <= 16'hdca0;
        src37 <= 16'he15c;
        src38 <= 16'h75ea;
        src39 <= 16'h705;
        src40 <= 16'h6320;
        src41 <= 16'hef7a;
        src42 <= 16'hb14b;
        src43 <= 16'h83a7;
        src44 <= 16'h7962;
        src45 <= 16'h9454;
        src46 <= 16'h226b;
        src47 <= 16'h9d51;
        src48 <= 16'h64a8;
        src49 <= 16'h4fd1;
        src50 <= 16'h5ae2;
        src51 <= 16'h5151;
        src52 <= 16'hf4b4;
        src53 <= 16'h6bb9;
        src54 <= 16'h5d7a;
        src55 <= 16'hc012;
        src56 <= 16'h693f;
        src57 <= 16'h4a8f;
        src58 <= 16'h609c;
        src59 <= 16'hf6b2;
        src60 <= 16'hc529;
        src61 <= 16'h8ba3;
        src62 <= 16'ha4a4;
        src63 <= 16'h1619;
        src64 <= 16'ha288;
        src65 <= 16'h8b5a;
        src66 <= 16'h17c;
        src67 <= 16'h959d;
        src68 <= 16'h1d88;
        src69 <= 16'hbf8d;
        src70 <= 16'h9b96;
        src71 <= 16'hd81c;
        src72 <= 16'hbd6e;
        src73 <= 16'hc16e;
        src74 <= 16'haf6;
        src75 <= 16'h526e;
        src76 <= 16'hdbcc;
        src77 <= 16'h2099;
        src78 <= 16'he963;
        src79 <= 16'h4fdb;
        src80 <= 16'h48f7;
        src81 <= 16'hb14;
        src82 <= 16'h5446;
        src83 <= 16'h7e79;
        src84 <= 16'h4fec;
        src85 <= 16'h90f1;
        src86 <= 16'h6544;
        src87 <= 16'hcaf6;
        src88 <= 16'h78a7;
        src89 <= 16'hc070;
        src90 <= 16'hf61e;
        src91 <= 16'ha151;
        src92 <= 16'hb0de;
        src93 <= 16'hf4b0;
        src94 <= 16'h155;
        src95 <= 16'h230a;
        src96 <= 16'hd8fd;
        src97 <= 16'hf124;
        src98 <= 16'h88b5;
        src99 <= 16'hba12;
        src100 <= 16'hb04d;
        src101 <= 16'h28e0;
        src102 <= 16'h1214;
        src103 <= 16'h65c9;
        src104 <= 16'h8c57;
        src105 <= 16'he287;
        src106 <= 16'h712d;
        src107 <= 16'h4ce6;
        src108 <= 16'h5ff1;
        src109 <= 16'h9273;
        src110 <= 16'h5df;
        src111 <= 16'h76ad;
        src112 <= 16'h8bf2;
        src113 <= 16'h5b0f;
        src114 <= 16'h4e6b;
        src115 <= 16'hbc26;
        src116 <= 16'h4ca9;
        src117 <= 16'h3ca4;
        src118 <= 16'h710b;
        src119 <= 16'h6116;
        src120 <= 16'h10cb;
        src121 <= 16'h4eb2;
        src122 <= 16'ha682;
        src123 <= 16'h1ea1;
        src124 <= 16'hac9d;
        src125 <= 16'h52d9;
        src126 <= 16'h2bf0;
        src127 <= 16'h65e1;
        src128 <= 16'h1f6e;
        src129 <= 16'h3f36;
        src130 <= 16'h2a28;
        src131 <= 16'h10ee;
        src132 <= 16'h7116;
        src133 <= 16'hb57e;
        src134 <= 16'hebe2;
        src135 <= 16'h3868;
        src136 <= 16'h8205;
        src137 <= 16'ha7dc;
        src138 <= 16'h683c;
        src139 <= 16'h6b62;
        src140 <= 16'ha29e;
        src141 <= 16'h773a;
        src142 <= 16'hc81f;
        src143 <= 16'h981c;
        src144 <= 16'hec86;
        src145 <= 16'hd1c9;
        src146 <= 16'hdbdd;
        src147 <= 16'h1638;
        src148 <= 16'h832f;
        src149 <= 16'h478f;
        src150 <= 16'h3bd2;
        src151 <= 16'h37d9;
        src152 <= 16'he751;
        src153 <= 16'hb7d6;
        src154 <= 16'hd80c;
        src155 <= 16'h1d15;
        src156 <= 16'h5171;
        src157 <= 16'hcd1b;
        src158 <= 16'hd099;
        src159 <= 16'hca72;
        src160 <= 16'h4cff;
        src161 <= 16'h1c0a;
        exp <= 24'h4c050a;
        #1
        src0 <= 16'h462e;
        src1 <= 16'h8964;
        src2 <= 16'h68dc;
        src3 <= 16'hafa;
        src4 <= 16'hc087;
        src5 <= 16'h7de3;
        src6 <= 16'ha726;
        src7 <= 16'hfe57;
        src8 <= 16'h107a;
        src9 <= 16'h3568;
        src10 <= 16'h9a07;
        src11 <= 16'h429b;
        src12 <= 16'h71c7;
        src13 <= 16'h2b36;
        src14 <= 16'h2da1;
        src15 <= 16'h7551;
        src16 <= 16'h77e1;
        src17 <= 16'hded0;
        src18 <= 16'hed76;
        src19 <= 16'hce30;
        src20 <= 16'hfd74;
        src21 <= 16'h29d5;
        src22 <= 16'h2830;
        src23 <= 16'h2e74;
        src24 <= 16'h35dc;
        src25 <= 16'h3fc2;
        src26 <= 16'h79a5;
        src27 <= 16'h21a;
        src28 <= 16'h3fe9;
        src29 <= 16'h357d;
        src30 <= 16'h9e78;
        src31 <= 16'hc913;
        src32 <= 16'h3d21;
        src33 <= 16'h576b;
        src34 <= 16'h25e0;
        src35 <= 16'h728b;
        src36 <= 16'h2d37;
        src37 <= 16'hcad8;
        src38 <= 16'h3f3c;
        src39 <= 16'h44dd;
        src40 <= 16'h528b;
        src41 <= 16'h3e13;
        src42 <= 16'h9215;
        src43 <= 16'h3e13;
        src44 <= 16'h526;
        src45 <= 16'h4347;
        src46 <= 16'hb2c9;
        src47 <= 16'h51cb;
        src48 <= 16'h1887;
        src49 <= 16'h7db1;
        src50 <= 16'heb70;
        src51 <= 16'hd71d;
        src52 <= 16'h599c;
        src53 <= 16'he73a;
        src54 <= 16'h2194;
        src55 <= 16'h1f8;
        src56 <= 16'hb822;
        src57 <= 16'h43e0;
        src58 <= 16'h8d0a;
        src59 <= 16'h787c;
        src60 <= 16'h4bbe;
        src61 <= 16'h73e3;
        src62 <= 16'hec6f;
        src63 <= 16'h2618;
        src64 <= 16'hd214;
        src65 <= 16'hc473;
        src66 <= 16'hccd6;
        src67 <= 16'h1731;
        src68 <= 16'h7d73;
        src69 <= 16'h3953;
        src70 <= 16'h2a7;
        src71 <= 16'h813e;
        src72 <= 16'h9ca3;
        src73 <= 16'h85e8;
        src74 <= 16'hc471;
        src75 <= 16'h3c6c;
        src76 <= 16'hb3b1;
        src77 <= 16'haf49;
        src78 <= 16'hbd6a;
        src79 <= 16'hf515;
        src80 <= 16'hb2be;
        src81 <= 16'hcd08;
        src82 <= 16'h23c;
        src83 <= 16'h26d6;
        src84 <= 16'hdf14;
        src85 <= 16'h2952;
        src86 <= 16'h2130;
        src87 <= 16'h993f;
        src88 <= 16'hc0ca;
        src89 <= 16'h184d;
        src90 <= 16'h83b4;
        src91 <= 16'h1fda;
        src92 <= 16'he39;
        src93 <= 16'h217a;
        src94 <= 16'ha900;
        src95 <= 16'hb5e;
        src96 <= 16'he20c;
        src97 <= 16'h4a1d;
        src98 <= 16'h1d69;
        src99 <= 16'ha4e6;
        src100 <= 16'hf9a6;
        src101 <= 16'h3c39;
        src102 <= 16'hb69b;
        src103 <= 16'h3279;
        src104 <= 16'h812f;
        src105 <= 16'h7098;
        src106 <= 16'hbde4;
        src107 <= 16'h590a;
        src108 <= 16'hb513;
        src109 <= 16'h18d5;
        src110 <= 16'hd19b;
        src111 <= 16'h9390;
        src112 <= 16'h777b;
        src113 <= 16'hf411;
        src114 <= 16'he29;
        src115 <= 16'h589e;
        src116 <= 16'h493a;
        src117 <= 16'hac5e;
        src118 <= 16'h3e07;
        src119 <= 16'h7514;
        src120 <= 16'h29e1;
        src121 <= 16'hcbaa;
        src122 <= 16'h923e;
        src123 <= 16'h2c9e;
        src124 <= 16'hc93c;
        src125 <= 16'h1487;
        src126 <= 16'h8a57;
        src127 <= 16'h442c;
        src128 <= 16'h6046;
        src129 <= 16'hb294;
        src130 <= 16'ha25e;
        src131 <= 16'h9a04;
        src132 <= 16'hc992;
        src133 <= 16'he3bf;
        src134 <= 16'h37fa;
        src135 <= 16'h8603;
        src136 <= 16'hfc74;
        src137 <= 16'h4220;
        src138 <= 16'hadb0;
        src139 <= 16'heed5;
        src140 <= 16'h7cc;
        src141 <= 16'h5ab8;
        src142 <= 16'h630a;
        src143 <= 16'h133b;
        src144 <= 16'h1166;
        src145 <= 16'h1bea;
        src146 <= 16'h7f84;
        src147 <= 16'he7e6;
        src148 <= 16'h7689;
        src149 <= 16'h9412;
        src150 <= 16'hd3a6;
        src151 <= 16'hd56;
        src152 <= 16'h2e38;
        src153 <= 16'hab97;
        src154 <= 16'h9744;
        src155 <= 16'h33ae;
        src156 <= 16'hc551;
        src157 <= 16'h3543;
        src158 <= 16'hccf2;
        src159 <= 16'h44a2;
        src160 <= 16'h1707;
        src161 <= 16'hfe95;
        exp <= 24'h4964b6;
        #1
        src0 <= 16'h6eed;
        src1 <= 16'h7804;
        src2 <= 16'hc68;
        src3 <= 16'h3d1a;
        src4 <= 16'h5b02;
        src5 <= 16'h1ec8;
        src6 <= 16'h70d8;
        src7 <= 16'ha4ef;
        src8 <= 16'haaab;
        src9 <= 16'had4e;
        src10 <= 16'he75a;
        src11 <= 16'hcb67;
        src12 <= 16'h27d0;
        src13 <= 16'h715f;
        src14 <= 16'hc0e6;
        src15 <= 16'hf1f7;
        src16 <= 16'h21de;
        src17 <= 16'h34a8;
        src18 <= 16'h8576;
        src19 <= 16'h54b9;
        src20 <= 16'hdd0b;
        src21 <= 16'h3558;
        src22 <= 16'h9059;
        src23 <= 16'h970b;
        src24 <= 16'h47df;
        src25 <= 16'h7b1c;
        src26 <= 16'h8b7f;
        src27 <= 16'he98a;
        src28 <= 16'he3c3;
        src29 <= 16'h5593;
        src30 <= 16'hd1d9;
        src31 <= 16'h6b2d;
        src32 <= 16'h8c73;
        src33 <= 16'haece;
        src34 <= 16'h3fee;
        src35 <= 16'hc3e8;
        src36 <= 16'h4806;
        src37 <= 16'hb4a6;
        src38 <= 16'he1a;
        src39 <= 16'hef92;
        src40 <= 16'habf0;
        src41 <= 16'hd667;
        src42 <= 16'h650a;
        src43 <= 16'h5005;
        src44 <= 16'ha0f9;
        src45 <= 16'h9fc5;
        src46 <= 16'hb5f9;
        src47 <= 16'h67a;
        src48 <= 16'he9c4;
        src49 <= 16'h868;
        src50 <= 16'h93e6;
        src51 <= 16'hd2e8;
        src52 <= 16'h2219;
        src53 <= 16'h7e82;
        src54 <= 16'h7625;
        src55 <= 16'hfab6;
        src56 <= 16'hf8cc;
        src57 <= 16'h6be7;
        src58 <= 16'h6af;
        src59 <= 16'h9a7b;
        src60 <= 16'hb1a9;
        src61 <= 16'h6da8;
        src62 <= 16'hf087;
        src63 <= 16'h8ce6;
        src64 <= 16'hf07d;
        src65 <= 16'h96e5;
        src66 <= 16'h604c;
        src67 <= 16'he4a9;
        src68 <= 16'h5e61;
        src69 <= 16'h28f7;
        src70 <= 16'h9f33;
        src71 <= 16'h5cab;
        src72 <= 16'h16c3;
        src73 <= 16'h7fa5;
        src74 <= 16'h349;
        src75 <= 16'h5783;
        src76 <= 16'haa5;
        src77 <= 16'hc5f4;
        src78 <= 16'h7dff;
        src79 <= 16'h6513;
        src80 <= 16'hc843;
        src81 <= 16'he6fa;
        src82 <= 16'h2588;
        src83 <= 16'ha3d9;
        src84 <= 16'hc052;
        src85 <= 16'had6b;
        src86 <= 16'hacab;
        src87 <= 16'h5c1b;
        src88 <= 16'hce6a;
        src89 <= 16'h439d;
        src90 <= 16'hf11c;
        src91 <= 16'ha462;
        src92 <= 16'h96f9;
        src93 <= 16'hbf10;
        src94 <= 16'ha6a9;
        src95 <= 16'h3342;
        src96 <= 16'hf19;
        src97 <= 16'h6012;
        src98 <= 16'hca50;
        src99 <= 16'h623f;
        src100 <= 16'h92c1;
        src101 <= 16'h784f;
        src102 <= 16'h3c44;
        src103 <= 16'h6aa5;
        src104 <= 16'h77e4;
        src105 <= 16'h49f7;
        src106 <= 16'ha0e4;
        src107 <= 16'h6a57;
        src108 <= 16'h602f;
        src109 <= 16'h7920;
        src110 <= 16'h4db;
        src111 <= 16'hd435;
        src112 <= 16'h6161;
        src113 <= 16'h10f0;
        src114 <= 16'h3825;
        src115 <= 16'hed51;
        src116 <= 16'h1d43;
        src117 <= 16'ha1ce;
        src118 <= 16'h9632;
        src119 <= 16'h1212;
        src120 <= 16'h7d3d;
        src121 <= 16'ha2a6;
        src122 <= 16'h55c0;
        src123 <= 16'h9509;
        src124 <= 16'h3f38;
        src125 <= 16'hbba3;
        src126 <= 16'h41b0;
        src127 <= 16'hb75e;
        src128 <= 16'hdb24;
        src129 <= 16'hab98;
        src130 <= 16'hfcf3;
        src131 <= 16'ha3f9;
        src132 <= 16'h9c4b;
        src133 <= 16'h3d39;
        src134 <= 16'hc7c8;
        src135 <= 16'h8502;
        src136 <= 16'hae37;
        src137 <= 16'h4aae;
        src138 <= 16'h5ee4;
        src139 <= 16'h750;
        src140 <= 16'h86ca;
        src141 <= 16'h1407;
        src142 <= 16'hdbd5;
        src143 <= 16'hc0fe;
        src144 <= 16'h88e3;
        src145 <= 16'h8456;
        src146 <= 16'h616e;
        src147 <= 16'h606d;
        src148 <= 16'hbe53;
        src149 <= 16'h8725;
        src150 <= 16'h83e3;
        src151 <= 16'h7c05;
        src152 <= 16'h20ef;
        src153 <= 16'h5325;
        src154 <= 16'hf208;
        src155 <= 16'hecb4;
        src156 <= 16'ha2ea;
        src157 <= 16'h5ce8;
        src158 <= 16'h4f96;
        src159 <= 16'h22e1;
        src160 <= 16'hb71b;
        src161 <= 16'h5760;
        exp <= 24'h51fd51;
        #1
        src0 <= 16'h8a45;
        src1 <= 16'hed61;
        src2 <= 16'h71dd;
        src3 <= 16'h6f8f;
        src4 <= 16'hb97c;
        src5 <= 16'h2dc5;
        src6 <= 16'h7506;
        src7 <= 16'h37ae;
        src8 <= 16'h1819;
        src9 <= 16'h6a0c;
        src10 <= 16'h809e;
        src11 <= 16'h183d;
        src12 <= 16'h5004;
        src13 <= 16'h1302;
        src14 <= 16'h1cf3;
        src15 <= 16'hdb9d;
        src16 <= 16'h4bbc;
        src17 <= 16'h8a75;
        src18 <= 16'h8b6a;
        src19 <= 16'h9a3;
        src20 <= 16'h9c6a;
        src21 <= 16'hf6a3;
        src22 <= 16'ha5f3;
        src23 <= 16'he91d;
        src24 <= 16'h2093;
        src25 <= 16'h6449;
        src26 <= 16'h25d;
        src27 <= 16'hc27b;
        src28 <= 16'ha666;
        src29 <= 16'h642a;
        src30 <= 16'h8a5d;
        src31 <= 16'hc41c;
        src32 <= 16'ha189;
        src33 <= 16'h3c12;
        src34 <= 16'hedeb;
        src35 <= 16'h7249;
        src36 <= 16'hb4e8;
        src37 <= 16'hf826;
        src38 <= 16'hd4d6;
        src39 <= 16'h38aa;
        src40 <= 16'h79ae;
        src41 <= 16'h8b4d;
        src42 <= 16'h7dbd;
        src43 <= 16'h4606;
        src44 <= 16'h3385;
        src45 <= 16'h2d49;
        src46 <= 16'h6d20;
        src47 <= 16'h8b2b;
        src48 <= 16'h255;
        src49 <= 16'h2ce5;
        src50 <= 16'hf329;
        src51 <= 16'h991d;
        src52 <= 16'he498;
        src53 <= 16'hfbc;
        src54 <= 16'h4fd5;
        src55 <= 16'h9fda;
        src56 <= 16'h593f;
        src57 <= 16'h650a;
        src58 <= 16'haa4c;
        src59 <= 16'h7e7f;
        src60 <= 16'h5002;
        src61 <= 16'h711c;
        src62 <= 16'h7b95;
        src63 <= 16'hc211;
        src64 <= 16'h3844;
        src65 <= 16'h9c5a;
        src66 <= 16'h4849;
        src67 <= 16'hb9d4;
        src68 <= 16'hb828;
        src69 <= 16'hc675;
        src70 <= 16'h98d6;
        src71 <= 16'hedfb;
        src72 <= 16'h60f0;
        src73 <= 16'h257;
        src74 <= 16'h61e;
        src75 <= 16'h4fe7;
        src76 <= 16'hcca7;
        src77 <= 16'hce03;
        src78 <= 16'hc92c;
        src79 <= 16'h8861;
        src80 <= 16'head0;
        src81 <= 16'h7402;
        src82 <= 16'hc628;
        src83 <= 16'h9a60;
        src84 <= 16'ha6d6;
        src85 <= 16'h5a1a;
        src86 <= 16'h9ca8;
        src87 <= 16'h5642;
        src88 <= 16'hb9e7;
        src89 <= 16'hf326;
        src90 <= 16'he7f1;
        src91 <= 16'h25ab;
        src92 <= 16'hb083;
        src93 <= 16'hc0b7;
        src94 <= 16'hf34f;
        src95 <= 16'h67fb;
        src96 <= 16'hd9b1;
        src97 <= 16'hccf1;
        src98 <= 16'h3566;
        src99 <= 16'h13b;
        src100 <= 16'hab59;
        src101 <= 16'h440c;
        src102 <= 16'h332d;
        src103 <= 16'he26a;
        src104 <= 16'h30aa;
        src105 <= 16'ha86f;
        src106 <= 16'hb439;
        src107 <= 16'h2d92;
        src108 <= 16'hffd7;
        src109 <= 16'h28b;
        src110 <= 16'h4809;
        src111 <= 16'hcd6a;
        src112 <= 16'hd199;
        src113 <= 16'h5092;
        src114 <= 16'hc4ff;
        src115 <= 16'hbe17;
        src116 <= 16'h1d6a;
        src117 <= 16'h45f4;
        src118 <= 16'hb025;
        src119 <= 16'h4f43;
        src120 <= 16'hec32;
        src121 <= 16'hc43a;
        src122 <= 16'h2603;
        src123 <= 16'hf1ef;
        src124 <= 16'he71f;
        src125 <= 16'h4bca;
        src126 <= 16'h3aea;
        src127 <= 16'h1886;
        src128 <= 16'hfb59;
        src129 <= 16'h82ec;
        src130 <= 16'h1cb4;
        src131 <= 16'ha104;
        src132 <= 16'h149d;
        src133 <= 16'h84e;
        src134 <= 16'h508f;
        src135 <= 16'hd4c0;
        src136 <= 16'h6fa5;
        src137 <= 16'ha8b5;
        src138 <= 16'ha566;
        src139 <= 16'ha40;
        src140 <= 16'h6c74;
        src141 <= 16'h6466;
        src142 <= 16'h8db2;
        src143 <= 16'h4c8c;
        src144 <= 16'h7f92;
        src145 <= 16'hd952;
        src146 <= 16'h5b1d;
        src147 <= 16'he220;
        src148 <= 16'h8d9d;
        src149 <= 16'hfbfc;
        src150 <= 16'h60e5;
        src151 <= 16'h7819;
        src152 <= 16'h8476;
        src153 <= 16'h5088;
        src154 <= 16'hdf8f;
        src155 <= 16'h5572;
        src156 <= 16'h49f8;
        src157 <= 16'hd71c;
        src158 <= 16'h8f6d;
        src159 <= 16'hbfa8;
        src160 <= 16'h48f7;
        src161 <= 16'h439f;
        exp <= 24'h51ebcc;
        #1
        src0 <= 16'ha31b;
        src1 <= 16'hd6b6;
        src2 <= 16'h95b8;
        src3 <= 16'ha331;
        src4 <= 16'h2184;
        src5 <= 16'h84a3;
        src6 <= 16'hace3;
        src7 <= 16'h2228;
        src8 <= 16'h9f1;
        src9 <= 16'hc328;
        src10 <= 16'h661d;
        src11 <= 16'hcb87;
        src12 <= 16'hbf4f;
        src13 <= 16'h5e6;
        src14 <= 16'h847a;
        src15 <= 16'hd864;
        src16 <= 16'h8310;
        src17 <= 16'he765;
        src18 <= 16'h5ae2;
        src19 <= 16'hc7ab;
        src20 <= 16'h742;
        src21 <= 16'h1569;
        src22 <= 16'h5323;
        src23 <= 16'h256d;
        src24 <= 16'hb54;
        src25 <= 16'hd9df;
        src26 <= 16'ha7b6;
        src27 <= 16'hc7e5;
        src28 <= 16'hb882;
        src29 <= 16'h5fe0;
        src30 <= 16'hdb49;
        src31 <= 16'h5024;
        src32 <= 16'h34e1;
        src33 <= 16'he7c7;
        src34 <= 16'h2b55;
        src35 <= 16'h2f2e;
        src36 <= 16'h1bd3;
        src37 <= 16'h9e27;
        src38 <= 16'ha776;
        src39 <= 16'hbf76;
        src40 <= 16'hbadb;
        src41 <= 16'h365c;
        src42 <= 16'hfac0;
        src43 <= 16'heff7;
        src44 <= 16'h5cd8;
        src45 <= 16'hbccf;
        src46 <= 16'h73ea;
        src47 <= 16'hf216;
        src48 <= 16'haa5f;
        src49 <= 16'haebf;
        src50 <= 16'h578;
        src51 <= 16'h7217;
        src52 <= 16'h7fd0;
        src53 <= 16'ha737;
        src54 <= 16'h6c59;
        src55 <= 16'hc269;
        src56 <= 16'h348;
        src57 <= 16'h54c0;
        src58 <= 16'h432f;
        src59 <= 16'hfb8f;
        src60 <= 16'hd146;
        src61 <= 16'h56fc;
        src62 <= 16'h7b02;
        src63 <= 16'h22bd;
        src64 <= 16'ha176;
        src65 <= 16'h5a01;
        src66 <= 16'hcb96;
        src67 <= 16'hba8a;
        src68 <= 16'h50a1;
        src69 <= 16'h92f8;
        src70 <= 16'hc276;
        src71 <= 16'hbca0;
        src72 <= 16'h656f;
        src73 <= 16'he0b9;
        src74 <= 16'h47b9;
        src75 <= 16'h3143;
        src76 <= 16'h1e0b;
        src77 <= 16'hdb66;
        src78 <= 16'h52a9;
        src79 <= 16'hc92f;
        src80 <= 16'heb4b;
        src81 <= 16'h683;
        src82 <= 16'h496e;
        src83 <= 16'he8b3;
        src84 <= 16'h2205;
        src85 <= 16'ha2e0;
        src86 <= 16'h9c4a;
        src87 <= 16'h7ef7;
        src88 <= 16'h9edc;
        src89 <= 16'h65dc;
        src90 <= 16'hc05e;
        src91 <= 16'h1990;
        src92 <= 16'h36eb;
        src93 <= 16'h4695;
        src94 <= 16'h4a0f;
        src95 <= 16'hfc52;
        src96 <= 16'h56a5;
        src97 <= 16'hb42c;
        src98 <= 16'h1299;
        src99 <= 16'h9b63;
        src100 <= 16'hc5f4;
        src101 <= 16'hfdf7;
        src102 <= 16'h37e0;
        src103 <= 16'h7fd9;
        src104 <= 16'hd432;
        src105 <= 16'he5aa;
        src106 <= 16'h70fc;
        src107 <= 16'h85bb;
        src108 <= 16'ha700;
        src109 <= 16'ha80e;
        src110 <= 16'h7be8;
        src111 <= 16'h920b;
        src112 <= 16'hc41f;
        src113 <= 16'h9b16;
        src114 <= 16'he633;
        src115 <= 16'hfaa3;
        src116 <= 16'hfec2;
        src117 <= 16'h2dc9;
        src118 <= 16'h442b;
        src119 <= 16'h57ae;
        src120 <= 16'h3254;
        src121 <= 16'h41af;
        src122 <= 16'hdfc5;
        src123 <= 16'hb17d;
        src124 <= 16'he892;
        src125 <= 16'hc094;
        src126 <= 16'hc135;
        src127 <= 16'h13c;
        src128 <= 16'h364d;
        src129 <= 16'h9f09;
        src130 <= 16'h82d7;
        src131 <= 16'h256f;
        src132 <= 16'h7853;
        src133 <= 16'h9cf2;
        src134 <= 16'h4e1;
        src135 <= 16'hff67;
        src136 <= 16'h2b97;
        src137 <= 16'h5b5a;
        src138 <= 16'h29cd;
        src139 <= 16'h8f4d;
        src140 <= 16'h4d51;
        src141 <= 16'hbae8;
        src142 <= 16'hd506;
        src143 <= 16'h8828;
        src144 <= 16'hb017;
        src145 <= 16'h99d1;
        src146 <= 16'h1565;
        src147 <= 16'hf840;
        src148 <= 16'h8f85;
        src149 <= 16'hf974;
        src150 <= 16'h9b41;
        src151 <= 16'h389b;
        src152 <= 16'hc97e;
        src153 <= 16'h8f3f;
        src154 <= 16'h8adf;
        src155 <= 16'h2a70;
        src156 <= 16'h1670;
        src157 <= 16'h7f22;
        src158 <= 16'h5fba;
        src159 <= 16'h184e;
        src160 <= 16'hbf16;
        src161 <= 16'h67e7;
        exp <= 24'h53c8b8;
        #1
        src0 <= 16'hb8d4;
        src1 <= 16'h2dff;
        src2 <= 16'h6826;
        src3 <= 16'hd0c2;
        src4 <= 16'heb89;
        src5 <= 16'h6034;
        src6 <= 16'h4eba;
        src7 <= 16'hdb00;
        src8 <= 16'h8c50;
        src9 <= 16'h4c7a;
        src10 <= 16'hdea0;
        src11 <= 16'h8a21;
        src12 <= 16'h84e8;
        src13 <= 16'h4c3e;
        src14 <= 16'h8a35;
        src15 <= 16'hb33;
        src16 <= 16'h1a8a;
        src17 <= 16'hf754;
        src18 <= 16'ha87c;
        src19 <= 16'hb9b1;
        src20 <= 16'h415c;
        src21 <= 16'h3c41;
        src22 <= 16'h4cf9;
        src23 <= 16'hc628;
        src24 <= 16'ha7c;
        src25 <= 16'he71c;
        src26 <= 16'h67a7;
        src27 <= 16'h87a;
        src28 <= 16'h61b6;
        src29 <= 16'h6cbc;
        src30 <= 16'h18;
        src31 <= 16'h802c;
        src32 <= 16'ha3ee;
        src33 <= 16'hf1c4;
        src34 <= 16'h1e10;
        src35 <= 16'hda76;
        src36 <= 16'hbdf1;
        src37 <= 16'h7f37;
        src38 <= 16'ha0a4;
        src39 <= 16'hb9d1;
        src40 <= 16'h1911;
        src41 <= 16'h131e;
        src42 <= 16'h7fd2;
        src43 <= 16'hf7f3;
        src44 <= 16'h23a6;
        src45 <= 16'h244b;
        src46 <= 16'h4dce;
        src47 <= 16'h6488;
        src48 <= 16'h3351;
        src49 <= 16'h27da;
        src50 <= 16'h6f62;
        src51 <= 16'he26c;
        src52 <= 16'hc303;
        src53 <= 16'hb297;
        src54 <= 16'h1536;
        src55 <= 16'hb7fb;
        src56 <= 16'h357a;
        src57 <= 16'h2f30;
        src58 <= 16'h3694;
        src59 <= 16'h2567;
        src60 <= 16'hcd1e;
        src61 <= 16'hfc93;
        src62 <= 16'hff3d;
        src63 <= 16'h113;
        src64 <= 16'h512a;
        src65 <= 16'hb11d;
        src66 <= 16'ha719;
        src67 <= 16'h31c;
        src68 <= 16'hf48f;
        src69 <= 16'h5128;
        src70 <= 16'h7283;
        src71 <= 16'h721e;
        src72 <= 16'h127e;
        src73 <= 16'h7446;
        src74 <= 16'h834;
        src75 <= 16'hb248;
        src76 <= 16'ha39d;
        src77 <= 16'hf800;
        src78 <= 16'h69af;
        src79 <= 16'hf32d;
        src80 <= 16'hbe69;
        src81 <= 16'h564c;
        src82 <= 16'hc17b;
        src83 <= 16'ha17;
        src84 <= 16'h8762;
        src85 <= 16'ha218;
        src86 <= 16'hddb5;
        src87 <= 16'h481e;
        src88 <= 16'h6a3d;
        src89 <= 16'h5f0e;
        src90 <= 16'h62bc;
        src91 <= 16'h710c;
        src92 <= 16'hca0c;
        src93 <= 16'h1b05;
        src94 <= 16'hdbb8;
        src95 <= 16'h31a9;
        src96 <= 16'ha802;
        src97 <= 16'h54f;
        src98 <= 16'hea34;
        src99 <= 16'h30e0;
        src100 <= 16'h370d;
        src101 <= 16'h5213;
        src102 <= 16'h3a6e;
        src103 <= 16'h60bc;
        src104 <= 16'h7dd5;
        src105 <= 16'h39d9;
        src106 <= 16'h648c;
        src107 <= 16'h568d;
        src108 <= 16'h6cff;
        src109 <= 16'h4bb9;
        src110 <= 16'hf58a;
        src111 <= 16'h29cf;
        src112 <= 16'h2a3;
        src113 <= 16'h7c5;
        src114 <= 16'hc1b2;
        src115 <= 16'h5cff;
        src116 <= 16'h5521;
        src117 <= 16'h2c62;
        src118 <= 16'h25aa;
        src119 <= 16'hb1eb;
        src120 <= 16'h2766;
        src121 <= 16'h8e60;
        src122 <= 16'h8b20;
        src123 <= 16'hcae3;
        src124 <= 16'hc4ad;
        src125 <= 16'h66cd;
        src126 <= 16'hc7fb;
        src127 <= 16'h8410;
        src128 <= 16'h1dd4;
        src129 <= 16'hb055;
        src130 <= 16'hf7b7;
        src131 <= 16'h8d36;
        src132 <= 16'h4150;
        src133 <= 16'h6d1;
        src134 <= 16'h1cea;
        src135 <= 16'ha758;
        src136 <= 16'h74ed;
        src137 <= 16'h5125;
        src138 <= 16'h22c5;
        src139 <= 16'he505;
        src140 <= 16'hf93c;
        src141 <= 16'ha9a;
        src142 <= 16'hc20f;
        src143 <= 16'h401b;
        src144 <= 16'h7d71;
        src145 <= 16'heb45;
        src146 <= 16'h5996;
        src147 <= 16'h5cb4;
        src148 <= 16'ha8c7;
        src149 <= 16'hcfd8;
        src150 <= 16'h4b4e;
        src151 <= 16'h837;
        src152 <= 16'h793;
        src153 <= 16'h31e3;
        src154 <= 16'he28e;
        src155 <= 16'h990a;
        src156 <= 16'h8321;
        src157 <= 16'h8c54;
        src158 <= 16'h57fb;
        src159 <= 16'h4cd0;
        src160 <= 16'hbc2d;
        src161 <= 16'h4178;
        exp <= 24'h4ac315;
        #1
        src0 <= 16'h3d58;
        src1 <= 16'he790;
        src2 <= 16'h565b;
        src3 <= 16'h4b2d;
        src4 <= 16'h70f3;
        src5 <= 16'h1124;
        src6 <= 16'hcf4d;
        src7 <= 16'h1254;
        src8 <= 16'hf08e;
        src9 <= 16'hc0dd;
        src10 <= 16'hf985;
        src11 <= 16'hbb62;
        src12 <= 16'h4594;
        src13 <= 16'hc64e;
        src14 <= 16'h3ec0;
        src15 <= 16'hf595;
        src16 <= 16'h5f8d;
        src17 <= 16'hee64;
        src18 <= 16'h729d;
        src19 <= 16'hb7a6;
        src20 <= 16'h79af;
        src21 <= 16'hdc99;
        src22 <= 16'h91b2;
        src23 <= 16'hed40;
        src24 <= 16'hc33e;
        src25 <= 16'haef4;
        src26 <= 16'h7dfd;
        src27 <= 16'h2b95;
        src28 <= 16'h22c3;
        src29 <= 16'h8950;
        src30 <= 16'he89b;
        src31 <= 16'heed8;
        src32 <= 16'hb2b4;
        src33 <= 16'hc884;
        src34 <= 16'heccb;
        src35 <= 16'h81ce;
        src36 <= 16'h563c;
        src37 <= 16'h4742;
        src38 <= 16'h1444;
        src39 <= 16'he628;
        src40 <= 16'h15b;
        src41 <= 16'hdfe7;
        src42 <= 16'hb9c2;
        src43 <= 16'h85b0;
        src44 <= 16'h7e29;
        src45 <= 16'hc500;
        src46 <= 16'h1510;
        src47 <= 16'hface;
        src48 <= 16'hc32;
        src49 <= 16'h304a;
        src50 <= 16'h140c;
        src51 <= 16'he3ca;
        src52 <= 16'h160a;
        src53 <= 16'hd875;
        src54 <= 16'hcc10;
        src55 <= 16'h8709;
        src56 <= 16'hfa1f;
        src57 <= 16'h7849;
        src58 <= 16'hd614;
        src59 <= 16'h8f3;
        src60 <= 16'hf587;
        src61 <= 16'h91c9;
        src62 <= 16'hf702;
        src63 <= 16'h994;
        src64 <= 16'h1771;
        src65 <= 16'h5c45;
        src66 <= 16'h75c6;
        src67 <= 16'h156f;
        src68 <= 16'h19f9;
        src69 <= 16'h5cef;
        src70 <= 16'h148c;
        src71 <= 16'h5a82;
        src72 <= 16'he7df;
        src73 <= 16'h8f18;
        src74 <= 16'hcb40;
        src75 <= 16'h90d6;
        src76 <= 16'h736c;
        src77 <= 16'h760a;
        src78 <= 16'h66c5;
        src79 <= 16'h3503;
        src80 <= 16'h5d9f;
        src81 <= 16'h34cb;
        src82 <= 16'hcb5a;
        src83 <= 16'hd9f6;
        src84 <= 16'hfd46;
        src85 <= 16'h4e59;
        src86 <= 16'h8435;
        src87 <= 16'h1d3e;
        src88 <= 16'hc4e8;
        src89 <= 16'h1415;
        src90 <= 16'h3eea;
        src91 <= 16'h8be7;
        src92 <= 16'h76b3;
        src93 <= 16'h34a;
        src94 <= 16'h71c6;
        src95 <= 16'h60c6;
        src96 <= 16'h4a49;
        src97 <= 16'he57;
        src98 <= 16'h5ffe;
        src99 <= 16'hbe4c;
        src100 <= 16'hee10;
        src101 <= 16'h2a7f;
        src102 <= 16'hb22e;
        src103 <= 16'h7e12;
        src104 <= 16'h8064;
        src105 <= 16'ha5f5;
        src106 <= 16'h792c;
        src107 <= 16'h4a27;
        src108 <= 16'hd566;
        src109 <= 16'h4f8e;
        src110 <= 16'h2902;
        src111 <= 16'hb741;
        src112 <= 16'h5ba;
        src113 <= 16'h5fc5;
        src114 <= 16'hb6d3;
        src115 <= 16'h29f4;
        src116 <= 16'h9dcd;
        src117 <= 16'h1b11;
        src118 <= 16'h5ec1;
        src119 <= 16'hc96c;
        src120 <= 16'ha983;
        src121 <= 16'hebe5;
        src122 <= 16'ha157;
        src123 <= 16'h17d2;
        src124 <= 16'hc951;
        src125 <= 16'he500;
        src126 <= 16'h87ed;
        src127 <= 16'h9da8;
        src128 <= 16'he17b;
        src129 <= 16'h4b7;
        src130 <= 16'hcae4;
        src131 <= 16'h4d06;
        src132 <= 16'hf9a8;
        src133 <= 16'h8223;
        src134 <= 16'had23;
        src135 <= 16'hf026;
        src136 <= 16'h543b;
        src137 <= 16'hd585;
        src138 <= 16'h1c1f;
        src139 <= 16'h15dd;
        src140 <= 16'hef69;
        src141 <= 16'hc680;
        src142 <= 16'hda14;
        src143 <= 16'hb97b;
        src144 <= 16'hb258;
        src145 <= 16'h5270;
        src146 <= 16'h8bf9;
        src147 <= 16'hff38;
        src148 <= 16'h89e0;
        src149 <= 16'h4c35;
        src150 <= 16'hffd7;
        src151 <= 16'hd35e;
        src152 <= 16'h7095;
        src153 <= 16'h4f13;
        src154 <= 16'hcce5;
        src155 <= 16'h4f90;
        src156 <= 16'haac0;
        src157 <= 16'hd226;
        src158 <= 16'h7949;
        src159 <= 16'ha007;
        src160 <= 16'h3149;
        src161 <= 16'h2175;
        exp <= 24'h550789;
        #1
        src0 <= 16'h82ca;
        src1 <= 16'h7ed;
        src2 <= 16'hf367;
        src3 <= 16'hdbd8;
        src4 <= 16'hb30d;
        src5 <= 16'hdee8;
        src6 <= 16'h6c62;
        src7 <= 16'h4fd4;
        src8 <= 16'h21c;
        src9 <= 16'h17db;
        src10 <= 16'ha4d6;
        src11 <= 16'heee;
        src12 <= 16'hd2d3;
        src13 <= 16'hdec4;
        src14 <= 16'h58e2;
        src15 <= 16'hdbec;
        src16 <= 16'h6419;
        src17 <= 16'h6e36;
        src18 <= 16'h83b1;
        src19 <= 16'h4814;
        src20 <= 16'hc2c8;
        src21 <= 16'h2abc;
        src22 <= 16'h8a13;
        src23 <= 16'hb8a5;
        src24 <= 16'hc58a;
        src25 <= 16'ha7f;
        src26 <= 16'hb0d5;
        src27 <= 16'h1dfa;
        src28 <= 16'h848f;
        src29 <= 16'h4a28;
        src30 <= 16'hd36b;
        src31 <= 16'hc671;
        src32 <= 16'h1b15;
        src33 <= 16'h6ee;
        src34 <= 16'hc2bb;
        src35 <= 16'he8da;
        src36 <= 16'hf5dc;
        src37 <= 16'ha6dc;
        src38 <= 16'hf8b7;
        src39 <= 16'h5187;
        src40 <= 16'ha908;
        src41 <= 16'hd080;
        src42 <= 16'h4560;
        src43 <= 16'h71ba;
        src44 <= 16'h8bbf;
        src45 <= 16'h9383;
        src46 <= 16'h26a0;
        src47 <= 16'h1f32;
        src48 <= 16'h1500;
        src49 <= 16'hb58c;
        src50 <= 16'h7a37;
        src51 <= 16'h101e;
        src52 <= 16'h5b5b;
        src53 <= 16'h84b2;
        src54 <= 16'hdb1;
        src55 <= 16'hb1b2;
        src56 <= 16'h9e49;
        src57 <= 16'h26a5;
        src58 <= 16'hb73e;
        src59 <= 16'h67c6;
        src60 <= 16'hccd0;
        src61 <= 16'h5e6c;
        src62 <= 16'h71b0;
        src63 <= 16'hd9a3;
        src64 <= 16'hdeed;
        src65 <= 16'h9bd4;
        src66 <= 16'h75e1;
        src67 <= 16'h5b60;
        src68 <= 16'hf18f;
        src69 <= 16'h1467;
        src70 <= 16'h8010;
        src71 <= 16'h3c3b;
        src72 <= 16'h3a06;
        src73 <= 16'h6bf0;
        src74 <= 16'hf6da;
        src75 <= 16'h73f7;
        src76 <= 16'hafdc;
        src77 <= 16'h8d14;
        src78 <= 16'h13eb;
        src79 <= 16'hcabd;
        src80 <= 16'hc3fe;
        src81 <= 16'hecc6;
        src82 <= 16'h9339;
        src83 <= 16'h883;
        src84 <= 16'h5ee6;
        src85 <= 16'hf7b2;
        src86 <= 16'h3ab2;
        src87 <= 16'hb88f;
        src88 <= 16'h692d;
        src89 <= 16'ha1d9;
        src90 <= 16'h6e2e;
        src91 <= 16'hc9be;
        src92 <= 16'h4192;
        src93 <= 16'hcdb4;
        src94 <= 16'h2d90;
        src95 <= 16'hd30d;
        src96 <= 16'h112b;
        src97 <= 16'h3a2b;
        src98 <= 16'h72a2;
        src99 <= 16'h6139;
        src100 <= 16'hb90f;
        src101 <= 16'hd5d0;
        src102 <= 16'hf2d8;
        src103 <= 16'h837d;
        src104 <= 16'h3d3e;
        src105 <= 16'had9d;
        src106 <= 16'h200b;
        src107 <= 16'h50c;
        src108 <= 16'h355f;
        src109 <= 16'h6cc8;
        src110 <= 16'h7e88;
        src111 <= 16'h5da8;
        src112 <= 16'hd117;
        src113 <= 16'h15c9;
        src114 <= 16'h6a71;
        src115 <= 16'h7ab0;
        src116 <= 16'h8a8a;
        src117 <= 16'h2c41;
        src118 <= 16'h88f7;
        src119 <= 16'h5ba2;
        src120 <= 16'h1013;
        src121 <= 16'hcac0;
        src122 <= 16'hf6f6;
        src123 <= 16'hee15;
        src124 <= 16'hdf86;
        src125 <= 16'he90f;
        src126 <= 16'h7a24;
        src127 <= 16'hc86e;
        src128 <= 16'hb069;
        src129 <= 16'hac61;
        src130 <= 16'hd842;
        src131 <= 16'h45f4;
        src132 <= 16'hb78d;
        src133 <= 16'h371e;
        src134 <= 16'heaa1;
        src135 <= 16'he982;
        src136 <= 16'hf84f;
        src137 <= 16'hfb82;
        src138 <= 16'hc4ce;
        src139 <= 16'h977c;
        src140 <= 16'h2c1d;
        src141 <= 16'he5d2;
        src142 <= 16'h2759;
        src143 <= 16'h82c4;
        src144 <= 16'h632e;
        src145 <= 16'heef2;
        src146 <= 16'hd9f2;
        src147 <= 16'h5008;
        src148 <= 16'he1bc;
        src149 <= 16'h5bd9;
        src150 <= 16'hedf7;
        src151 <= 16'he0f0;
        src152 <= 16'h1633;
        src153 <= 16'hd565;
        src154 <= 16'h1d85;
        src155 <= 16'hd186;
        src156 <= 16'hed89;
        src157 <= 16'h57cb;
        src158 <= 16'h32c;
        src159 <= 16'he6b1;
        src160 <= 16'h3ade;
        src161 <= 16'hfe78;
        exp <= 24'h55e9af;
        #1
        src0 <= 16'hba26;
        src1 <= 16'hd8d;
        src2 <= 16'h72a6;
        src3 <= 16'ha461;
        src4 <= 16'h397;
        src5 <= 16'he1c7;
        src6 <= 16'h85f3;
        src7 <= 16'h8a9d;
        src8 <= 16'hd2b0;
        src9 <= 16'h64e;
        src10 <= 16'hee7;
        src11 <= 16'ha871;
        src12 <= 16'ha930;
        src13 <= 16'h9115;
        src14 <= 16'h5e4f;
        src15 <= 16'hfab;
        src16 <= 16'h8d9e;
        src17 <= 16'h5f72;
        src18 <= 16'hef7d;
        src19 <= 16'h94db;
        src20 <= 16'h8696;
        src21 <= 16'h1418;
        src22 <= 16'h943b;
        src23 <= 16'hee87;
        src24 <= 16'hba6c;
        src25 <= 16'hec31;
        src26 <= 16'h6c6;
        src27 <= 16'h4ab1;
        src28 <= 16'h9c0;
        src29 <= 16'h787d;
        src30 <= 16'h79ad;
        src31 <= 16'hc4c1;
        src32 <= 16'h9157;
        src33 <= 16'h1483;
        src34 <= 16'h40fb;
        src35 <= 16'h3b7b;
        src36 <= 16'h3541;
        src37 <= 16'hfe90;
        src38 <= 16'h996b;
        src39 <= 16'h2e3d;
        src40 <= 16'hdb96;
        src41 <= 16'ha32e;
        src42 <= 16'ha900;
        src43 <= 16'h4056;
        src44 <= 16'he26e;
        src45 <= 16'h898f;
        src46 <= 16'h56de;
        src47 <= 16'ha05a;
        src48 <= 16'h88f3;
        src49 <= 16'h788e;
        src50 <= 16'h4f29;
        src51 <= 16'h2fb8;
        src52 <= 16'hcabc;
        src53 <= 16'h9b99;
        src54 <= 16'hec85;
        src55 <= 16'heef9;
        src56 <= 16'h136;
        src57 <= 16'h9206;
        src58 <= 16'h1b08;
        src59 <= 16'h3c80;
        src60 <= 16'h229f;
        src61 <= 16'hcb35;
        src62 <= 16'heba3;
        src63 <= 16'ha604;
        src64 <= 16'h5904;
        src65 <= 16'he314;
        src66 <= 16'hb777;
        src67 <= 16'hf9ca;
        src68 <= 16'hd8ea;
        src69 <= 16'h495a;
        src70 <= 16'he580;
        src71 <= 16'h3ca2;
        src72 <= 16'h638d;
        src73 <= 16'ha7cd;
        src74 <= 16'h31dd;
        src75 <= 16'he75c;
        src76 <= 16'h4b11;
        src77 <= 16'hd8f4;
        src78 <= 16'h489d;
        src79 <= 16'h5cfc;
        src80 <= 16'hed8d;
        src81 <= 16'ha1d9;
        src82 <= 16'h3d8c;
        src83 <= 16'he237;
        src84 <= 16'h14d9;
        src85 <= 16'h12ea;
        src86 <= 16'hde7a;
        src87 <= 16'hfb41;
        src88 <= 16'hbb3;
        src89 <= 16'hee92;
        src90 <= 16'hd00f;
        src91 <= 16'h6b5f;
        src92 <= 16'hee44;
        src93 <= 16'hff44;
        src94 <= 16'h1a63;
        src95 <= 16'h3933;
        src96 <= 16'h72f8;
        src97 <= 16'h7de4;
        src98 <= 16'h6bce;
        src99 <= 16'h75e2;
        src100 <= 16'hc2d6;
        src101 <= 16'h2537;
        src102 <= 16'h1da3;
        src103 <= 16'h81dc;
        src104 <= 16'h62ab;
        src105 <= 16'hfeaa;
        src106 <= 16'ha347;
        src107 <= 16'h8397;
        src108 <= 16'hf78c;
        src109 <= 16'haad0;
        src110 <= 16'h1552;
        src111 <= 16'h532f;
        src112 <= 16'h745a;
        src113 <= 16'h28b6;
        src114 <= 16'h7869;
        src115 <= 16'h26b2;
        src116 <= 16'h5e47;
        src117 <= 16'h5893;
        src118 <= 16'h5f1e;
        src119 <= 16'h7624;
        src120 <= 16'hade7;
        src121 <= 16'hec3a;
        src122 <= 16'he95d;
        src123 <= 16'h24fb;
        src124 <= 16'he9fe;
        src125 <= 16'h6181;
        src126 <= 16'h2029;
        src127 <= 16'hdcd5;
        src128 <= 16'h1fe;
        src129 <= 16'he163;
        src130 <= 16'h90ca;
        src131 <= 16'ha6fd;
        src132 <= 16'h4f62;
        src133 <= 16'hbd97;
        src134 <= 16'h8e04;
        src135 <= 16'h98f1;
        src136 <= 16'hc2fa;
        src137 <= 16'he7d3;
        src138 <= 16'h9bbe;
        src139 <= 16'he09c;
        src140 <= 16'he656;
        src141 <= 16'hd19e;
        src142 <= 16'hf3e5;
        src143 <= 16'h52b2;
        src144 <= 16'hbce;
        src145 <= 16'hd8a6;
        src146 <= 16'h4c6b;
        src147 <= 16'h2cde;
        src148 <= 16'h9290;
        src149 <= 16'heeb5;
        src150 <= 16'hf35d;
        src151 <= 16'h2ab8;
        src152 <= 16'h43b9;
        src153 <= 16'h7597;
        src154 <= 16'he6f0;
        src155 <= 16'hab99;
        src156 <= 16'hf833;
        src157 <= 16'hbbdb;
        src158 <= 16'h4a0b;
        src159 <= 16'hca16;
        src160 <= 16'h3c46;
        src161 <= 16'h37ba;
        exp <= 24'h555214;
        #1
        src0 <= 16'h6669;
        src1 <= 16'h4c81;
        src2 <= 16'haa19;
        src3 <= 16'h9e9a;
        src4 <= 16'hd24d;
        src5 <= 16'hf1c1;
        src6 <= 16'h3b82;
        src7 <= 16'h8c7d;
        src8 <= 16'h269c;
        src9 <= 16'h84f;
        src10 <= 16'hb750;
        src11 <= 16'ha400;
        src12 <= 16'hea6f;
        src13 <= 16'hd7c0;
        src14 <= 16'h6b42;
        src15 <= 16'ha90;
        src16 <= 16'h16f5;
        src17 <= 16'h38f1;
        src18 <= 16'h5ab1;
        src19 <= 16'hbbe4;
        src20 <= 16'h25bb;
        src21 <= 16'had1c;
        src22 <= 16'ha372;
        src23 <= 16'hf9eb;
        src24 <= 16'hfb7b;
        src25 <= 16'h3409;
        src26 <= 16'h734b;
        src27 <= 16'hfff8;
        src28 <= 16'hfc58;
        src29 <= 16'hd049;
        src30 <= 16'h3e04;
        src31 <= 16'h96cf;
        src32 <= 16'hf8e8;
        src33 <= 16'hf69b;
        src34 <= 16'h9058;
        src35 <= 16'h7b91;
        src36 <= 16'hf8b6;
        src37 <= 16'h7be3;
        src38 <= 16'h46b6;
        src39 <= 16'h19cf;
        src40 <= 16'h2446;
        src41 <= 16'he40c;
        src42 <= 16'h268e;
        src43 <= 16'h5c94;
        src44 <= 16'h4cdd;
        src45 <= 16'h3b8c;
        src46 <= 16'h94da;
        src47 <= 16'h95c4;
        src48 <= 16'h8be2;
        src49 <= 16'h21d1;
        src50 <= 16'h3f75;
        src51 <= 16'hbffb;
        src52 <= 16'h56c0;
        src53 <= 16'h9aaa;
        src54 <= 16'ha0ba;
        src55 <= 16'h9b45;
        src56 <= 16'hd81e;
        src57 <= 16'h9197;
        src58 <= 16'h8089;
        src59 <= 16'hb86a;
        src60 <= 16'hc375;
        src61 <= 16'h910b;
        src62 <= 16'hf5a7;
        src63 <= 16'hef6f;
        src64 <= 16'h4c43;
        src65 <= 16'h5018;
        src66 <= 16'h4132;
        src67 <= 16'h65bf;
        src68 <= 16'hc00a;
        src69 <= 16'h2a1a;
        src70 <= 16'hf4fc;
        src71 <= 16'h62a9;
        src72 <= 16'h49dc;
        src73 <= 16'hf6c8;
        src74 <= 16'h3d4;
        src75 <= 16'hd21f;
        src76 <= 16'hf15c;
        src77 <= 16'h8c8f;
        src78 <= 16'h63c4;
        src79 <= 16'h54f6;
        src80 <= 16'h4771;
        src81 <= 16'h8575;
        src82 <= 16'ha410;
        src83 <= 16'ha796;
        src84 <= 16'h5b38;
        src85 <= 16'h3ec4;
        src86 <= 16'h4588;
        src87 <= 16'h55f9;
        src88 <= 16'h7e00;
        src89 <= 16'h2f44;
        src90 <= 16'h9df3;
        src91 <= 16'h57bd;
        src92 <= 16'h5655;
        src93 <= 16'ha379;
        src94 <= 16'hc18a;
        src95 <= 16'hd18d;
        src96 <= 16'h80f3;
        src97 <= 16'hbc72;
        src98 <= 16'h3d56;
        src99 <= 16'hfbac;
        src100 <= 16'h62e0;
        src101 <= 16'hebbf;
        src102 <= 16'h400d;
        src103 <= 16'h9ed2;
        src104 <= 16'h81e9;
        src105 <= 16'hc2d;
        src106 <= 16'hdd5f;
        src107 <= 16'h2189;
        src108 <= 16'hcd00;
        src109 <= 16'h634a;
        src110 <= 16'h6c48;
        src111 <= 16'hff4b;
        src112 <= 16'h44c5;
        src113 <= 16'h1120;
        src114 <= 16'h40aa;
        src115 <= 16'hde87;
        src116 <= 16'hb7ae;
        src117 <= 16'h9372;
        src118 <= 16'h95fd;
        src119 <= 16'hb374;
        src120 <= 16'h4cbf;
        src121 <= 16'h12ad;
        src122 <= 16'h33ba;
        src123 <= 16'h48d9;
        src124 <= 16'hb04a;
        src125 <= 16'hfbed;
        src126 <= 16'haf03;
        src127 <= 16'h94b;
        src128 <= 16'h3cd4;
        src129 <= 16'hef58;
        src130 <= 16'hbbda;
        src131 <= 16'hbc79;
        src132 <= 16'h8153;
        src133 <= 16'h171d;
        src134 <= 16'h977d;
        src135 <= 16'h35ca;
        src136 <= 16'hc4c8;
        src137 <= 16'h276;
        src138 <= 16'h7cf7;
        src139 <= 16'h9db8;
        src140 <= 16'h75b5;
        src141 <= 16'h7198;
        src142 <= 16'h8cb;
        src143 <= 16'hd138;
        src144 <= 16'h4647;
        src145 <= 16'hcf28;
        src146 <= 16'h4df2;
        src147 <= 16'h9a1b;
        src148 <= 16'hdb5;
        src149 <= 16'h270f;
        src150 <= 16'h9d3b;
        src151 <= 16'hd1be;
        src152 <= 16'hb4c4;
        src153 <= 16'h99aa;
        src154 <= 16'h74a4;
        src155 <= 16'h4845;
        src156 <= 16'h47c5;
        src157 <= 16'h784a;
        src158 <= 16'h18e8;
        src159 <= 16'hb63d;
        src160 <= 16'hcda1;
        src161 <= 16'h591d;
        exp <= 24'h52a1b2;
        #1
        src0 <= 16'hc97f;
        src1 <= 16'h7101;
        src2 <= 16'h89f8;
        src3 <= 16'h1cbb;
        src4 <= 16'h66f0;
        src5 <= 16'hb356;
        src6 <= 16'he70c;
        src7 <= 16'h58c5;
        src8 <= 16'h81bf;
        src9 <= 16'ha404;
        src10 <= 16'hcb86;
        src11 <= 16'h5fe6;
        src12 <= 16'hdc7e;
        src13 <= 16'hfc9c;
        src14 <= 16'hbff0;
        src15 <= 16'h3855;
        src16 <= 16'hf2ba;
        src17 <= 16'h2c21;
        src18 <= 16'hcbb0;
        src19 <= 16'ha54e;
        src20 <= 16'hd7bb;
        src21 <= 16'hd4c7;
        src22 <= 16'h91af;
        src23 <= 16'hdc28;
        src24 <= 16'h89c3;
        src25 <= 16'h4a82;
        src26 <= 16'h32b2;
        src27 <= 16'hd9fd;
        src28 <= 16'h859e;
        src29 <= 16'h6616;
        src30 <= 16'hf1f9;
        src31 <= 16'h94fb;
        src32 <= 16'hc275;
        src33 <= 16'heeef;
        src34 <= 16'h352d;
        src35 <= 16'hc3fa;
        src36 <= 16'hd17e;
        src37 <= 16'he9ce;
        src38 <= 16'h2d95;
        src39 <= 16'hdf0f;
        src40 <= 16'h19fc;
        src41 <= 16'hd400;
        src42 <= 16'h1033;
        src43 <= 16'hc1e1;
        src44 <= 16'hf9d4;
        src45 <= 16'ha9fc;
        src46 <= 16'h9eb4;
        src47 <= 16'h4a3;
        src48 <= 16'h4684;
        src49 <= 16'hc4a4;
        src50 <= 16'hfc86;
        src51 <= 16'h129b;
        src52 <= 16'h8005;
        src53 <= 16'h9ef2;
        src54 <= 16'h7eb4;
        src55 <= 16'h4328;
        src56 <= 16'h9eca;
        src57 <= 16'h7bdd;
        src58 <= 16'hc672;
        src59 <= 16'h8741;
        src60 <= 16'hac48;
        src61 <= 16'hd90c;
        src62 <= 16'h5022;
        src63 <= 16'h7f06;
        src64 <= 16'h9f81;
        src65 <= 16'h46ff;
        src66 <= 16'had49;
        src67 <= 16'h69b6;
        src68 <= 16'hec8e;
        src69 <= 16'hacc4;
        src70 <= 16'h210b;
        src71 <= 16'hd10e;
        src72 <= 16'hf3c2;
        src73 <= 16'h9935;
        src74 <= 16'h19d7;
        src75 <= 16'h96a8;
        src76 <= 16'h2a73;
        src77 <= 16'hb178;
        src78 <= 16'hc9a7;
        src79 <= 16'h12ac;
        src80 <= 16'hf8d;
        src81 <= 16'hbbda;
        src82 <= 16'h7816;
        src83 <= 16'hd8d2;
        src84 <= 16'ha7e8;
        src85 <= 16'h7c5e;
        src86 <= 16'hc170;
        src87 <= 16'h7876;
        src88 <= 16'h778f;
        src89 <= 16'hf7a8;
        src90 <= 16'hf67;
        src91 <= 16'hacb6;
        src92 <= 16'hdb07;
        src93 <= 16'h7a66;
        src94 <= 16'h7df9;
        src95 <= 16'h1ede;
        src96 <= 16'hec37;
        src97 <= 16'h22a4;
        src98 <= 16'hc4d9;
        src99 <= 16'hf178;
        src100 <= 16'h6bd9;
        src101 <= 16'h7719;
        src102 <= 16'h93d3;
        src103 <= 16'h29c9;
        src104 <= 16'h5d05;
        src105 <= 16'h8dfa;
        src106 <= 16'h328f;
        src107 <= 16'h3abb;
        src108 <= 16'h189c;
        src109 <= 16'hfe6;
        src110 <= 16'hb128;
        src111 <= 16'hb383;
        src112 <= 16'h6b58;
        src113 <= 16'hce03;
        src114 <= 16'hecd0;
        src115 <= 16'hb5c4;
        src116 <= 16'h2b65;
        src117 <= 16'hd973;
        src118 <= 16'h982c;
        src119 <= 16'hd7e3;
        src120 <= 16'hc1b5;
        src121 <= 16'hb77c;
        src122 <= 16'he40b;
        src123 <= 16'hd72;
        src124 <= 16'h381a;
        src125 <= 16'h8cee;
        src126 <= 16'h3929;
        src127 <= 16'h8371;
        src128 <= 16'h7618;
        src129 <= 16'h885c;
        src130 <= 16'h4e6f;
        src131 <= 16'ha61c;
        src132 <= 16'hf8f6;
        src133 <= 16'he4e6;
        src134 <= 16'hd5ef;
        src135 <= 16'h9c5;
        src136 <= 16'h81dc;
        src137 <= 16'h2274;
        src138 <= 16'h8536;
        src139 <= 16'h71e6;
        src140 <= 16'hd93e;
        src141 <= 16'h7f8d;
        src142 <= 16'hb174;
        src143 <= 16'hff76;
        src144 <= 16'h1f54;
        src145 <= 16'h64a8;
        src146 <= 16'h6121;
        src147 <= 16'h9a4e;
        src148 <= 16'h4d74;
        src149 <= 16'h3e8d;
        src150 <= 16'hcfb5;
        src151 <= 16'h1da5;
        src152 <= 16'hba2;
        src153 <= 16'h28e7;
        src154 <= 16'h3b3e;
        src155 <= 16'hab44;
        src156 <= 16'h3580;
        src157 <= 16'h93a0;
        src158 <= 16'h35c7;
        src159 <= 16'h4462;
        src160 <= 16'h1c48;
        src161 <= 16'h3517;
        exp <= 24'h562a7a;
        #1
        src0 <= 16'h61be;
        src1 <= 16'h87e;
        src2 <= 16'he01a;
        src3 <= 16'h5083;
        src4 <= 16'h1123;
        src5 <= 16'hf9c4;
        src6 <= 16'h8fd2;
        src7 <= 16'hd273;
        src8 <= 16'h91e4;
        src9 <= 16'hbcac;
        src10 <= 16'h6c52;
        src11 <= 16'h5cf2;
        src12 <= 16'h3645;
        src13 <= 16'h813a;
        src14 <= 16'h190e;
        src15 <= 16'h1ae2;
        src16 <= 16'hc1da;
        src17 <= 16'h833b;
        src18 <= 16'h79ac;
        src19 <= 16'hc7ff;
        src20 <= 16'h539;
        src21 <= 16'h580;
        src22 <= 16'h5d6b;
        src23 <= 16'hfb5a;
        src24 <= 16'h8929;
        src25 <= 16'h7541;
        src26 <= 16'h5ab6;
        src27 <= 16'he537;
        src28 <= 16'ha0f1;
        src29 <= 16'hb395;
        src30 <= 16'h94d7;
        src31 <= 16'h8f2c;
        src32 <= 16'h2fdd;
        src33 <= 16'h87e2;
        src34 <= 16'hb3b5;
        src35 <= 16'hb43f;
        src36 <= 16'hdfc0;
        src37 <= 16'h4bd;
        src38 <= 16'h9f84;
        src39 <= 16'hffa4;
        src40 <= 16'h5fd4;
        src41 <= 16'h8fd0;
        src42 <= 16'h7e0f;
        src43 <= 16'h43c4;
        src44 <= 16'hfc1e;
        src45 <= 16'hba39;
        src46 <= 16'h169d;
        src47 <= 16'h6be;
        src48 <= 16'h4460;
        src49 <= 16'hdf58;
        src50 <= 16'h8de2;
        src51 <= 16'h5548;
        src52 <= 16'hd230;
        src53 <= 16'h82b0;
        src54 <= 16'h73fc;
        src55 <= 16'hb33d;
        src56 <= 16'h1db3;
        src57 <= 16'hd1de;
        src58 <= 16'h8ae4;
        src59 <= 16'h80fb;
        src60 <= 16'hb6c8;
        src61 <= 16'h856d;
        src62 <= 16'hb063;
        src63 <= 16'h61e8;
        src64 <= 16'h5754;
        src65 <= 16'h7bec;
        src66 <= 16'h863a;
        src67 <= 16'hc2dd;
        src68 <= 16'h50;
        src69 <= 16'heed4;
        src70 <= 16'hfac1;
        src71 <= 16'h74f8;
        src72 <= 16'hdb8a;
        src73 <= 16'hc039;
        src74 <= 16'hca28;
        src75 <= 16'h69f4;
        src76 <= 16'h7a3e;
        src77 <= 16'hbab;
        src78 <= 16'h602;
        src79 <= 16'h5f8c;
        src80 <= 16'hdbef;
        src81 <= 16'h3839;
        src82 <= 16'he4c5;
        src83 <= 16'hb1f8;
        src84 <= 16'hfa18;
        src85 <= 16'hd33b;
        src86 <= 16'hadd2;
        src87 <= 16'h4532;
        src88 <= 16'hc6e5;
        src89 <= 16'hc465;
        src90 <= 16'h532c;
        src91 <= 16'haacc;
        src92 <= 16'h52ba;
        src93 <= 16'habab;
        src94 <= 16'h86a;
        src95 <= 16'h9099;
        src96 <= 16'h79ee;
        src97 <= 16'h4c42;
        src98 <= 16'h2b00;
        src99 <= 16'h84b6;
        src100 <= 16'hadc4;
        src101 <= 16'h71f8;
        src102 <= 16'hc7d5;
        src103 <= 16'h1eb1;
        src104 <= 16'h5127;
        src105 <= 16'h1bfa;
        src106 <= 16'h2a6e;
        src107 <= 16'h799b;
        src108 <= 16'h14be;
        src109 <= 16'hdfec;
        src110 <= 16'he227;
        src111 <= 16'h78c6;
        src112 <= 16'hb2b4;
        src113 <= 16'h3c57;
        src114 <= 16'h673e;
        src115 <= 16'h9abe;
        src116 <= 16'h617e;
        src117 <= 16'h3fd3;
        src118 <= 16'hd205;
        src119 <= 16'he26b;
        src120 <= 16'h52fc;
        src121 <= 16'h4211;
        src122 <= 16'hb67a;
        src123 <= 16'h98e8;
        src124 <= 16'h2c90;
        src125 <= 16'h7d4d;
        src126 <= 16'hf993;
        src127 <= 16'he20d;
        src128 <= 16'h6f4a;
        src129 <= 16'hf892;
        src130 <= 16'hdeb2;
        src131 <= 16'hbf78;
        src132 <= 16'h68ba;
        src133 <= 16'h3220;
        src134 <= 16'h1bd0;
        src135 <= 16'h95f3;
        src136 <= 16'h9398;
        src137 <= 16'h4886;
        src138 <= 16'h10f0;
        src139 <= 16'h9d21;
        src140 <= 16'hfc3c;
        src141 <= 16'hbe6;
        src142 <= 16'h24a4;
        src143 <= 16'hdb55;
        src144 <= 16'h2d7a;
        src145 <= 16'h7f52;
        src146 <= 16'h2dec;
        src147 <= 16'h353f;
        src148 <= 16'h1498;
        src149 <= 16'h5892;
        src150 <= 16'hed84;
        src151 <= 16'h8f7f;
        src152 <= 16'hf127;
        src153 <= 16'hf02f;
        src154 <= 16'h6a01;
        src155 <= 16'h561;
        src156 <= 16'h3ab4;
        src157 <= 16'hf6b9;
        src158 <= 16'ha1a4;
        src159 <= 16'hc71d;
        src160 <= 16'h8e7a;
        src161 <= 16'hd928;
        exp <= 24'h532378;
        #1
        src0 <= 16'h9901;
        src1 <= 16'h9131;
        src2 <= 16'h147a;
        src3 <= 16'h1a1c;
        src4 <= 16'hca27;
        src5 <= 16'h3574;
        src6 <= 16'hdfe8;
        src7 <= 16'hdf78;
        src8 <= 16'h389a;
        src9 <= 16'h3b96;
        src10 <= 16'hffb;
        src11 <= 16'h5f02;
        src12 <= 16'hc982;
        src13 <= 16'h32b2;
        src14 <= 16'h7a0a;
        src15 <= 16'h784a;
        src16 <= 16'h5af6;
        src17 <= 16'h2d9;
        src18 <= 16'h691c;
        src19 <= 16'h60e6;
        src20 <= 16'h68d1;
        src21 <= 16'ha432;
        src22 <= 16'h8cea;
        src23 <= 16'he4d9;
        src24 <= 16'h6373;
        src25 <= 16'ha597;
        src26 <= 16'hdc56;
        src27 <= 16'h49f3;
        src28 <= 16'hf6c0;
        src29 <= 16'h96b0;
        src30 <= 16'hbdfe;
        src31 <= 16'h3a25;
        src32 <= 16'haaaa;
        src33 <= 16'h1097;
        src34 <= 16'h9259;
        src35 <= 16'h23ba;
        src36 <= 16'hd099;
        src37 <= 16'h7045;
        src38 <= 16'ha9cd;
        src39 <= 16'h8c4b;
        src40 <= 16'h9ecb;
        src41 <= 16'h8edc;
        src42 <= 16'h8643;
        src43 <= 16'hb50;
        src44 <= 16'h5554;
        src45 <= 16'hd8e0;
        src46 <= 16'h32a;
        src47 <= 16'h6bb6;
        src48 <= 16'h7ece;
        src49 <= 16'h5a28;
        src50 <= 16'h794e;
        src51 <= 16'h15a7;
        src52 <= 16'ha390;
        src53 <= 16'h6e;
        src54 <= 16'hb923;
        src55 <= 16'hd80c;
        src56 <= 16'h5f18;
        src57 <= 16'h26cd;
        src58 <= 16'hf3e3;
        src59 <= 16'h8bcc;
        src60 <= 16'hab85;
        src61 <= 16'ha7d3;
        src62 <= 16'ha214;
        src63 <= 16'h3b21;
        src64 <= 16'h6631;
        src65 <= 16'h6c80;
        src66 <= 16'hacbb;
        src67 <= 16'h66ea;
        src68 <= 16'h312b;
        src69 <= 16'h1a42;
        src70 <= 16'hda7b;
        src71 <= 16'h782b;
        src72 <= 16'h4458;
        src73 <= 16'hc3c8;
        src74 <= 16'hd2c1;
        src75 <= 16'hc73c;
        src76 <= 16'hf11c;
        src77 <= 16'h8293;
        src78 <= 16'haff5;
        src79 <= 16'h256a;
        src80 <= 16'hec17;
        src81 <= 16'h6a7e;
        src82 <= 16'hbd7c;
        src83 <= 16'h3898;
        src84 <= 16'h769c;
        src85 <= 16'h7bbb;
        src86 <= 16'h8685;
        src87 <= 16'h7ec9;
        src88 <= 16'heb6e;
        src89 <= 16'hffb6;
        src90 <= 16'h2ec4;
        src91 <= 16'h68f1;
        src92 <= 16'h3d12;
        src93 <= 16'hbaeb;
        src94 <= 16'h5051;
        src95 <= 16'hec3;
        src96 <= 16'h3f33;
        src97 <= 16'h90e0;
        src98 <= 16'h44f7;
        src99 <= 16'h7b12;
        src100 <= 16'h2d9c;
        src101 <= 16'habb7;
        src102 <= 16'h1a55;
        src103 <= 16'h5282;
        src104 <= 16'haff1;
        src105 <= 16'h3ac3;
        src106 <= 16'he5d9;
        src107 <= 16'he5e8;
        src108 <= 16'h224f;
        src109 <= 16'h3545;
        src110 <= 16'hdf0;
        src111 <= 16'h8e66;
        src112 <= 16'h5c1f;
        src113 <= 16'he383;
        src114 <= 16'hd84c;
        src115 <= 16'h934b;
        src116 <= 16'hc96e;
        src117 <= 16'ha28d;
        src118 <= 16'h313;
        src119 <= 16'hb8b7;
        src120 <= 16'h6703;
        src121 <= 16'hc602;
        src122 <= 16'hc559;
        src123 <= 16'h1eae;
        src124 <= 16'hb8c1;
        src125 <= 16'h42bc;
        src126 <= 16'hc42f;
        src127 <= 16'he191;
        src128 <= 16'h5b50;
        src129 <= 16'h4791;
        src130 <= 16'he62d;
        src131 <= 16'hb7c8;
        src132 <= 16'h1b49;
        src133 <= 16'h867a;
        src134 <= 16'hf210;
        src135 <= 16'h9c6d;
        src136 <= 16'hc1b6;
        src137 <= 16'h6446;
        src138 <= 16'h31b6;
        src139 <= 16'h2ab9;
        src140 <= 16'hb1d9;
        src141 <= 16'h3de6;
        src142 <= 16'h668a;
        src143 <= 16'h227a;
        src144 <= 16'hf2c;
        src145 <= 16'hb857;
        src146 <= 16'h5983;
        src147 <= 16'h6643;
        src148 <= 16'hd734;
        src149 <= 16'h866e;
        src150 <= 16'h6cb9;
        src151 <= 16'h49b5;
        src152 <= 16'h293c;
        src153 <= 16'he829;
        src154 <= 16'h16b2;
        src155 <= 16'h73fc;
        src156 <= 16'h792;
        src157 <= 16'h94c9;
        src158 <= 16'h3cfa;
        src159 <= 16'hf738;
        src160 <= 16'hfbfb;
        src161 <= 16'ha1f4;
        exp <= 24'h4f02aa;
        #1
        src0 <= 16'hc1c4;
        src1 <= 16'h4d25;
        src2 <= 16'h6a1d;
        src3 <= 16'hf241;
        src4 <= 16'hdaf7;
        src5 <= 16'h53ff;
        src6 <= 16'h9b1;
        src7 <= 16'ha5af;
        src8 <= 16'hd14c;
        src9 <= 16'ha8dd;
        src10 <= 16'h46ce;
        src11 <= 16'hda96;
        src12 <= 16'h7150;
        src13 <= 16'haffc;
        src14 <= 16'hf9ac;
        src15 <= 16'h4b45;
        src16 <= 16'h3d39;
        src17 <= 16'hb9;
        src18 <= 16'h7878;
        src19 <= 16'h9d85;
        src20 <= 16'h7a8d;
        src21 <= 16'hc464;
        src22 <= 16'h51b7;
        src23 <= 16'h469e;
        src24 <= 16'hc06d;
        src25 <= 16'hdebf;
        src26 <= 16'hfb53;
        src27 <= 16'h3e4e;
        src28 <= 16'h2803;
        src29 <= 16'hba58;
        src30 <= 16'h4cf5;
        src31 <= 16'he59d;
        src32 <= 16'hd67a;
        src33 <= 16'h2;
        src34 <= 16'habba;
        src35 <= 16'h746c;
        src36 <= 16'h16cf;
        src37 <= 16'h3732;
        src38 <= 16'hc812;
        src39 <= 16'h1fbf;
        src40 <= 16'h2f30;
        src41 <= 16'h3f7;
        src42 <= 16'h7835;
        src43 <= 16'h58b9;
        src44 <= 16'h67f3;
        src45 <= 16'h7b7e;
        src46 <= 16'h47e2;
        src47 <= 16'hf2cb;
        src48 <= 16'hc2d4;
        src49 <= 16'h419c;
        src50 <= 16'h5ee6;
        src51 <= 16'h2fa4;
        src52 <= 16'he58e;
        src53 <= 16'hcdc9;
        src54 <= 16'h4f67;
        src55 <= 16'hf40f;
        src56 <= 16'hc665;
        src57 <= 16'h26dd;
        src58 <= 16'hd998;
        src59 <= 16'hc5db;
        src60 <= 16'h2240;
        src61 <= 16'hde24;
        src62 <= 16'h9ed9;
        src63 <= 16'h7e07;
        src64 <= 16'hf0f;
        src65 <= 16'h2305;
        src66 <= 16'hf502;
        src67 <= 16'h671e;
        src68 <= 16'h9c7b;
        src69 <= 16'h6b31;
        src70 <= 16'hba6b;
        src71 <= 16'ha257;
        src72 <= 16'h7daa;
        src73 <= 16'haf2e;
        src74 <= 16'hb9cf;
        src75 <= 16'h36e6;
        src76 <= 16'hd6c8;
        src77 <= 16'h8418;
        src78 <= 16'h3a5f;
        src79 <= 16'hf7b0;
        src80 <= 16'hcedc;
        src81 <= 16'h4775;
        src82 <= 16'hc3a2;
        src83 <= 16'heae1;
        src84 <= 16'ha8f6;
        src85 <= 16'he765;
        src86 <= 16'h3160;
        src87 <= 16'h9a78;
        src88 <= 16'hdbbd;
        src89 <= 16'h1c00;
        src90 <= 16'h7265;
        src91 <= 16'ha336;
        src92 <= 16'h3a9b;
        src93 <= 16'h6031;
        src94 <= 16'hc350;
        src95 <= 16'h8b9a;
        src96 <= 16'h34f0;
        src97 <= 16'h14cd;
        src98 <= 16'hdcf0;
        src99 <= 16'h559d;
        src100 <= 16'h1f1f;
        src101 <= 16'he901;
        src102 <= 16'hd99d;
        src103 <= 16'h6600;
        src104 <= 16'h4354;
        src105 <= 16'h3ada;
        src106 <= 16'hf67f;
        src107 <= 16'heec1;
        src108 <= 16'h84ff;
        src109 <= 16'hb95;
        src110 <= 16'h28d1;
        src111 <= 16'h600c;
        src112 <= 16'h13b9;
        src113 <= 16'hb53d;
        src114 <= 16'h7a54;
        src115 <= 16'hc1d5;
        src116 <= 16'ha6fc;
        src117 <= 16'h55a0;
        src118 <= 16'h2c92;
        src119 <= 16'h190a;
        src120 <= 16'h1a7e;
        src121 <= 16'h725a;
        src122 <= 16'h63dd;
        src123 <= 16'heca6;
        src124 <= 16'h4a36;
        src125 <= 16'h5e0e;
        src126 <= 16'hc0be;
        src127 <= 16'h4188;
        src128 <= 16'hf10c;
        src129 <= 16'h55dd;
        src130 <= 16'hee6f;
        src131 <= 16'he7d9;
        src132 <= 16'h62ac;
        src133 <= 16'h4f4b;
        src134 <= 16'hc9f9;
        src135 <= 16'he911;
        src136 <= 16'he62;
        src137 <= 16'hdab5;
        src138 <= 16'h41b9;
        src139 <= 16'hc7;
        src140 <= 16'h6e1f;
        src141 <= 16'h4178;
        src142 <= 16'h7017;
        src143 <= 16'hbb11;
        src144 <= 16'h2623;
        src145 <= 16'h4b13;
        src146 <= 16'h8cdd;
        src147 <= 16'h5239;
        src148 <= 16'hf492;
        src149 <= 16'h1035;
        src150 <= 16'hf83d;
        src151 <= 16'h1e9f;
        src152 <= 16'he7f4;
        src153 <= 16'h7839;
        src154 <= 16'h8116;
        src155 <= 16'h665;
        src156 <= 16'h8e4a;
        src157 <= 16'hffed;
        src158 <= 16'h7331;
        src159 <= 16'hc5c9;
        src160 <= 16'hc745;
        src161 <= 16'h1eb5;
        exp <= 24'h52355c;
        #1
        src0 <= 16'h8483;
        src1 <= 16'h826f;
        src2 <= 16'h9e37;
        src3 <= 16'h82a4;
        src4 <= 16'h4eb1;
        src5 <= 16'h2b34;
        src6 <= 16'h8c17;
        src7 <= 16'h70f9;
        src8 <= 16'hb1f3;
        src9 <= 16'h4a12;
        src10 <= 16'h9c61;
        src11 <= 16'haa22;
        src12 <= 16'hedd4;
        src13 <= 16'h46d8;
        src14 <= 16'he0a4;
        src15 <= 16'hfa3e;
        src16 <= 16'h96b9;
        src17 <= 16'h17d;
        src18 <= 16'h900a;
        src19 <= 16'hd258;
        src20 <= 16'h5f05;
        src21 <= 16'hd8eb;
        src22 <= 16'h98bc;
        src23 <= 16'h1a24;
        src24 <= 16'he4d5;
        src25 <= 16'h1962;
        src26 <= 16'hf720;
        src27 <= 16'h6924;
        src28 <= 16'h2e00;
        src29 <= 16'hf3a4;
        src30 <= 16'h5b54;
        src31 <= 16'h350f;
        src32 <= 16'hf05c;
        src33 <= 16'h413f;
        src34 <= 16'h8dff;
        src35 <= 16'he596;
        src36 <= 16'h39e4;
        src37 <= 16'h7791;
        src38 <= 16'h65d1;
        src39 <= 16'h56d2;
        src40 <= 16'h3ef4;
        src41 <= 16'h1aee;
        src42 <= 16'h3243;
        src43 <= 16'he2a4;
        src44 <= 16'h1483;
        src45 <= 16'h2afd;
        src46 <= 16'hfcbb;
        src47 <= 16'hfa2d;
        src48 <= 16'h358d;
        src49 <= 16'h476f;
        src50 <= 16'h7aa3;
        src51 <= 16'hf5dd;
        src52 <= 16'h70dc;
        src53 <= 16'h8652;
        src54 <= 16'h2131;
        src55 <= 16'hab7b;
        src56 <= 16'h173d;
        src57 <= 16'h3502;
        src58 <= 16'hebc8;
        src59 <= 16'he017;
        src60 <= 16'h917b;
        src61 <= 16'h239;
        src62 <= 16'h7ba5;
        src63 <= 16'h3a3;
        src64 <= 16'h13b1;
        src65 <= 16'hec2e;
        src66 <= 16'h3451;
        src67 <= 16'h350b;
        src68 <= 16'ha1b6;
        src69 <= 16'h8162;
        src70 <= 16'hd819;
        src71 <= 16'he620;
        src72 <= 16'h6049;
        src73 <= 16'h1a31;
        src74 <= 16'hdf90;
        src75 <= 16'hb8b3;
        src76 <= 16'hde1e;
        src77 <= 16'ha019;
        src78 <= 16'he572;
        src79 <= 16'h3e39;
        src80 <= 16'h42d8;
        src81 <= 16'he0a1;
        src82 <= 16'ha5;
        src83 <= 16'h33d4;
        src84 <= 16'h2e7e;
        src85 <= 16'h57ed;
        src86 <= 16'h5165;
        src87 <= 16'h97c1;
        src88 <= 16'hece9;
        src89 <= 16'ha471;
        src90 <= 16'h517f;
        src91 <= 16'h8f90;
        src92 <= 16'hfb92;
        src93 <= 16'haa4d;
        src94 <= 16'hacc9;
        src95 <= 16'h1715;
        src96 <= 16'hcf0f;
        src97 <= 16'h1d32;
        src98 <= 16'hb37d;
        src99 <= 16'hbbf3;
        src100 <= 16'h2b2d;
        src101 <= 16'h8ce3;
        src102 <= 16'h3584;
        src103 <= 16'h5c62;
        src104 <= 16'h64a3;
        src105 <= 16'hcd2;
        src106 <= 16'h27d5;
        src107 <= 16'hbd49;
        src108 <= 16'h9f2f;
        src109 <= 16'h4cbb;
        src110 <= 16'hac5f;
        src111 <= 16'h9bf3;
        src112 <= 16'h876c;
        src113 <= 16'h2157;
        src114 <= 16'h3d75;
        src115 <= 16'h12be;
        src116 <= 16'he85b;
        src117 <= 16'h1737;
        src118 <= 16'h1a69;
        src119 <= 16'h31be;
        src120 <= 16'h186f;
        src121 <= 16'hff4;
        src122 <= 16'ha671;
        src123 <= 16'h9af7;
        src124 <= 16'h37a1;
        src125 <= 16'hc0ee;
        src126 <= 16'h8540;
        src127 <= 16'he6a1;
        src128 <= 16'hac34;
        src129 <= 16'h9a06;
        src130 <= 16'hd928;
        src131 <= 16'h259f;
        src132 <= 16'h3112;
        src133 <= 16'ha09c;
        src134 <= 16'h5002;
        src135 <= 16'h7442;
        src136 <= 16'h9fd3;
        src137 <= 16'hb539;
        src138 <= 16'hd3f9;
        src139 <= 16'h5b25;
        src140 <= 16'he66c;
        src141 <= 16'h7548;
        src142 <= 16'h93de;
        src143 <= 16'haab9;
        src144 <= 16'hf629;
        src145 <= 16'hfc47;
        src146 <= 16'hb765;
        src147 <= 16'h4eb1;
        src148 <= 16'h674a;
        src149 <= 16'hcf5d;
        src150 <= 16'h989;
        src151 <= 16'h668d;
        src152 <= 16'h2eb2;
        src153 <= 16'h38cd;
        src154 <= 16'hc8d8;
        src155 <= 16'h9d5c;
        src156 <= 16'h73e2;
        src157 <= 16'h5775;
        src158 <= 16'h3dbc;
        src159 <= 16'hceb8;
        src160 <= 16'h554e;
        src161 <= 16'hbc6c;
        exp <= 24'h4fb1c2;
        #1
        src0 <= 16'h7bde;
        src1 <= 16'h8827;
        src2 <= 16'h3db4;
        src3 <= 16'hc241;
        src4 <= 16'h2eb1;
        src5 <= 16'he49f;
        src6 <= 16'h497a;
        src7 <= 16'hcb66;
        src8 <= 16'h5aff;
        src9 <= 16'hf10d;
        src10 <= 16'h2656;
        src11 <= 16'he11c;
        src12 <= 16'h3603;
        src13 <= 16'h9328;
        src14 <= 16'h2d46;
        src15 <= 16'h29d2;
        src16 <= 16'h8be0;
        src17 <= 16'h2843;
        src18 <= 16'h107a;
        src19 <= 16'h5b0d;
        src20 <= 16'h7a;
        src21 <= 16'h99e3;
        src22 <= 16'h8ffb;
        src23 <= 16'h8389;
        src24 <= 16'h75ee;
        src25 <= 16'h717a;
        src26 <= 16'h6033;
        src27 <= 16'hedb1;
        src28 <= 16'h6d05;
        src29 <= 16'h897e;
        src30 <= 16'he323;
        src31 <= 16'h3e0;
        src32 <= 16'he41e;
        src33 <= 16'hf6c7;
        src34 <= 16'h79e5;
        src35 <= 16'hefc2;
        src36 <= 16'h58e6;
        src37 <= 16'h7681;
        src38 <= 16'h9e8d;
        src39 <= 16'hcae3;
        src40 <= 16'hd110;
        src41 <= 16'hdc2b;
        src42 <= 16'h1774;
        src43 <= 16'h9f0a;
        src44 <= 16'h6d85;
        src45 <= 16'h9b34;
        src46 <= 16'h8be5;
        src47 <= 16'hcb3;
        src48 <= 16'habc9;
        src49 <= 16'h2197;
        src50 <= 16'h74aa;
        src51 <= 16'h774;
        src52 <= 16'hfaf5;
        src53 <= 16'h9704;
        src54 <= 16'h3f27;
        src55 <= 16'h833f;
        src56 <= 16'h7fac;
        src57 <= 16'h1a71;
        src58 <= 16'hd3df;
        src59 <= 16'hb002;
        src60 <= 16'h4d7b;
        src61 <= 16'ha7a1;
        src62 <= 16'h3035;
        src63 <= 16'hdf2b;
        src64 <= 16'he49c;
        src65 <= 16'h1682;
        src66 <= 16'h7d70;
        src67 <= 16'ha828;
        src68 <= 16'hf85c;
        src69 <= 16'hff24;
        src70 <= 16'h30ad;
        src71 <= 16'h118a;
        src72 <= 16'h4718;
        src73 <= 16'h3b5c;
        src74 <= 16'h4056;
        src75 <= 16'h92e3;
        src76 <= 16'hd23d;
        src77 <= 16'h8a3b;
        src78 <= 16'h5502;
        src79 <= 16'h66c6;
        src80 <= 16'hde0;
        src81 <= 16'ha85;
        src82 <= 16'h2adc;
        src83 <= 16'h7cbf;
        src84 <= 16'he63b;
        src85 <= 16'he15e;
        src86 <= 16'h8a6c;
        src87 <= 16'h7bc6;
        src88 <= 16'hbfec;
        src89 <= 16'h2347;
        src90 <= 16'h3ab7;
        src91 <= 16'h33dd;
        src92 <= 16'h926f;
        src93 <= 16'h2f4a;
        src94 <= 16'h6e1e;
        src95 <= 16'h1417;
        src96 <= 16'hbf3a;
        src97 <= 16'h48b9;
        src98 <= 16'h9482;
        src99 <= 16'h8ef1;
        src100 <= 16'hb3f0;
        src101 <= 16'h4c22;
        src102 <= 16'hcb59;
        src103 <= 16'h8fb5;
        src104 <= 16'h3a51;
        src105 <= 16'he383;
        src106 <= 16'h5df0;
        src107 <= 16'hdb62;
        src108 <= 16'h9b5a;
        src109 <= 16'h7c83;
        src110 <= 16'h3494;
        src111 <= 16'hec55;
        src112 <= 16'hca30;
        src113 <= 16'h51e5;
        src114 <= 16'h5750;
        src115 <= 16'h7724;
        src116 <= 16'hfb7a;
        src117 <= 16'hfb2b;
        src118 <= 16'h268b;
        src119 <= 16'h7219;
        src120 <= 16'hedff;
        src121 <= 16'he206;
        src122 <= 16'hfa5c;
        src123 <= 16'hffd5;
        src124 <= 16'hb944;
        src125 <= 16'hdda1;
        src126 <= 16'he59;
        src127 <= 16'h2157;
        src128 <= 16'h10c3;
        src129 <= 16'hdec5;
        src130 <= 16'h3072;
        src131 <= 16'h77a0;
        src132 <= 16'hff92;
        src133 <= 16'h9949;
        src134 <= 16'h5693;
        src135 <= 16'h6535;
        src136 <= 16'h826e;
        src137 <= 16'h76f7;
        src138 <= 16'hecee;
        src139 <= 16'h8c18;
        src140 <= 16'h4e3e;
        src141 <= 16'h3b38;
        src142 <= 16'h640c;
        src143 <= 16'h878c;
        src144 <= 16'h97b;
        src145 <= 16'h90b8;
        src146 <= 16'hc010;
        src147 <= 16'hc805;
        src148 <= 16'hc21c;
        src149 <= 16'h2d54;
        src150 <= 16'h18e3;
        src151 <= 16'ha12a;
        src152 <= 16'hfc0b;
        src153 <= 16'hffc1;
        src154 <= 16'h452b;
        src155 <= 16'h7d9;
        src156 <= 16'h60e3;
        src157 <= 16'h22e5;
        src158 <= 16'h1b84;
        src159 <= 16'had77;
        src160 <= 16'hb568;
        src161 <= 16'hc63d;
        exp <= 24'h5180a8;
        #1
        src0 <= 16'h48d2;
        src1 <= 16'h2748;
        src2 <= 16'hbfca;
        src3 <= 16'hd1d8;
        src4 <= 16'h169f;
        src5 <= 16'hdbbe;
        src6 <= 16'hbff4;
        src7 <= 16'h5f17;
        src8 <= 16'h6a58;
        src9 <= 16'h22dc;
        src10 <= 16'h60ae;
        src11 <= 16'h34ee;
        src12 <= 16'hcc2e;
        src13 <= 16'ha34d;
        src14 <= 16'ha337;
        src15 <= 16'h79d;
        src16 <= 16'h1b9f;
        src17 <= 16'heb08;
        src18 <= 16'h82f5;
        src19 <= 16'h5860;
        src20 <= 16'habef;
        src21 <= 16'hc754;
        src22 <= 16'h9276;
        src23 <= 16'h65e;
        src24 <= 16'hf6b7;
        src25 <= 16'h162d;
        src26 <= 16'h3f3b;
        src27 <= 16'h94b7;
        src28 <= 16'hb0d6;
        src29 <= 16'hf74;
        src30 <= 16'he860;
        src31 <= 16'h98cb;
        src32 <= 16'h7a0c;
        src33 <= 16'h9cf4;
        src34 <= 16'h2ceb;
        src35 <= 16'h4dd9;
        src36 <= 16'h529d;
        src37 <= 16'hc61f;
        src38 <= 16'h9431;
        src39 <= 16'hc116;
        src40 <= 16'hac33;
        src41 <= 16'h446a;
        src42 <= 16'h2faf;
        src43 <= 16'hc775;
        src44 <= 16'h1335;
        src45 <= 16'ha357;
        src46 <= 16'hb7ad;
        src47 <= 16'h61b1;
        src48 <= 16'h9147;
        src49 <= 16'h22f2;
        src50 <= 16'hd6c5;
        src51 <= 16'h1be1;
        src52 <= 16'h7700;
        src53 <= 16'h5b74;
        src54 <= 16'h5da2;
        src55 <= 16'h558e;
        src56 <= 16'hf6cb;
        src57 <= 16'h8d97;
        src58 <= 16'h37b5;
        src59 <= 16'hfeb;
        src60 <= 16'h9a7e;
        src61 <= 16'he688;
        src62 <= 16'h1ead;
        src63 <= 16'hdb54;
        src64 <= 16'hd975;
        src65 <= 16'hef1d;
        src66 <= 16'h27a6;
        src67 <= 16'h3c82;
        src68 <= 16'he9d;
        src69 <= 16'hc611;
        src70 <= 16'hbed4;
        src71 <= 16'hf390;
        src72 <= 16'hf9b5;
        src73 <= 16'hc178;
        src74 <= 16'hb79b;
        src75 <= 16'hdbdb;
        src76 <= 16'hd8af;
        src77 <= 16'h4be9;
        src78 <= 16'he6a;
        src79 <= 16'hc1e6;
        src80 <= 16'h2bce;
        src81 <= 16'h4b8a;
        src82 <= 16'hfea9;
        src83 <= 16'h34c9;
        src84 <= 16'h7edb;
        src85 <= 16'h50cc;
        src86 <= 16'h5451;
        src87 <= 16'h1a8a;
        src88 <= 16'h91db;
        src89 <= 16'h43d3;
        src90 <= 16'h6c50;
        src91 <= 16'h59ec;
        src92 <= 16'hb385;
        src93 <= 16'h30bc;
        src94 <= 16'ha027;
        src95 <= 16'h5259;
        src96 <= 16'ha75b;
        src97 <= 16'hcf90;
        src98 <= 16'h688d;
        src99 <= 16'hd665;
        src100 <= 16'hf952;
        src101 <= 16'h58d0;
        src102 <= 16'h9c0f;
        src103 <= 16'h5994;
        src104 <= 16'h8b;
        src105 <= 16'he8b0;
        src106 <= 16'h5492;
        src107 <= 16'hc63d;
        src108 <= 16'hdf6;
        src109 <= 16'hc7e6;
        src110 <= 16'h16c9;
        src111 <= 16'h64ce;
        src112 <= 16'hfd47;
        src113 <= 16'hade3;
        src114 <= 16'h483a;
        src115 <= 16'h7294;
        src116 <= 16'h28b8;
        src117 <= 16'h3780;
        src118 <= 16'h7328;
        src119 <= 16'h5210;
        src120 <= 16'hfe00;
        src121 <= 16'he859;
        src122 <= 16'h5700;
        src123 <= 16'h5336;
        src124 <= 16'h399d;
        src125 <= 16'hd0e8;
        src126 <= 16'h4f55;
        src127 <= 16'h8002;
        src128 <= 16'heeb6;
        src129 <= 16'h222;
        src130 <= 16'h433e;
        src131 <= 16'hd56e;
        src132 <= 16'h85c9;
        src133 <= 16'h6c99;
        src134 <= 16'h21c1;
        src135 <= 16'h8ed9;
        src136 <= 16'h4b25;
        src137 <= 16'h3271;
        src138 <= 16'hacf4;
        src139 <= 16'h5c54;
        src140 <= 16'hff50;
        src141 <= 16'ha28;
        src142 <= 16'h8269;
        src143 <= 16'h78f2;
        src144 <= 16'h60da;
        src145 <= 16'h9b09;
        src146 <= 16'h3de1;
        src147 <= 16'ha599;
        src148 <= 16'h48cb;
        src149 <= 16'hbed3;
        src150 <= 16'hae73;
        src151 <= 16'hf141;
        src152 <= 16'h1b46;
        src153 <= 16'hb7db;
        src154 <= 16'hf3cf;
        src155 <= 16'h79e1;
        src156 <= 16'h5c6f;
        src157 <= 16'hef22;
        src158 <= 16'h42cc;
        src159 <= 16'h5dee;
        src160 <= 16'h544b;
        src161 <= 16'hf9e6;
        exp <= 24'h50620c;
        #1
        src0 <= 16'hca6c;
        src1 <= 16'hc495;
        src2 <= 16'h9929;
        src3 <= 16'hc3a6;
        src4 <= 16'he4ac;
        src5 <= 16'hdcd;
        src6 <= 16'hcee4;
        src7 <= 16'hcaa7;
        src8 <= 16'h1959;
        src9 <= 16'hb585;
        src10 <= 16'h60d2;
        src11 <= 16'h5752;
        src12 <= 16'h7a56;
        src13 <= 16'h21ac;
        src14 <= 16'h9c9d;
        src15 <= 16'hcae1;
        src16 <= 16'h3bd2;
        src17 <= 16'he652;
        src18 <= 16'hc6fa;
        src19 <= 16'hfb8a;
        src20 <= 16'h7f63;
        src21 <= 16'hb65e;
        src22 <= 16'hacc8;
        src23 <= 16'h62e5;
        src24 <= 16'hf2ef;
        src25 <= 16'hafa0;
        src26 <= 16'hc297;
        src27 <= 16'hecbf;
        src28 <= 16'hc2b0;
        src29 <= 16'hb019;
        src30 <= 16'h8e9d;
        src31 <= 16'h1ea1;
        src32 <= 16'h3990;
        src33 <= 16'ha2d2;
        src34 <= 16'hc4fa;
        src35 <= 16'h4fc0;
        src36 <= 16'h899e;
        src37 <= 16'h1791;
        src38 <= 16'hb7c5;
        src39 <= 16'h31d1;
        src40 <= 16'h3651;
        src41 <= 16'h644e;
        src42 <= 16'h2417;
        src43 <= 16'hd868;
        src44 <= 16'h502;
        src45 <= 16'h1f12;
        src46 <= 16'hdece;
        src47 <= 16'hed75;
        src48 <= 16'h26c4;
        src49 <= 16'hd58e;
        src50 <= 16'hda4e;
        src51 <= 16'h340;
        src52 <= 16'hdc06;
        src53 <= 16'hed2a;
        src54 <= 16'h9d0b;
        src55 <= 16'h8b92;
        src56 <= 16'h1792;
        src57 <= 16'h7952;
        src58 <= 16'h4925;
        src59 <= 16'h3576;
        src60 <= 16'hbfad;
        src61 <= 16'h334b;
        src62 <= 16'hb828;
        src63 <= 16'hd3d3;
        src64 <= 16'he2ef;
        src65 <= 16'h2939;
        src66 <= 16'h2a3f;
        src67 <= 16'he2d7;
        src68 <= 16'he80d;
        src69 <= 16'h4343;
        src70 <= 16'hf472;
        src71 <= 16'h943a;
        src72 <= 16'h7369;
        src73 <= 16'hc4de;
        src74 <= 16'h4587;
        src75 <= 16'hf152;
        src76 <= 16'h94b2;
        src77 <= 16'hc259;
        src78 <= 16'h852;
        src79 <= 16'h8ab2;
        src80 <= 16'ha0ee;
        src81 <= 16'h61e4;
        src82 <= 16'h5162;
        src83 <= 16'h5d22;
        src84 <= 16'h8ad7;
        src85 <= 16'h39f4;
        src86 <= 16'h2eae;
        src87 <= 16'h14f8;
        src88 <= 16'hc1f4;
        src89 <= 16'hdcc5;
        src90 <= 16'hf2ae;
        src91 <= 16'h40d6;
        src92 <= 16'ha565;
        src93 <= 16'h1d36;
        src94 <= 16'hf214;
        src95 <= 16'ha7cd;
        src96 <= 16'h52cd;
        src97 <= 16'h4794;
        src98 <= 16'hbbe8;
        src99 <= 16'hf99;
        src100 <= 16'h6dfc;
        src101 <= 16'hc74d;
        src102 <= 16'hcc55;
        src103 <= 16'h1785;
        src104 <= 16'h8ec0;
        src105 <= 16'h8f3a;
        src106 <= 16'h3509;
        src107 <= 16'h1461;
        src108 <= 16'h97da;
        src109 <= 16'h16c3;
        src110 <= 16'h3cc9;
        src111 <= 16'he85d;
        src112 <= 16'h7707;
        src113 <= 16'h34b2;
        src114 <= 16'hb834;
        src115 <= 16'hcf2f;
        src116 <= 16'hbb8f;
        src117 <= 16'hf9ef;
        src118 <= 16'h6db;
        src119 <= 16'ha50d;
        src120 <= 16'h593d;
        src121 <= 16'h1649;
        src122 <= 16'h2125;
        src123 <= 16'h8237;
        src124 <= 16'h626a;
        src125 <= 16'h6575;
        src126 <= 16'h6302;
        src127 <= 16'h23f2;
        src128 <= 16'h6108;
        src129 <= 16'h3741;
        src130 <= 16'h9749;
        src131 <= 16'h3485;
        src132 <= 16'hfaf7;
        src133 <= 16'h253c;
        src134 <= 16'he4a2;
        src135 <= 16'h303f;
        src136 <= 16'hc883;
        src137 <= 16'h996a;
        src138 <= 16'hdd72;
        src139 <= 16'h3ac8;
        src140 <= 16'hf5f4;
        src141 <= 16'h950;
        src142 <= 16'h988c;
        src143 <= 16'h81d3;
        src144 <= 16'h224d;
        src145 <= 16'h128f;
        src146 <= 16'ha2c1;
        src147 <= 16'h4bc4;
        src148 <= 16'h96eb;
        src149 <= 16'h1c32;
        src150 <= 16'h2c37;
        src151 <= 16'h63e2;
        src152 <= 16'h26cd;
        src153 <= 16'h8c37;
        src154 <= 16'he37d;
        src155 <= 16'h4f55;
        src156 <= 16'hd13e;
        src157 <= 16'hd6a5;
        src158 <= 16'he2f2;
        src159 <= 16'h3dcc;
        src160 <= 16'h55df;
        src161 <= 16'hade4;
        exp <= 24'h5200df;
        #1
        src0 <= 16'hf1ee;
        src1 <= 16'h5bf0;
        src2 <= 16'hed9d;
        src3 <= 16'h7a26;
        src4 <= 16'h4b81;
        src5 <= 16'h2a27;
        src6 <= 16'h4b12;
        src7 <= 16'h5098;
        src8 <= 16'h3eef;
        src9 <= 16'he6e5;
        src10 <= 16'ha0ad;
        src11 <= 16'h21e0;
        src12 <= 16'h4cc;
        src13 <= 16'hc8ad;
        src14 <= 16'h1bd9;
        src15 <= 16'hbf96;
        src16 <= 16'h6096;
        src17 <= 16'hd495;
        src18 <= 16'h7f9f;
        src19 <= 16'h8d86;
        src20 <= 16'h7d1d;
        src21 <= 16'hfda0;
        src22 <= 16'h1688;
        src23 <= 16'h1abf;
        src24 <= 16'h460;
        src25 <= 16'h799;
        src26 <= 16'ha511;
        src27 <= 16'hde54;
        src28 <= 16'hed36;
        src29 <= 16'h73e8;
        src30 <= 16'h78a7;
        src31 <= 16'hc2aa;
        src32 <= 16'h8240;
        src33 <= 16'h3510;
        src34 <= 16'h3830;
        src35 <= 16'ha00a;
        src36 <= 16'h156e;
        src37 <= 16'h657e;
        src38 <= 16'hff20;
        src39 <= 16'h73ac;
        src40 <= 16'hed44;
        src41 <= 16'h5cdb;
        src42 <= 16'hce55;
        src43 <= 16'hf600;
        src44 <= 16'hbccb;
        src45 <= 16'h4352;
        src46 <= 16'h610f;
        src47 <= 16'h4d25;
        src48 <= 16'h512e;
        src49 <= 16'h4fb9;
        src50 <= 16'h61bd;
        src51 <= 16'h144a;
        src52 <= 16'ha44;
        src53 <= 16'h3587;
        src54 <= 16'hd8bc;
        src55 <= 16'h6e5;
        src56 <= 16'hc4d9;
        src57 <= 16'h6416;
        src58 <= 16'h3f4;
        src59 <= 16'h12eb;
        src60 <= 16'hd8a7;
        src61 <= 16'h2fc7;
        src62 <= 16'hf122;
        src63 <= 16'h797a;
        src64 <= 16'h62e1;
        src65 <= 16'h4119;
        src66 <= 16'h2cf0;
        src67 <= 16'h139d;
        src68 <= 16'h9ac2;
        src69 <= 16'h66df;
        src70 <= 16'h815c;
        src71 <= 16'h5a40;
        src72 <= 16'h40b5;
        src73 <= 16'h29b1;
        src74 <= 16'he133;
        src75 <= 16'h228d;
        src76 <= 16'hafef;
        src77 <= 16'h2903;
        src78 <= 16'hcfe7;
        src79 <= 16'hc36;
        src80 <= 16'he728;
        src81 <= 16'hd7d3;
        src82 <= 16'h3670;
        src83 <= 16'hdbbf;
        src84 <= 16'h8419;
        src85 <= 16'h610e;
        src86 <= 16'hccc6;
        src87 <= 16'h724f;
        src88 <= 16'hb52e;
        src89 <= 16'hd8d;
        src90 <= 16'h4e49;
        src91 <= 16'h670a;
        src92 <= 16'h63fc;
        src93 <= 16'hd763;
        src94 <= 16'hb45c;
        src95 <= 16'h801d;
        src96 <= 16'hddb7;
        src97 <= 16'h9741;
        src98 <= 16'h1fe;
        src99 <= 16'hdd90;
        src100 <= 16'h74f8;
        src101 <= 16'h620c;
        src102 <= 16'h37ee;
        src103 <= 16'h1601;
        src104 <= 16'hec59;
        src105 <= 16'heca4;
        src106 <= 16'hf19b;
        src107 <= 16'hf3f6;
        src108 <= 16'h66d9;
        src109 <= 16'h28b1;
        src110 <= 16'h4751;
        src111 <= 16'h614e;
        src112 <= 16'h9998;
        src113 <= 16'hf6a5;
        src114 <= 16'h2153;
        src115 <= 16'h72a;
        src116 <= 16'h1101;
        src117 <= 16'he944;
        src118 <= 16'haf4c;
        src119 <= 16'h4979;
        src120 <= 16'hd164;
        src121 <= 16'h19a1;
        src122 <= 16'h1de5;
        src123 <= 16'h4a5f;
        src124 <= 16'h2bd8;
        src125 <= 16'hc6d4;
        src126 <= 16'h346a;
        src127 <= 16'h5ede;
        src128 <= 16'h5c75;
        src129 <= 16'h6166;
        src130 <= 16'hda6b;
        src131 <= 16'he068;
        src132 <= 16'h473a;
        src133 <= 16'h9f5c;
        src134 <= 16'h4fe1;
        src135 <= 16'hc06;
        src136 <= 16'h7519;
        src137 <= 16'h4b0;
        src138 <= 16'hc4df;
        src139 <= 16'hd407;
        src140 <= 16'hec6b;
        src141 <= 16'hb3a8;
        src142 <= 16'h425;
        src143 <= 16'he2bb;
        src144 <= 16'had79;
        src145 <= 16'ha4c3;
        src146 <= 16'h9c93;
        src147 <= 16'hf85;
        src148 <= 16'h8069;
        src149 <= 16'h1075;
        src150 <= 16'hd8a5;
        src151 <= 16'hd493;
        src152 <= 16'h8603;
        src153 <= 16'h597f;
        src154 <= 16'h4d7b;
        src155 <= 16'he1b8;
        src156 <= 16'hf424;
        src157 <= 16'hdce3;
        src158 <= 16'hae31;
        src159 <= 16'h28f3;
        src160 <= 16'h1c1a;
        src161 <= 16'hb537;
        exp <= 24'h4d6674;
        #1
        src0 <= 16'h1ea;
        src1 <= 16'ha1dc;
        src2 <= 16'had8a;
        src3 <= 16'h803f;
        src4 <= 16'ha20c;
        src5 <= 16'h2035;
        src6 <= 16'hc20f;
        src7 <= 16'h8d3f;
        src8 <= 16'h9e05;
        src9 <= 16'ha716;
        src10 <= 16'hf60;
        src11 <= 16'hc3e1;
        src12 <= 16'hd582;
        src13 <= 16'h76e5;
        src14 <= 16'h4ea6;
        src15 <= 16'h7f9d;
        src16 <= 16'ha8da;
        src17 <= 16'h3eac;
        src18 <= 16'h8411;
        src19 <= 16'h8802;
        src20 <= 16'h872e;
        src21 <= 16'hd801;
        src22 <= 16'h985f;
        src23 <= 16'h47ed;
        src24 <= 16'h4caa;
        src25 <= 16'h6478;
        src26 <= 16'hc9a2;
        src27 <= 16'h1360;
        src28 <= 16'h3d7e;
        src29 <= 16'h3a4f;
        src30 <= 16'h4ee0;
        src31 <= 16'h8300;
        src32 <= 16'hfd25;
        src33 <= 16'h9fea;
        src34 <= 16'ha0a7;
        src35 <= 16'hd177;
        src36 <= 16'hf209;
        src37 <= 16'h4a5e;
        src38 <= 16'hbb0a;
        src39 <= 16'h3bf5;
        src40 <= 16'h5fdf;
        src41 <= 16'h87ff;
        src42 <= 16'h8384;
        src43 <= 16'h9a37;
        src44 <= 16'h9adc;
        src45 <= 16'h4adf;
        src46 <= 16'hde9b;
        src47 <= 16'hc1f0;
        src48 <= 16'h2c8d;
        src49 <= 16'hb2a7;
        src50 <= 16'hc4b3;
        src51 <= 16'h7543;
        src52 <= 16'hb3a3;
        src53 <= 16'h1680;
        src54 <= 16'h680c;
        src55 <= 16'hf413;
        src56 <= 16'h4c68;
        src57 <= 16'hf436;
        src58 <= 16'hf582;
        src59 <= 16'h9325;
        src60 <= 16'h2feb;
        src61 <= 16'h929e;
        src62 <= 16'hee7b;
        src63 <= 16'h4cdc;
        src64 <= 16'hbf9b;
        src65 <= 16'h7c45;
        src66 <= 16'he14a;
        src67 <= 16'hb784;
        src68 <= 16'hf597;
        src69 <= 16'he6db;
        src70 <= 16'h2a74;
        src71 <= 16'h33ff;
        src72 <= 16'hfcaf;
        src73 <= 16'hecaa;
        src74 <= 16'hcb92;
        src75 <= 16'hbd2f;
        src76 <= 16'h2fee;
        src77 <= 16'hb0b8;
        src78 <= 16'h56af;
        src79 <= 16'h68cb;
        src80 <= 16'h510b;
        src81 <= 16'h48f9;
        src82 <= 16'h6338;
        src83 <= 16'h2c11;
        src84 <= 16'heecf;
        src85 <= 16'hc3c2;
        src86 <= 16'h69b;
        src87 <= 16'h4407;
        src88 <= 16'hae50;
        src89 <= 16'hf1f9;
        src90 <= 16'h557e;
        src91 <= 16'ha3fb;
        src92 <= 16'h55d2;
        src93 <= 16'hbe80;
        src94 <= 16'h1ed0;
        src95 <= 16'h84d2;
        src96 <= 16'h5fc;
        src97 <= 16'h9bc0;
        src98 <= 16'h6148;
        src99 <= 16'h2570;
        src100 <= 16'hdd64;
        src101 <= 16'h8997;
        src102 <= 16'h4768;
        src103 <= 16'h167c;
        src104 <= 16'h7993;
        src105 <= 16'h528a;
        src106 <= 16'h656b;
        src107 <= 16'h44be;
        src108 <= 16'h6e1b;
        src109 <= 16'haf85;
        src110 <= 16'hce2b;
        src111 <= 16'hb81c;
        src112 <= 16'hfbb5;
        src113 <= 16'h4055;
        src114 <= 16'hcaa;
        src115 <= 16'h9f0c;
        src116 <= 16'hc43d;
        src117 <= 16'h6faf;
        src118 <= 16'h59a7;
        src119 <= 16'hc2d1;
        src120 <= 16'h8e9;
        src121 <= 16'h1fb9;
        src122 <= 16'hb445;
        src123 <= 16'he3c;
        src124 <= 16'h85b3;
        src125 <= 16'hca4c;
        src126 <= 16'hea22;
        src127 <= 16'ha303;
        src128 <= 16'h9d4b;
        src129 <= 16'h47e5;
        src130 <= 16'hde58;
        src131 <= 16'hb7b2;
        src132 <= 16'h686c;
        src133 <= 16'hf07d;
        src134 <= 16'hfa63;
        src135 <= 16'hdf42;
        src136 <= 16'h85a8;
        src137 <= 16'h26ab;
        src138 <= 16'hfe83;
        src139 <= 16'h9b37;
        src140 <= 16'h7f75;
        src141 <= 16'h48f7;
        src142 <= 16'hdee0;
        src143 <= 16'h3c43;
        src144 <= 16'hb6e6;
        src145 <= 16'h571a;
        src146 <= 16'h7335;
        src147 <= 16'hc516;
        src148 <= 16'h2795;
        src149 <= 16'h4a0f;
        src150 <= 16'hfcbc;
        src151 <= 16'hc50c;
        src152 <= 16'h96fd;
        src153 <= 16'hc305;
        src154 <= 16'hb3d6;
        src155 <= 16'h89e8;
        src156 <= 16'h321b;
        src157 <= 16'h424a;
        src158 <= 16'h80d4;
        src159 <= 16'h7130;
        src160 <= 16'h3e91;
        src161 <= 16'h9564;
        exp <= 24'h55bb33;
        #1
        src0 <= 16'h804b;
        src1 <= 16'h9889;
        src2 <= 16'h268d;
        src3 <= 16'h7837;
        src4 <= 16'hb973;
        src5 <= 16'h41fa;
        src6 <= 16'h98ef;
        src7 <= 16'h7810;
        src8 <= 16'h4156;
        src9 <= 16'h19bb;
        src10 <= 16'ha63b;
        src11 <= 16'h6852;
        src12 <= 16'h444b;
        src13 <= 16'h9acb;
        src14 <= 16'hc060;
        src15 <= 16'h517d;
        src16 <= 16'h756b;
        src17 <= 16'h3372;
        src18 <= 16'he953;
        src19 <= 16'h23fd;
        src20 <= 16'he350;
        src21 <= 16'he3d0;
        src22 <= 16'heb9e;
        src23 <= 16'h27a9;
        src24 <= 16'h9aea;
        src25 <= 16'hf53f;
        src26 <= 16'hb4c7;
        src27 <= 16'hb3b4;
        src28 <= 16'h87;
        src29 <= 16'h6184;
        src30 <= 16'h63e0;
        src31 <= 16'hf6d8;
        src32 <= 16'he270;
        src33 <= 16'h5355;
        src34 <= 16'h6016;
        src35 <= 16'h7cc3;
        src36 <= 16'h6e23;
        src37 <= 16'hc521;
        src38 <= 16'h3a6c;
        src39 <= 16'h21ca;
        src40 <= 16'hc103;
        src41 <= 16'had9c;
        src42 <= 16'hfaeb;
        src43 <= 16'hddcc;
        src44 <= 16'h5da9;
        src45 <= 16'hd9ef;
        src46 <= 16'h695a;
        src47 <= 16'he0eb;
        src48 <= 16'h9e08;
        src49 <= 16'h6f9a;
        src50 <= 16'hb5ab;
        src51 <= 16'he31c;
        src52 <= 16'h1a86;
        src53 <= 16'hb037;
        src54 <= 16'h2649;
        src55 <= 16'hab14;
        src56 <= 16'hefa4;
        src57 <= 16'hb4e6;
        src58 <= 16'h1b17;
        src59 <= 16'h2d98;
        src60 <= 16'h8649;
        src61 <= 16'h6572;
        src62 <= 16'h2bfb;
        src63 <= 16'h798e;
        src64 <= 16'h76ab;
        src65 <= 16'hbbd5;
        src66 <= 16'h74f7;
        src67 <= 16'h64c0;
        src68 <= 16'hee88;
        src69 <= 16'he709;
        src70 <= 16'h4bf5;
        src71 <= 16'hf9d7;
        src72 <= 16'hf6b4;
        src73 <= 16'h5410;
        src74 <= 16'ha419;
        src75 <= 16'hed26;
        src76 <= 16'h4639;
        src77 <= 16'h6b7b;
        src78 <= 16'h3b5b;
        src79 <= 16'h1d4c;
        src80 <= 16'ha2cf;
        src81 <= 16'hee64;
        src82 <= 16'h2cc6;
        src83 <= 16'h79c;
        src84 <= 16'h4440;
        src85 <= 16'hd45d;
        src86 <= 16'h9b22;
        src87 <= 16'h7dad;
        src88 <= 16'he1ce;
        src89 <= 16'h94c7;
        src90 <= 16'h2460;
        src91 <= 16'hfaa6;
        src92 <= 16'hcf31;
        src93 <= 16'hec89;
        src94 <= 16'hc57b;
        src95 <= 16'hc697;
        src96 <= 16'h4eab;
        src97 <= 16'h9aaa;
        src98 <= 16'h917f;
        src99 <= 16'hbd6f;
        src100 <= 16'h7dc9;
        src101 <= 16'hae78;
        src102 <= 16'hbac4;
        src103 <= 16'h127f;
        src104 <= 16'h7c45;
        src105 <= 16'h367b;
        src106 <= 16'heb9c;
        src107 <= 16'hd33d;
        src108 <= 16'h71b3;
        src109 <= 16'hbc0;
        src110 <= 16'hbc89;
        src111 <= 16'h9895;
        src112 <= 16'h4271;
        src113 <= 16'hf478;
        src114 <= 16'he97;
        src115 <= 16'h2730;
        src116 <= 16'h7d73;
        src117 <= 16'h848;
        src118 <= 16'ha17;
        src119 <= 16'hce8c;
        src120 <= 16'h951f;
        src121 <= 16'hf2b8;
        src122 <= 16'hd047;
        src123 <= 16'h1226;
        src124 <= 16'hae0;
        src125 <= 16'hafc;
        src126 <= 16'hf9ec;
        src127 <= 16'hcd3e;
        src128 <= 16'heb4c;
        src129 <= 16'hd9a0;
        src130 <= 16'h7920;
        src131 <= 16'h300a;
        src132 <= 16'hdcb5;
        src133 <= 16'h4ef6;
        src134 <= 16'hb5f;
        src135 <= 16'h4079;
        src136 <= 16'hc323;
        src137 <= 16'h4e55;
        src138 <= 16'h71ef;
        src139 <= 16'h6e74;
        src140 <= 16'h55a6;
        src141 <= 16'hfc46;
        src142 <= 16'h2414;
        src143 <= 16'hfa25;
        src144 <= 16'he10d;
        src145 <= 16'hcb7b;
        src146 <= 16'h215f;
        src147 <= 16'h24c5;
        src148 <= 16'hde11;
        src149 <= 16'hee7a;
        src150 <= 16'h4658;
        src151 <= 16'hd2c5;
        src152 <= 16'hacc7;
        src153 <= 16'h2c59;
        src154 <= 16'hf0b5;
        src155 <= 16'h6c01;
        src156 <= 16'h2ab1;
        src157 <= 16'hce5e;
        src158 <= 16'ha63a;
        src159 <= 16'h216a;
        src160 <= 16'h5a64;
        src161 <= 16'h772a;
        exp <= 24'h55e382;
        #1
        src0 <= 16'hf470;
        src1 <= 16'h117b;
        src2 <= 16'hb2ee;
        src3 <= 16'h1995;
        src4 <= 16'h122f;
        src5 <= 16'h64b9;
        src6 <= 16'h19e;
        src7 <= 16'hc0d8;
        src8 <= 16'hc4c4;
        src9 <= 16'h4bcd;
        src10 <= 16'h61b7;
        src11 <= 16'h4c97;
        src12 <= 16'h3121;
        src13 <= 16'ha006;
        src14 <= 16'h824;
        src15 <= 16'hf04f;
        src16 <= 16'had4;
        src17 <= 16'h6e8d;
        src18 <= 16'hfbaf;
        src19 <= 16'h29d9;
        src20 <= 16'h610d;
        src21 <= 16'h76f4;
        src22 <= 16'h4628;
        src23 <= 16'h3a96;
        src24 <= 16'h38cc;
        src25 <= 16'h51a3;
        src26 <= 16'h4267;
        src27 <= 16'he9d0;
        src28 <= 16'hc1a1;
        src29 <= 16'h9d5e;
        src30 <= 16'hd9b8;
        src31 <= 16'h5ec7;
        src32 <= 16'h2334;
        src33 <= 16'h850e;
        src34 <= 16'h6dc0;
        src35 <= 16'h6e9a;
        src36 <= 16'hc641;
        src37 <= 16'hd07b;
        src38 <= 16'h9662;
        src39 <= 16'h503c;
        src40 <= 16'hcdaa;
        src41 <= 16'h411a;
        src42 <= 16'h895b;
        src43 <= 16'hfceb;
        src44 <= 16'h3e43;
        src45 <= 16'h567c;
        src46 <= 16'h4f00;
        src47 <= 16'hc3e4;
        src48 <= 16'hc4b0;
        src49 <= 16'h7738;
        src50 <= 16'h939e;
        src51 <= 16'hc091;
        src52 <= 16'hbff;
        src53 <= 16'h5201;
        src54 <= 16'hb672;
        src55 <= 16'h7035;
        src56 <= 16'hfe57;
        src57 <= 16'h2477;
        src58 <= 16'h2973;
        src59 <= 16'h9cab;
        src60 <= 16'h11d3;
        src61 <= 16'hd9a;
        src62 <= 16'h1f8;
        src63 <= 16'h8b6b;
        src64 <= 16'hab34;
        src65 <= 16'h33b3;
        src66 <= 16'h5060;
        src67 <= 16'hd1a7;
        src68 <= 16'h97c7;
        src69 <= 16'h450f;
        src70 <= 16'hf6c6;
        src71 <= 16'h7e42;
        src72 <= 16'ha2a8;
        src73 <= 16'h85db;
        src74 <= 16'h9471;
        src75 <= 16'hb198;
        src76 <= 16'hf963;
        src77 <= 16'h3940;
        src78 <= 16'hec79;
        src79 <= 16'h5864;
        src80 <= 16'h4f86;
        src81 <= 16'h2431;
        src82 <= 16'h613f;
        src83 <= 16'h6b24;
        src84 <= 16'hf66;
        src85 <= 16'he98f;
        src86 <= 16'h7962;
        src87 <= 16'h63d6;
        src88 <= 16'h777a;
        src89 <= 16'ha036;
        src90 <= 16'hd5d4;
        src91 <= 16'h6e11;
        src92 <= 16'h81e;
        src93 <= 16'ha0e;
        src94 <= 16'h4f6c;
        src95 <= 16'h8b82;
        src96 <= 16'h575f;
        src97 <= 16'heebd;
        src98 <= 16'h2443;
        src99 <= 16'he606;
        src100 <= 16'hd7c8;
        src101 <= 16'hefb6;
        src102 <= 16'hb891;
        src103 <= 16'hf818;
        src104 <= 16'h639d;
        src105 <= 16'hb171;
        src106 <= 16'h950a;
        src107 <= 16'h1161;
        src108 <= 16'hc5e7;
        src109 <= 16'hf0ef;
        src110 <= 16'h7767;
        src111 <= 16'h5afe;
        src112 <= 16'h8930;
        src113 <= 16'hc7ad;
        src114 <= 16'hc2af;
        src115 <= 16'h5ac4;
        src116 <= 16'hdd8c;
        src117 <= 16'hda8d;
        src118 <= 16'h1f7d;
        src119 <= 16'h4924;
        src120 <= 16'hbc29;
        src121 <= 16'h7432;
        src122 <= 16'h5cbc;
        src123 <= 16'h9453;
        src124 <= 16'h2703;
        src125 <= 16'h7d79;
        src126 <= 16'h8c56;
        src127 <= 16'hb58;
        src128 <= 16'hd1a9;
        src129 <= 16'hda18;
        src130 <= 16'h1f06;
        src131 <= 16'hb7c7;
        src132 <= 16'h13de;
        src133 <= 16'h99d7;
        src134 <= 16'hc44e;
        src135 <= 16'h5fc3;
        src136 <= 16'h3de;
        src137 <= 16'h43fc;
        src138 <= 16'h2ebf;
        src139 <= 16'h82c4;
        src140 <= 16'h72fa;
        src141 <= 16'hbf75;
        src142 <= 16'h2276;
        src143 <= 16'h84b3;
        src144 <= 16'h223e;
        src145 <= 16'h7e8f;
        src146 <= 16'h4cbc;
        src147 <= 16'h5b8a;
        src148 <= 16'h589c;
        src149 <= 16'h2e0a;
        src150 <= 16'h2ae0;
        src151 <= 16'h14da;
        src152 <= 16'he1f2;
        src153 <= 16'h3621;
        src154 <= 16'hce88;
        src155 <= 16'he10e;
        src156 <= 16'hfa7e;
        src157 <= 16'h1869;
        src158 <= 16'h66d5;
        src159 <= 16'ha8e3;
        src160 <= 16'hfd80;
        src161 <= 16'hcb1c;
        exp <= 24'h4e3e7a;
        #1
        src0 <= 16'h9a85;
        src1 <= 16'hba42;
        src2 <= 16'h6a88;
        src3 <= 16'h6d74;
        src4 <= 16'hc6af;
        src5 <= 16'h439b;
        src6 <= 16'h57ce;
        src7 <= 16'h6fec;
        src8 <= 16'hd8f2;
        src9 <= 16'h31f3;
        src10 <= 16'h5229;
        src11 <= 16'hc1cf;
        src12 <= 16'hd437;
        src13 <= 16'h1c96;
        src14 <= 16'h153e;
        src15 <= 16'haad9;
        src16 <= 16'he0e9;
        src17 <= 16'ha362;
        src18 <= 16'he1b0;
        src19 <= 16'hc96e;
        src20 <= 16'haa99;
        src21 <= 16'h536e;
        src22 <= 16'hbeb6;
        src23 <= 16'hdf9;
        src24 <= 16'hd34;
        src25 <= 16'hc6cd;
        src26 <= 16'hc8d9;
        src27 <= 16'ha33;
        src28 <= 16'h987a;
        src29 <= 16'h3826;
        src30 <= 16'hd9ae;
        src31 <= 16'h7f8f;
        src32 <= 16'h6609;
        src33 <= 16'h701f;
        src34 <= 16'h350b;
        src35 <= 16'h5a02;
        src36 <= 16'hba13;
        src37 <= 16'hd132;
        src38 <= 16'h5e9;
        src39 <= 16'ha500;
        src40 <= 16'h7a31;
        src41 <= 16'h9b8b;
        src42 <= 16'heecb;
        src43 <= 16'h3446;
        src44 <= 16'h9a41;
        src45 <= 16'h2caa;
        src46 <= 16'h9ba;
        src47 <= 16'ha33a;
        src48 <= 16'h418b;
        src49 <= 16'h279a;
        src50 <= 16'h815f;
        src51 <= 16'ha9d3;
        src52 <= 16'hfb18;
        src53 <= 16'h512a;
        src54 <= 16'he5b8;
        src55 <= 16'hfd0b;
        src56 <= 16'hba8c;
        src57 <= 16'h88ca;
        src58 <= 16'hd39d;
        src59 <= 16'hff31;
        src60 <= 16'h54b1;
        src61 <= 16'h2968;
        src62 <= 16'h4ab;
        src63 <= 16'h62e7;
        src64 <= 16'hd887;
        src65 <= 16'h4d84;
        src66 <= 16'h796f;
        src67 <= 16'h2e5;
        src68 <= 16'hbfaf;
        src69 <= 16'h3d3a;
        src70 <= 16'hb10e;
        src71 <= 16'h5e6b;
        src72 <= 16'h7e;
        src73 <= 16'h9604;
        src74 <= 16'h9d95;
        src75 <= 16'he7b6;
        src76 <= 16'hb672;
        src77 <= 16'hac9a;
        src78 <= 16'hcab4;
        src79 <= 16'h4ce6;
        src80 <= 16'hb4c1;
        src81 <= 16'h927a;
        src82 <= 16'h431f;
        src83 <= 16'hb1f9;
        src84 <= 16'hb687;
        src85 <= 16'h53a0;
        src86 <= 16'hcd0;
        src87 <= 16'h93fe;
        src88 <= 16'he93e;
        src89 <= 16'h34ea;
        src90 <= 16'hcdca;
        src91 <= 16'h233f;
        src92 <= 16'h4451;
        src93 <= 16'h56fa;
        src94 <= 16'hc1b5;
        src95 <= 16'h7c60;
        src96 <= 16'hd5fc;
        src97 <= 16'h241f;
        src98 <= 16'h5436;
        src99 <= 16'h8d31;
        src100 <= 16'h5672;
        src101 <= 16'hef37;
        src102 <= 16'h9820;
        src103 <= 16'h1118;
        src104 <= 16'h41de;
        src105 <= 16'h60ac;
        src106 <= 16'h14f7;
        src107 <= 16'hf191;
        src108 <= 16'h5bf;
        src109 <= 16'h6ed6;
        src110 <= 16'ha513;
        src111 <= 16'h56a9;
        src112 <= 16'h8165;
        src113 <= 16'h712e;
        src114 <= 16'h7572;
        src115 <= 16'hcc2c;
        src116 <= 16'h5012;
        src117 <= 16'hcac7;
        src118 <= 16'hbbd4;
        src119 <= 16'h2a05;
        src120 <= 16'h8ddf;
        src121 <= 16'hd603;
        src122 <= 16'h211e;
        src123 <= 16'h2a85;
        src124 <= 16'haa3c;
        src125 <= 16'h38ce;
        src126 <= 16'h2b0;
        src127 <= 16'hb84;
        src128 <= 16'h722b;
        src129 <= 16'h7f2a;
        src130 <= 16'hf5f4;
        src131 <= 16'h88d1;
        src132 <= 16'hf89d;
        src133 <= 16'hac6d;
        src134 <= 16'hd75;
        src135 <= 16'h5750;
        src136 <= 16'h3e9b;
        src137 <= 16'h9cc5;
        src138 <= 16'hb789;
        src139 <= 16'h9262;
        src140 <= 16'h5f2a;
        src141 <= 16'ha201;
        src142 <= 16'h83fc;
        src143 <= 16'hfabb;
        src144 <= 16'he3c2;
        src145 <= 16'h8232;
        src146 <= 16'hac1f;
        src147 <= 16'h5904;
        src148 <= 16'hb1fa;
        src149 <= 16'h9b13;
        src150 <= 16'h1a5;
        src151 <= 16'h4986;
        src152 <= 16'h2dde;
        src153 <= 16'h4e8a;
        src154 <= 16'hf864;
        src155 <= 16'ha339;
        src156 <= 16'h6ee3;
        src157 <= 16'h4ec4;
        src158 <= 16'hd152;
        src159 <= 16'h79ce;
        src160 <= 16'h346e;
        src161 <= 16'h89de;
        exp <= 24'h5070c1;
        #1
        src0 <= 16'hd3f2;
        src1 <= 16'hdc1c;
        src2 <= 16'h93c;
        src3 <= 16'h6a18;
        src4 <= 16'h9e01;
        src5 <= 16'hf90c;
        src6 <= 16'h6a36;
        src7 <= 16'h41e1;
        src8 <= 16'ha5c1;
        src9 <= 16'hdd39;
        src10 <= 16'h993e;
        src11 <= 16'ha672;
        src12 <= 16'hc50f;
        src13 <= 16'h592a;
        src14 <= 16'ha118;
        src15 <= 16'hfc70;
        src16 <= 16'h8c69;
        src17 <= 16'hcfe7;
        src18 <= 16'hb925;
        src19 <= 16'hcb7a;
        src20 <= 16'h9c2c;
        src21 <= 16'hae54;
        src22 <= 16'h7cc2;
        src23 <= 16'h78ab;
        src24 <= 16'h3e4e;
        src25 <= 16'h524c;
        src26 <= 16'he450;
        src27 <= 16'h2e39;
        src28 <= 16'hd489;
        src29 <= 16'h4faa;
        src30 <= 16'h42d6;
        src31 <= 16'hd77f;
        src32 <= 16'h7727;
        src33 <= 16'h9c63;
        src34 <= 16'hb1ef;
        src35 <= 16'h293e;
        src36 <= 16'hd6b6;
        src37 <= 16'h7535;
        src38 <= 16'h8774;
        src39 <= 16'h4149;
        src40 <= 16'h8e2a;
        src41 <= 16'hc442;
        src42 <= 16'hf4e4;
        src43 <= 16'hc638;
        src44 <= 16'h84a;
        src45 <= 16'h6993;
        src46 <= 16'h9f3f;
        src47 <= 16'h7c9b;
        src48 <= 16'h736c;
        src49 <= 16'h69ca;
        src50 <= 16'haa97;
        src51 <= 16'h31b;
        src52 <= 16'h4153;
        src53 <= 16'he23c;
        src54 <= 16'hb594;
        src55 <= 16'h9d41;
        src56 <= 16'he1a7;
        src57 <= 16'hee3f;
        src58 <= 16'h7811;
        src59 <= 16'ha398;
        src60 <= 16'h4564;
        src61 <= 16'h9ffe;
        src62 <= 16'h3672;
        src63 <= 16'h8500;
        src64 <= 16'h7848;
        src65 <= 16'h84e;
        src66 <= 16'h7fca;
        src67 <= 16'h7152;
        src68 <= 16'ha3a;
        src69 <= 16'hd054;
        src70 <= 16'h3d9;
        src71 <= 16'h720f;
        src72 <= 16'h770c;
        src73 <= 16'h9719;
        src74 <= 16'hb92;
        src75 <= 16'hf3c0;
        src76 <= 16'hba5d;
        src77 <= 16'h18ab;
        src78 <= 16'h74ab;
        src79 <= 16'hc24a;
        src80 <= 16'hb3;
        src81 <= 16'h1f9f;
        src82 <= 16'h4b4;
        src83 <= 16'hf998;
        src84 <= 16'h9510;
        src85 <= 16'h3c76;
        src86 <= 16'he7c6;
        src87 <= 16'hfd03;
        src88 <= 16'h3ed9;
        src89 <= 16'h9b08;
        src90 <= 16'h4ab7;
        src91 <= 16'hd8c4;
        src92 <= 16'h9422;
        src93 <= 16'hd3c5;
        src94 <= 16'hb8f7;
        src95 <= 16'hf15c;
        src96 <= 16'heec3;
        src97 <= 16'hf3e4;
        src98 <= 16'hd0ed;
        src99 <= 16'h74fe;
        src100 <= 16'ha133;
        src101 <= 16'h896c;
        src102 <= 16'hf669;
        src103 <= 16'h8179;
        src104 <= 16'h3701;
        src105 <= 16'hd563;
        src106 <= 16'h2451;
        src107 <= 16'h3ab6;
        src108 <= 16'hb0b4;
        src109 <= 16'hc71c;
        src110 <= 16'h68d1;
        src111 <= 16'ha6ee;
        src112 <= 16'h53ab;
        src113 <= 16'h514b;
        src114 <= 16'h4c19;
        src115 <= 16'heea4;
        src116 <= 16'h46d7;
        src117 <= 16'h7e55;
        src118 <= 16'hb98d;
        src119 <= 16'h859;
        src120 <= 16'h4a4a;
        src121 <= 16'hd95b;
        src122 <= 16'h2496;
        src123 <= 16'h1e3b;
        src124 <= 16'h27e8;
        src125 <= 16'hd411;
        src126 <= 16'h8e53;
        src127 <= 16'h5afa;
        src128 <= 16'h42cc;
        src129 <= 16'hc3fb;
        src130 <= 16'h656;
        src131 <= 16'h5ef9;
        src132 <= 16'hc464;
        src133 <= 16'hef7e;
        src134 <= 16'h3306;
        src135 <= 16'h65e2;
        src136 <= 16'hc928;
        src137 <= 16'h7f04;
        src138 <= 16'h1d4a;
        src139 <= 16'hbf9b;
        src140 <= 16'h876f;
        src141 <= 16'h8ae6;
        src142 <= 16'h2193;
        src143 <= 16'hbfdb;
        src144 <= 16'h4e7e;
        src145 <= 16'h84b5;
        src146 <= 16'h5be8;
        src147 <= 16'h9277;
        src148 <= 16'h9dfe;
        src149 <= 16'hdc25;
        src150 <= 16'hafd6;
        src151 <= 16'hb8c3;
        src152 <= 16'had0c;
        src153 <= 16'hd7a2;
        src154 <= 16'h6a31;
        src155 <= 16'hebc1;
        src156 <= 16'h7ab3;
        src157 <= 16'haa1e;
        src158 <= 16'h9996;
        src159 <= 16'hc529;
        src160 <= 16'h6e9f;
        src161 <= 16'h3568;
        exp <= 24'h56baab;
        #1
        src0 <= 16'h4779;
        src1 <= 16'h4a5f;
        src2 <= 16'h523f;
        src3 <= 16'h5c4e;
        src4 <= 16'hfe74;
        src5 <= 16'hdeba;
        src6 <= 16'h2614;
        src7 <= 16'hc4a6;
        src8 <= 16'h24f7;
        src9 <= 16'h9fa8;
        src10 <= 16'h1f4a;
        src11 <= 16'h83ba;
        src12 <= 16'hd4f5;
        src13 <= 16'h5596;
        src14 <= 16'hfc8a;
        src15 <= 16'h501c;
        src16 <= 16'h9045;
        src17 <= 16'h4ecf;
        src18 <= 16'ha3a4;
        src19 <= 16'hb707;
        src20 <= 16'h9eb8;
        src21 <= 16'h4cd;
        src22 <= 16'h2ca7;
        src23 <= 16'hcc20;
        src24 <= 16'h6f74;
        src25 <= 16'h2a4e;
        src26 <= 16'h8d86;
        src27 <= 16'h4f89;
        src28 <= 16'h272;
        src29 <= 16'hfa51;
        src30 <= 16'h8ac3;
        src31 <= 16'he315;
        src32 <= 16'h20e8;
        src33 <= 16'h7402;
        src34 <= 16'h4a22;
        src35 <= 16'h9769;
        src36 <= 16'h4246;
        src37 <= 16'he4d;
        src38 <= 16'h65f;
        src39 <= 16'h68e;
        src40 <= 16'hb072;
        src41 <= 16'he8f4;
        src42 <= 16'h8cda;
        src43 <= 16'h441a;
        src44 <= 16'h3746;
        src45 <= 16'he4be;
        src46 <= 16'hb4d9;
        src47 <= 16'hcb18;
        src48 <= 16'h2da0;
        src49 <= 16'hee90;
        src50 <= 16'h4a56;
        src51 <= 16'hb87b;
        src52 <= 16'h64da;
        src53 <= 16'hff5d;
        src54 <= 16'hb388;
        src55 <= 16'h6263;
        src56 <= 16'hd5ca;
        src57 <= 16'h66aa;
        src58 <= 16'h7125;
        src59 <= 16'h6464;
        src60 <= 16'h8ef5;
        src61 <= 16'hb4c;
        src62 <= 16'h52cb;
        src63 <= 16'h761d;
        src64 <= 16'h5507;
        src65 <= 16'h6b17;
        src66 <= 16'h2dce;
        src67 <= 16'habeb;
        src68 <= 16'h2d39;
        src69 <= 16'hf798;
        src70 <= 16'h499d;
        src71 <= 16'hb152;
        src72 <= 16'h64e2;
        src73 <= 16'h9dfa;
        src74 <= 16'h6568;
        src75 <= 16'h180;
        src76 <= 16'heee9;
        src77 <= 16'hefe1;
        src78 <= 16'hc41e;
        src79 <= 16'h4cc0;
        src80 <= 16'h1122;
        src81 <= 16'hf34e;
        src82 <= 16'h5d78;
        src83 <= 16'hcfa9;
        src84 <= 16'he6b2;
        src85 <= 16'hc989;
        src86 <= 16'hb1c7;
        src87 <= 16'hfd37;
        src88 <= 16'h29;
        src89 <= 16'h644;
        src90 <= 16'h2ea;
        src91 <= 16'h6768;
        src92 <= 16'h46c2;
        src93 <= 16'h74bc;
        src94 <= 16'h289c;
        src95 <= 16'he8df;
        src96 <= 16'h7936;
        src97 <= 16'hd43e;
        src98 <= 16'h888a;
        src99 <= 16'ha652;
        src100 <= 16'hb644;
        src101 <= 16'h92a8;
        src102 <= 16'h2be9;
        src103 <= 16'h9911;
        src104 <= 16'h853c;
        src105 <= 16'hef3;
        src106 <= 16'h8c69;
        src107 <= 16'h1132;
        src108 <= 16'ha4ab;
        src109 <= 16'h7afc;
        src110 <= 16'h6ddd;
        src111 <= 16'hfcab;
        src112 <= 16'hf92;
        src113 <= 16'ha230;
        src114 <= 16'hb0da;
        src115 <= 16'hceef;
        src116 <= 16'hbf8c;
        src117 <= 16'h46f8;
        src118 <= 16'h7be0;
        src119 <= 16'h58ac;
        src120 <= 16'hbff9;
        src121 <= 16'h53ba;
        src122 <= 16'h6fe9;
        src123 <= 16'h2649;
        src124 <= 16'h4350;
        src125 <= 16'hc09d;
        src126 <= 16'he84;
        src127 <= 16'hc254;
        src128 <= 16'h1c2a;
        src129 <= 16'h3554;
        src130 <= 16'hf55;
        src131 <= 16'he723;
        src132 <= 16'hd473;
        src133 <= 16'h2643;
        src134 <= 16'hbeb0;
        src135 <= 16'haa56;
        src136 <= 16'hf73d;
        src137 <= 16'hfa2b;
        src138 <= 16'h3efd;
        src139 <= 16'h4dd8;
        src140 <= 16'hdf97;
        src141 <= 16'h6218;
        src142 <= 16'habde;
        src143 <= 16'hf2f6;
        src144 <= 16'h21e3;
        src145 <= 16'hd584;
        src146 <= 16'h3f66;
        src147 <= 16'had21;
        src148 <= 16'hb709;
        src149 <= 16'h5f5;
        src150 <= 16'hae95;
        src151 <= 16'h6ccb;
        src152 <= 16'h169b;
        src153 <= 16'hf53a;
        src154 <= 16'h54d8;
        src155 <= 16'ha2bd;
        src156 <= 16'hee83;
        src157 <= 16'h5cf3;
        src158 <= 16'h5a27;
        src159 <= 16'h9921;
        src160 <= 16'heeb7;
        src161 <= 16'hddc9;
        exp <= 24'h510f84;
        #1
        src0 <= 16'heda1;
        src1 <= 16'hfe6e;
        src2 <= 16'hc224;
        src3 <= 16'h6817;
        src4 <= 16'h5930;
        src5 <= 16'h4688;
        src6 <= 16'h597;
        src7 <= 16'h11f5;
        src8 <= 16'h29e6;
        src9 <= 16'h9cc0;
        src10 <= 16'he248;
        src11 <= 16'h6f8c;
        src12 <= 16'ha3b1;
        src13 <= 16'h6d72;
        src14 <= 16'h68c4;
        src15 <= 16'h8f49;
        src16 <= 16'h66ad;
        src17 <= 16'h2d4c;
        src18 <= 16'hcbc3;
        src19 <= 16'h4977;
        src20 <= 16'hc0b0;
        src21 <= 16'h15f0;
        src22 <= 16'hc8db;
        src23 <= 16'h98ae;
        src24 <= 16'h3e42;
        src25 <= 16'hb6db;
        src26 <= 16'h6250;
        src27 <= 16'h98bf;
        src28 <= 16'h2c32;
        src29 <= 16'h970a;
        src30 <= 16'h3be3;
        src31 <= 16'h94e2;
        src32 <= 16'h9b9e;
        src33 <= 16'h81f0;
        src34 <= 16'hb92e;
        src35 <= 16'h9799;
        src36 <= 16'ha872;
        src37 <= 16'h1339;
        src38 <= 16'h9e18;
        src39 <= 16'h222a;
        src40 <= 16'h2025;
        src41 <= 16'h8bec;
        src42 <= 16'h104d;
        src43 <= 16'haa60;
        src44 <= 16'h682c;
        src45 <= 16'h98d4;
        src46 <= 16'h9d1c;
        src47 <= 16'hf2fe;
        src48 <= 16'h902a;
        src49 <= 16'he588;
        src50 <= 16'h581e;
        src51 <= 16'hdb6f;
        src52 <= 16'h809a;
        src53 <= 16'h3f9e;
        src54 <= 16'hf1dc;
        src55 <= 16'h355f;
        src56 <= 16'h44f6;
        src57 <= 16'h1d46;
        src58 <= 16'h7eb6;
        src59 <= 16'h3e0c;
        src60 <= 16'hc09;
        src61 <= 16'h37f;
        src62 <= 16'hd4da;
        src63 <= 16'h69ec;
        src64 <= 16'hd6b;
        src65 <= 16'hed2d;
        src66 <= 16'h2853;
        src67 <= 16'h8a7a;
        src68 <= 16'h4952;
        src69 <= 16'hf7cd;
        src70 <= 16'h10a4;
        src71 <= 16'h5019;
        src72 <= 16'h8ada;
        src73 <= 16'h93b6;
        src74 <= 16'haf6e;
        src75 <= 16'h106a;
        src76 <= 16'h4e2e;
        src77 <= 16'h4fd;
        src78 <= 16'h72a7;
        src79 <= 16'hfdce;
        src80 <= 16'h2031;
        src81 <= 16'h30a7;
        src82 <= 16'h55a0;
        src83 <= 16'h5f85;
        src84 <= 16'h5118;
        src85 <= 16'h3b70;
        src86 <= 16'hdaf;
        src87 <= 16'h3c8a;
        src88 <= 16'ha499;
        src89 <= 16'hf0d6;
        src90 <= 16'h60c1;
        src91 <= 16'h9959;
        src92 <= 16'h5581;
        src93 <= 16'h69d7;
        src94 <= 16'hf226;
        src95 <= 16'h7f91;
        src96 <= 16'hb139;
        src97 <= 16'h6352;
        src98 <= 16'h24f6;
        src99 <= 16'h7f01;
        src100 <= 16'h35e3;
        src101 <= 16'ha511;
        src102 <= 16'he6c0;
        src103 <= 16'h9f92;
        src104 <= 16'h3082;
        src105 <= 16'ha3f3;
        src106 <= 16'h3b43;
        src107 <= 16'h5f22;
        src108 <= 16'hee53;
        src109 <= 16'h49f;
        src110 <= 16'h705e;
        src111 <= 16'hf8ac;
        src112 <= 16'h259f;
        src113 <= 16'ha4ef;
        src114 <= 16'hdea5;
        src115 <= 16'hb7bf;
        src116 <= 16'hce19;
        src117 <= 16'h49f0;
        src118 <= 16'hc522;
        src119 <= 16'h50d5;
        src120 <= 16'h236f;
        src121 <= 16'h894;
        src122 <= 16'h4e95;
        src123 <= 16'h8837;
        src124 <= 16'hc12d;
        src125 <= 16'h5818;
        src126 <= 16'h480b;
        src127 <= 16'h92a;
        src128 <= 16'h6346;
        src129 <= 16'hec34;
        src130 <= 16'he35a;
        src131 <= 16'h5df5;
        src132 <= 16'hc0bd;
        src133 <= 16'hd8b4;
        src134 <= 16'hc43b;
        src135 <= 16'h52e8;
        src136 <= 16'hf6e0;
        src137 <= 16'hb87b;
        src138 <= 16'hd056;
        src139 <= 16'h7692;
        src140 <= 16'h16d;
        src141 <= 16'hf7b7;
        src142 <= 16'h2f;
        src143 <= 16'h750;
        src144 <= 16'h7b1d;
        src145 <= 16'hf500;
        src146 <= 16'h50e5;
        src147 <= 16'hb900;
        src148 <= 16'hd88d;
        src149 <= 16'h7536;
        src150 <= 16'h4cc5;
        src151 <= 16'hdf96;
        src152 <= 16'h7695;
        src153 <= 16'h8986;
        src154 <= 16'h9e98;
        src155 <= 16'h52d7;
        src156 <= 16'hada5;
        src157 <= 16'h2848;
        src158 <= 16'h8e28;
        src159 <= 16'hb095;
        src160 <= 16'h9803;
        src161 <= 16'hfa25;
        exp <= 24'h4e6910;
        #1
        src0 <= 16'hd3f5;
        src1 <= 16'hedef;
        src2 <= 16'h28e4;
        src3 <= 16'hce9;
        src4 <= 16'hfc87;
        src5 <= 16'hb410;
        src6 <= 16'h938f;
        src7 <= 16'h51c4;
        src8 <= 16'hc19f;
        src9 <= 16'hca77;
        src10 <= 16'h630f;
        src11 <= 16'hcba2;
        src12 <= 16'h32e;
        src13 <= 16'h437f;
        src14 <= 16'h4fb3;
        src15 <= 16'h8eee;
        src16 <= 16'hc74f;
        src17 <= 16'h6c50;
        src18 <= 16'h60ab;
        src19 <= 16'h7587;
        src20 <= 16'h3a8f;
        src21 <= 16'h8835;
        src22 <= 16'h3bad;
        src23 <= 16'h8752;
        src24 <= 16'h5fb0;
        src25 <= 16'h6e48;
        src26 <= 16'hcd12;
        src27 <= 16'hf99d;
        src28 <= 16'h38aa;
        src29 <= 16'h56da;
        src30 <= 16'h5beb;
        src31 <= 16'h634e;
        src32 <= 16'h6800;
        src33 <= 16'h147b;
        src34 <= 16'hd89c;
        src35 <= 16'h86d7;
        src36 <= 16'hea27;
        src37 <= 16'h3925;
        src38 <= 16'h10bf;
        src39 <= 16'ha6be;
        src40 <= 16'h2d74;
        src41 <= 16'h4fca;
        src42 <= 16'he05a;
        src43 <= 16'hc87d;
        src44 <= 16'h56a0;
        src45 <= 16'he74c;
        src46 <= 16'h356d;
        src47 <= 16'h8fa9;
        src48 <= 16'h184c;
        src49 <= 16'ha69e;
        src50 <= 16'hee33;
        src51 <= 16'h3cbc;
        src52 <= 16'h9385;
        src53 <= 16'hac24;
        src54 <= 16'haf1f;
        src55 <= 16'h20e5;
        src56 <= 16'hf3e5;
        src57 <= 16'h175b;
        src58 <= 16'h74df;
        src59 <= 16'h4583;
        src60 <= 16'h2906;
        src61 <= 16'hb4f5;
        src62 <= 16'hbbff;
        src63 <= 16'h115;
        src64 <= 16'hb1f4;
        src65 <= 16'h5754;
        src66 <= 16'he8be;
        src67 <= 16'hd75f;
        src68 <= 16'h42f4;
        src69 <= 16'hff2;
        src70 <= 16'h1356;
        src71 <= 16'hc64f;
        src72 <= 16'h5bbe;
        src73 <= 16'ha465;
        src74 <= 16'h7011;
        src75 <= 16'h3a00;
        src76 <= 16'hf2fb;
        src77 <= 16'hea46;
        src78 <= 16'h2489;
        src79 <= 16'h348c;
        src80 <= 16'hd186;
        src81 <= 16'h9a4f;
        src82 <= 16'hae14;
        src83 <= 16'h9100;
        src84 <= 16'h38b9;
        src85 <= 16'hb3d6;
        src86 <= 16'ha62d;
        src87 <= 16'hdb8e;
        src88 <= 16'hcf29;
        src89 <= 16'hbd8;
        src90 <= 16'h1663;
        src91 <= 16'h2309;
        src92 <= 16'hb308;
        src93 <= 16'he91f;
        src94 <= 16'h67dd;
        src95 <= 16'h7e58;
        src96 <= 16'hf18f;
        src97 <= 16'hfd0a;
        src98 <= 16'h8d19;
        src99 <= 16'h974b;
        src100 <= 16'hd334;
        src101 <= 16'h3cc3;
        src102 <= 16'h5505;
        src103 <= 16'h5bd8;
        src104 <= 16'hc656;
        src105 <= 16'h382e;
        src106 <= 16'h4f23;
        src107 <= 16'h49f3;
        src108 <= 16'he26a;
        src109 <= 16'h4d3b;
        src110 <= 16'hcd70;
        src111 <= 16'h2e4e;
        src112 <= 16'h9511;
        src113 <= 16'h50b2;
        src114 <= 16'h946f;
        src115 <= 16'h1d02;
        src116 <= 16'hb0a;
        src117 <= 16'h3f0c;
        src118 <= 16'hc819;
        src119 <= 16'h484d;
        src120 <= 16'h337b;
        src121 <= 16'h6525;
        src122 <= 16'h4e30;
        src123 <= 16'hbbf8;
        src124 <= 16'ha3c;
        src125 <= 16'hfae6;
        src126 <= 16'h6250;
        src127 <= 16'h9e9e;
        src128 <= 16'h4438;
        src129 <= 16'h4d80;
        src130 <= 16'h688f;
        src131 <= 16'hda68;
        src132 <= 16'h65cf;
        src133 <= 16'hc0e6;
        src134 <= 16'h6bb4;
        src135 <= 16'h9552;
        src136 <= 16'h85b5;
        src137 <= 16'h2f5;
        src138 <= 16'h9a81;
        src139 <= 16'hf28;
        src140 <= 16'h8d7e;
        src141 <= 16'hcf81;
        src142 <= 16'h3493;
        src143 <= 16'h2580;
        src144 <= 16'hee4f;
        src145 <= 16'h3e41;
        src146 <= 16'h2d03;
        src147 <= 16'hdeb1;
        src148 <= 16'h5e5d;
        src149 <= 16'h7a55;
        src150 <= 16'h1c59;
        src151 <= 16'hb8ac;
        src152 <= 16'hd540;
        src153 <= 16'ha490;
        src154 <= 16'he567;
        src155 <= 16'h48a4;
        src156 <= 16'hb7c2;
        src157 <= 16'h95d5;
        src158 <= 16'h8354;
        src159 <= 16'h7355;
        src160 <= 16'h6e49;
        src161 <= 16'h95ca;
        exp <= 24'h4f8e71;
        #1
        src0 <= 16'hd546;
        src1 <= 16'h58e3;
        src2 <= 16'hbe0c;
        src3 <= 16'h7a8f;
        src4 <= 16'hee87;
        src5 <= 16'h9246;
        src6 <= 16'hdba2;
        src7 <= 16'hb48d;
        src8 <= 16'hbf43;
        src9 <= 16'h779c;
        src10 <= 16'h1c28;
        src11 <= 16'h9866;
        src12 <= 16'h5b3a;
        src13 <= 16'h66e5;
        src14 <= 16'h1434;
        src15 <= 16'h6201;
        src16 <= 16'h600e;
        src17 <= 16'h7185;
        src18 <= 16'h5bac;
        src19 <= 16'h60d8;
        src20 <= 16'h26b7;
        src21 <= 16'h9d1f;
        src22 <= 16'hdfde;
        src23 <= 16'he7be;
        src24 <= 16'h8aa7;
        src25 <= 16'hda1f;
        src26 <= 16'h68ea;
        src27 <= 16'hf692;
        src28 <= 16'hf5ad;
        src29 <= 16'hca7;
        src30 <= 16'h2c5c;
        src31 <= 16'h7b40;
        src32 <= 16'ha184;
        src33 <= 16'hbde5;
        src34 <= 16'h5df6;
        src35 <= 16'h8f35;
        src36 <= 16'h2828;
        src37 <= 16'he29a;
        src38 <= 16'hf179;
        src39 <= 16'hed2e;
        src40 <= 16'hf45c;
        src41 <= 16'hdca2;
        src42 <= 16'h6df1;
        src43 <= 16'ha032;
        src44 <= 16'hd6a7;
        src45 <= 16'hcecf;
        src46 <= 16'h54f6;
        src47 <= 16'h147f;
        src48 <= 16'hb16;
        src49 <= 16'h9db8;
        src50 <= 16'h7a8f;
        src51 <= 16'h4c8c;
        src52 <= 16'h409a;
        src53 <= 16'h6424;
        src54 <= 16'hcc63;
        src55 <= 16'h50bc;
        src56 <= 16'hf856;
        src57 <= 16'h5098;
        src58 <= 16'h77df;
        src59 <= 16'hd4b7;
        src60 <= 16'h3d31;
        src61 <= 16'h6399;
        src62 <= 16'h300;
        src63 <= 16'h33b5;
        src64 <= 16'hd8ff;
        src65 <= 16'hfdc7;
        src66 <= 16'hf21c;
        src67 <= 16'hf638;
        src68 <= 16'hb5bd;
        src69 <= 16'h7627;
        src70 <= 16'hf9b;
        src71 <= 16'hb3a4;
        src72 <= 16'hde75;
        src73 <= 16'h6fb7;
        src74 <= 16'hc729;
        src75 <= 16'h5167;
        src76 <= 16'h2608;
        src77 <= 16'he0d0;
        src78 <= 16'hed78;
        src79 <= 16'h300d;
        src80 <= 16'h954a;
        src81 <= 16'ha8c5;
        src82 <= 16'h5937;
        src83 <= 16'h2eff;
        src84 <= 16'hc25;
        src85 <= 16'h9e7e;
        src86 <= 16'ha493;
        src87 <= 16'hefb1;
        src88 <= 16'hbc7c;
        src89 <= 16'ha845;
        src90 <= 16'h802b;
        src91 <= 16'hecf7;
        src92 <= 16'h4e99;
        src93 <= 16'hf6a3;
        src94 <= 16'he125;
        src95 <= 16'he4b9;
        src96 <= 16'hf37f;
        src97 <= 16'h12f;
        src98 <= 16'h263e;
        src99 <= 16'he457;
        src100 <= 16'h3f04;
        src101 <= 16'hf6dd;
        src102 <= 16'h1445;
        src103 <= 16'h1e14;
        src104 <= 16'h16f0;
        src105 <= 16'h151c;
        src106 <= 16'h399f;
        src107 <= 16'h6631;
        src108 <= 16'h71e5;
        src109 <= 16'h5385;
        src110 <= 16'h7e3e;
        src111 <= 16'h382d;
        src112 <= 16'h79b0;
        src113 <= 16'hff8b;
        src114 <= 16'hf244;
        src115 <= 16'h6aa6;
        src116 <= 16'hc24a;
        src117 <= 16'hf729;
        src118 <= 16'h7f7;
        src119 <= 16'hb86f;
        src120 <= 16'hf7c6;
        src121 <= 16'hd186;
        src122 <= 16'hca64;
        src123 <= 16'h9434;
        src124 <= 16'h94d5;
        src125 <= 16'h5c8a;
        src126 <= 16'h6a87;
        src127 <= 16'h69d3;
        src128 <= 16'hc57a;
        src129 <= 16'ha225;
        src130 <= 16'h2e0d;
        src131 <= 16'hb096;
        src132 <= 16'h7900;
        src133 <= 16'h216e;
        src134 <= 16'he8b8;
        src135 <= 16'hf1c2;
        src136 <= 16'hc0af;
        src137 <= 16'hd1bf;
        src138 <= 16'h7f69;
        src139 <= 16'h85c2;
        src140 <= 16'h6952;
        src141 <= 16'h5c72;
        src142 <= 16'h3435;
        src143 <= 16'hdbbf;
        src144 <= 16'hbc43;
        src145 <= 16'h4750;
        src146 <= 16'hf680;
        src147 <= 16'h5e57;
        src148 <= 16'h2efe;
        src149 <= 16'h3997;
        src150 <= 16'h3314;
        src151 <= 16'h55df;
        src152 <= 16'h680f;
        src153 <= 16'hf692;
        src154 <= 16'he9a1;
        src155 <= 16'h2f14;
        src156 <= 16'h34f8;
        src157 <= 16'hfd4e;
        src158 <= 16'ha340;
        src159 <= 16'he7a8;
        src160 <= 16'he591;
        src161 <= 16'h9b96;
        exp <= 24'h59166e;
        #1
        src0 <= 16'h674f;
        src1 <= 16'h1259;
        src2 <= 16'hda4d;
        src3 <= 16'he8a2;
        src4 <= 16'h43e2;
        src5 <= 16'haef6;
        src6 <= 16'hb5a3;
        src7 <= 16'ha98c;
        src8 <= 16'he1f0;
        src9 <= 16'h789b;
        src10 <= 16'hde0b;
        src11 <= 16'haa91;
        src12 <= 16'h8905;
        src13 <= 16'h3b30;
        src14 <= 16'hf80e;
        src15 <= 16'h2646;
        src16 <= 16'h5040;
        src17 <= 16'h331f;
        src18 <= 16'h7229;
        src19 <= 16'h9f6b;
        src20 <= 16'h1073;
        src21 <= 16'h8807;
        src22 <= 16'h7d3b;
        src23 <= 16'h9896;
        src24 <= 16'h7621;
        src25 <= 16'h3f20;
        src26 <= 16'h475a;
        src27 <= 16'hc7a9;
        src28 <= 16'hddd8;
        src29 <= 16'h6ce3;
        src30 <= 16'hd50d;
        src31 <= 16'h6fd3;
        src32 <= 16'hadf1;
        src33 <= 16'hf0;
        src34 <= 16'h2097;
        src35 <= 16'hb43d;
        src36 <= 16'h92eb;
        src37 <= 16'hecce;
        src38 <= 16'h1f5e;
        src39 <= 16'h80ad;
        src40 <= 16'h55e8;
        src41 <= 16'h3985;
        src42 <= 16'h6c38;
        src43 <= 16'h2e50;
        src44 <= 16'hc523;
        src45 <= 16'h6572;
        src46 <= 16'h7074;
        src47 <= 16'h67f8;
        src48 <= 16'h108d;
        src49 <= 16'h151e;
        src50 <= 16'hc520;
        src51 <= 16'h8939;
        src52 <= 16'he5ed;
        src53 <= 16'h9af3;
        src54 <= 16'h3152;
        src55 <= 16'h2877;
        src56 <= 16'h84c6;
        src57 <= 16'hca5f;
        src58 <= 16'hb25;
        src59 <= 16'hcb45;
        src60 <= 16'h3e8a;
        src61 <= 16'hb44b;
        src62 <= 16'hdc13;
        src63 <= 16'h667f;
        src64 <= 16'h854d;
        src65 <= 16'h808b;
        src66 <= 16'hd40f;
        src67 <= 16'h77d5;
        src68 <= 16'h38d3;
        src69 <= 16'h8549;
        src70 <= 16'he670;
        src71 <= 16'hc6fc;
        src72 <= 16'hff11;
        src73 <= 16'ha73d;
        src74 <= 16'h6496;
        src75 <= 16'ha28f;
        src76 <= 16'h6b95;
        src77 <= 16'hd191;
        src78 <= 16'h3099;
        src79 <= 16'h6cc0;
        src80 <= 16'hbcdd;
        src81 <= 16'hc979;
        src82 <= 16'he031;
        src83 <= 16'hf280;
        src84 <= 16'hc001;
        src85 <= 16'hbcc6;
        src86 <= 16'hd4f7;
        src87 <= 16'h1148;
        src88 <= 16'hbee0;
        src89 <= 16'h5d57;
        src90 <= 16'h354d;
        src91 <= 16'h298;
        src92 <= 16'hd8e;
        src93 <= 16'h2ec2;
        src94 <= 16'h9374;
        src95 <= 16'hfef7;
        src96 <= 16'h8908;
        src97 <= 16'ha7c6;
        src98 <= 16'hb043;
        src99 <= 16'h6dfd;
        src100 <= 16'hf22e;
        src101 <= 16'h9fe3;
        src102 <= 16'ha8ee;
        src103 <= 16'h50f2;
        src104 <= 16'ha1d2;
        src105 <= 16'hf7e3;
        src106 <= 16'h8b4c;
        src107 <= 16'h78ee;
        src108 <= 16'hcb3a;
        src109 <= 16'habb8;
        src110 <= 16'h13a8;
        src111 <= 16'hf68c;
        src112 <= 16'h2372;
        src113 <= 16'heea6;
        src114 <= 16'h893b;
        src115 <= 16'h9ae4;
        src116 <= 16'hace4;
        src117 <= 16'h39c0;
        src118 <= 16'h3dc1;
        src119 <= 16'ha25b;
        src120 <= 16'hec7f;
        src121 <= 16'h47c6;
        src122 <= 16'hbd38;
        src123 <= 16'hfc83;
        src124 <= 16'h9624;
        src125 <= 16'h9f7d;
        src126 <= 16'hb60b;
        src127 <= 16'hb4f1;
        src128 <= 16'hadfa;
        src129 <= 16'h259d;
        src130 <= 16'hac3b;
        src131 <= 16'hea21;
        src132 <= 16'hb7b0;
        src133 <= 16'hac7b;
        src134 <= 16'h1aea;
        src135 <= 16'h856a;
        src136 <= 16'h97c8;
        src137 <= 16'h4d31;
        src138 <= 16'h38aa;
        src139 <= 16'h17f8;
        src140 <= 16'hbe5d;
        src141 <= 16'h9ba2;
        src142 <= 16'h1db5;
        src143 <= 16'h2c98;
        src144 <= 16'h1e7f;
        src145 <= 16'hedf0;
        src146 <= 16'h712d;
        src147 <= 16'h9f18;
        src148 <= 16'h4d24;
        src149 <= 16'h6a3f;
        src150 <= 16'h5cce;
        src151 <= 16'h88a8;
        src152 <= 16'hfe3d;
        src153 <= 16'h5c90;
        src154 <= 16'heb42;
        src155 <= 16'h6f06;
        src156 <= 16'haefe;
        src157 <= 16'h4de7;
        src158 <= 16'h962e;
        src159 <= 16'h4edf;
        src160 <= 16'h1575;
        src161 <= 16'h7091;
        exp <= 24'h552e32;
        #1
        src0 <= 16'he1f6;
        src1 <= 16'h8f07;
        src2 <= 16'hded8;
        src3 <= 16'hf1dd;
        src4 <= 16'h577c;
        src5 <= 16'h592d;
        src6 <= 16'h4d89;
        src7 <= 16'hdb8f;
        src8 <= 16'h54aa;
        src9 <= 16'hce87;
        src10 <= 16'h86b4;
        src11 <= 16'h1ce5;
        src12 <= 16'h4fc6;
        src13 <= 16'h5dec;
        src14 <= 16'h4e66;
        src15 <= 16'hf4aa;
        src16 <= 16'h5abd;
        src17 <= 16'h15bb;
        src18 <= 16'h9e60;
        src19 <= 16'hbf1d;
        src20 <= 16'h852e;
        src21 <= 16'h7b48;
        src22 <= 16'h9d07;
        src23 <= 16'hab22;
        src24 <= 16'hfeb;
        src25 <= 16'h44d8;
        src26 <= 16'h269f;
        src27 <= 16'he7d3;
        src28 <= 16'he4b7;
        src29 <= 16'hf47d;
        src30 <= 16'h584f;
        src31 <= 16'h1ed2;
        src32 <= 16'h179a;
        src33 <= 16'h3d19;
        src34 <= 16'hba3b;
        src35 <= 16'hb64e;
        src36 <= 16'hec2e;
        src37 <= 16'hf4a4;
        src38 <= 16'h7d59;
        src39 <= 16'he94c;
        src40 <= 16'h4f8e;
        src41 <= 16'h81b3;
        src42 <= 16'h1587;
        src43 <= 16'h5d32;
        src44 <= 16'he1cc;
        src45 <= 16'h2ef6;
        src46 <= 16'h48f2;
        src47 <= 16'hadb1;
        src48 <= 16'h853b;
        src49 <= 16'h3e30;
        src50 <= 16'h76b1;
        src51 <= 16'hdf0;
        src52 <= 16'hed35;
        src53 <= 16'h5266;
        src54 <= 16'h1256;
        src55 <= 16'h6395;
        src56 <= 16'h83b7;
        src57 <= 16'h9614;
        src58 <= 16'hd67f;
        src59 <= 16'h25fe;
        src60 <= 16'hd81e;
        src61 <= 16'h6321;
        src62 <= 16'h3cfd;
        src63 <= 16'h59ad;
        src64 <= 16'h51da;
        src65 <= 16'hbb8a;
        src66 <= 16'h5cfd;
        src67 <= 16'h8bee;
        src68 <= 16'hf5ed;
        src69 <= 16'hc2fe;
        src70 <= 16'h7971;
        src71 <= 16'h5ca0;
        src72 <= 16'h6da;
        src73 <= 16'h11fe;
        src74 <= 16'h5936;
        src75 <= 16'h7f7d;
        src76 <= 16'h3f53;
        src77 <= 16'h7ff1;
        src78 <= 16'h802;
        src79 <= 16'h76af;
        src80 <= 16'h3c67;
        src81 <= 16'hd447;
        src82 <= 16'hc17d;
        src83 <= 16'hab7e;
        src84 <= 16'h773b;
        src85 <= 16'h93c8;
        src86 <= 16'he951;
        src87 <= 16'h159b;
        src88 <= 16'h7c42;
        src89 <= 16'h39f2;
        src90 <= 16'h532;
        src91 <= 16'h3dc5;
        src92 <= 16'h5af3;
        src93 <= 16'hf50c;
        src94 <= 16'h8b12;
        src95 <= 16'hbe29;
        src96 <= 16'hc77e;
        src97 <= 16'h29d4;
        src98 <= 16'h4f8e;
        src99 <= 16'h48c9;
        src100 <= 16'hb5ef;
        src101 <= 16'h2674;
        src102 <= 16'h20f2;
        src103 <= 16'h7bd3;
        src104 <= 16'h28fa;
        src105 <= 16'hb7f0;
        src106 <= 16'h7700;
        src107 <= 16'hf9f8;
        src108 <= 16'h64db;
        src109 <= 16'hb858;
        src110 <= 16'h8aa9;
        src111 <= 16'h3f40;
        src112 <= 16'h9f36;
        src113 <= 16'h88d1;
        src114 <= 16'h7bad;
        src115 <= 16'hcc99;
        src116 <= 16'h80aa;
        src117 <= 16'h59d6;
        src118 <= 16'h5957;
        src119 <= 16'he3ad;
        src120 <= 16'hfbb;
        src121 <= 16'h7e6a;
        src122 <= 16'h3921;
        src123 <= 16'h923c;
        src124 <= 16'h4b0e;
        src125 <= 16'hab1c;
        src126 <= 16'hfd3;
        src127 <= 16'h6296;
        src128 <= 16'hedfd;
        src129 <= 16'h4e8a;
        src130 <= 16'h53d0;
        src131 <= 16'h7a16;
        src132 <= 16'hef7b;
        src133 <= 16'h7ca6;
        src134 <= 16'hb1f7;
        src135 <= 16'he029;
        src136 <= 16'hfa9e;
        src137 <= 16'heab0;
        src138 <= 16'ha6a2;
        src139 <= 16'hb8b3;
        src140 <= 16'hb757;
        src141 <= 16'h8a3;
        src142 <= 16'h3eb8;
        src143 <= 16'h9435;
        src144 <= 16'hf091;
        src145 <= 16'h5e7b;
        src146 <= 16'hb48c;
        src147 <= 16'h83eb;
        src148 <= 16'h789f;
        src149 <= 16'h9a1b;
        src150 <= 16'h2a3a;
        src151 <= 16'hc52c;
        src152 <= 16'h33d3;
        src153 <= 16'hecfa;
        src154 <= 16'hdb35;
        src155 <= 16'h53c4;
        src156 <= 16'he1de;
        src157 <= 16'hd9e8;
        src158 <= 16'h7564;
        src159 <= 16'he888;
        src160 <= 16'h2783;
        src161 <= 16'hc4a4;
        exp <= 24'h51eee9;
        #1
        src0 <= 16'hd22d;
        src1 <= 16'h2c40;
        src2 <= 16'h4ccf;
        src3 <= 16'hd3b6;
        src4 <= 16'h6591;
        src5 <= 16'hf35e;
        src6 <= 16'hd995;
        src7 <= 16'h7d6d;
        src8 <= 16'h623a;
        src9 <= 16'had8b;
        src10 <= 16'hb50d;
        src11 <= 16'h2d11;
        src12 <= 16'he41b;
        src13 <= 16'hb09f;
        src14 <= 16'h4677;
        src15 <= 16'hd610;
        src16 <= 16'hfc1f;
        src17 <= 16'hf0ed;
        src18 <= 16'h22d4;
        src19 <= 16'hf5b2;
        src20 <= 16'hfad;
        src21 <= 16'h9411;
        src22 <= 16'he44f;
        src23 <= 16'h45c2;
        src24 <= 16'hdbb8;
        src25 <= 16'h6ae1;
        src26 <= 16'h2365;
        src27 <= 16'h589f;
        src28 <= 16'h7b3;
        src29 <= 16'h55ed;
        src30 <= 16'hc489;
        src31 <= 16'hd06b;
        src32 <= 16'ha139;
        src33 <= 16'heab2;
        src34 <= 16'hc97a;
        src35 <= 16'hf0f;
        src36 <= 16'ha0e;
        src37 <= 16'hc74d;
        src38 <= 16'h2ca9;
        src39 <= 16'hde8f;
        src40 <= 16'h4a10;
        src41 <= 16'h6195;
        src42 <= 16'h1d4f;
        src43 <= 16'hd55;
        src44 <= 16'hc913;
        src45 <= 16'h1fb0;
        src46 <= 16'h951;
        src47 <= 16'h2d6c;
        src48 <= 16'h8ece;
        src49 <= 16'hff90;
        src50 <= 16'hbdc9;
        src51 <= 16'h70d1;
        src52 <= 16'hbb07;
        src53 <= 16'had14;
        src54 <= 16'hb5cd;
        src55 <= 16'ha1b;
        src56 <= 16'h9967;
        src57 <= 16'hd23d;
        src58 <= 16'h15e0;
        src59 <= 16'h1f82;
        src60 <= 16'h608c;
        src61 <= 16'h1d9b;
        src62 <= 16'hc8c3;
        src63 <= 16'he0a5;
        src64 <= 16'hde1c;
        src65 <= 16'h2a2c;
        src66 <= 16'hb56e;
        src67 <= 16'h5381;
        src68 <= 16'hf19d;
        src69 <= 16'ha60a;
        src70 <= 16'h7d59;
        src71 <= 16'hd34e;
        src72 <= 16'h3f4b;
        src73 <= 16'h9dd6;
        src74 <= 16'h911e;
        src75 <= 16'h8d67;
        src76 <= 16'h2d6b;
        src77 <= 16'h315e;
        src78 <= 16'haeda;
        src79 <= 16'h9e17;
        src80 <= 16'hcaeb;
        src81 <= 16'h82f6;
        src82 <= 16'h3721;
        src83 <= 16'h2de2;
        src84 <= 16'he03a;
        src85 <= 16'h1eee;
        src86 <= 16'h1a0e;
        src87 <= 16'h42f7;
        src88 <= 16'h5160;
        src89 <= 16'hb1c4;
        src90 <= 16'he08e;
        src91 <= 16'h1b19;
        src92 <= 16'hf04a;
        src93 <= 16'h6503;
        src94 <= 16'h328f;
        src95 <= 16'hb830;
        src96 <= 16'hc02;
        src97 <= 16'h1a05;
        src98 <= 16'h9ccc;
        src99 <= 16'hd55b;
        src100 <= 16'h6f35;
        src101 <= 16'h9f23;
        src102 <= 16'h95f1;
        src103 <= 16'hc523;
        src104 <= 16'ha002;
        src105 <= 16'h986;
        src106 <= 16'h4f0;
        src107 <= 16'hca31;
        src108 <= 16'h872;
        src109 <= 16'h965e;
        src110 <= 16'h2e15;
        src111 <= 16'he732;
        src112 <= 16'h216c;
        src113 <= 16'h5a6b;
        src114 <= 16'h1aad;
        src115 <= 16'h780b;
        src116 <= 16'h5e4b;
        src117 <= 16'h2779;
        src118 <= 16'h6610;
        src119 <= 16'h7b2e;
        src120 <= 16'ha815;
        src121 <= 16'h9ece;
        src122 <= 16'h12b2;
        src123 <= 16'hfda5;
        src124 <= 16'h5af1;
        src125 <= 16'h6e8a;
        src126 <= 16'h679f;
        src127 <= 16'h46e2;
        src128 <= 16'hd810;
        src129 <= 16'h184;
        src130 <= 16'h8a22;
        src131 <= 16'h39df;
        src132 <= 16'h6862;
        src133 <= 16'h4177;
        src134 <= 16'h2a;
        src135 <= 16'h6b8f;
        src136 <= 16'h8c1b;
        src137 <= 16'ha8a8;
        src138 <= 16'h6a76;
        src139 <= 16'h47d3;
        src140 <= 16'h2c6c;
        src141 <= 16'hf985;
        src142 <= 16'h2d73;
        src143 <= 16'hf691;
        src144 <= 16'h3f59;
        src145 <= 16'h7516;
        src146 <= 16'hd9da;
        src147 <= 16'hfc97;
        src148 <= 16'h9027;
        src149 <= 16'h1bf2;
        src150 <= 16'hd195;
        src151 <= 16'h5e79;
        src152 <= 16'h2c7d;
        src153 <= 16'h2bb1;
        src154 <= 16'hdce6;
        src155 <= 16'hca4d;
        src156 <= 16'h50a;
        src157 <= 16'hacc9;
        src158 <= 16'hd8e8;
        src159 <= 16'h4ea5;
        src160 <= 16'h5464;
        src161 <= 16'h2465;
        exp <= 24'h4ddda0;
        #1
        src0 <= 16'h6403;
        src1 <= 16'hd4c;
        src2 <= 16'h80b8;
        src3 <= 16'hcd8b;
        src4 <= 16'ha345;
        src5 <= 16'h9f6a;
        src6 <= 16'hdd5e;
        src7 <= 16'h70d3;
        src8 <= 16'hefc2;
        src9 <= 16'h860c;
        src10 <= 16'h7ac1;
        src11 <= 16'h6006;
        src12 <= 16'hc885;
        src13 <= 16'hb2e0;
        src14 <= 16'hacf4;
        src15 <= 16'h5c7b;
        src16 <= 16'h2fea;
        src17 <= 16'h8847;
        src18 <= 16'h867;
        src19 <= 16'hbbf5;
        src20 <= 16'hea26;
        src21 <= 16'hb0d6;
        src22 <= 16'h4bbb;
        src23 <= 16'h637c;
        src24 <= 16'hb75a;
        src25 <= 16'hbcda;
        src26 <= 16'hb362;
        src27 <= 16'h4d73;
        src28 <= 16'h6110;
        src29 <= 16'h67fa;
        src30 <= 16'h2760;
        src31 <= 16'haa6;
        src32 <= 16'h6581;
        src33 <= 16'h2d5f;
        src34 <= 16'hea23;
        src35 <= 16'hd9ea;
        src36 <= 16'hb685;
        src37 <= 16'h9f9c;
        src38 <= 16'hc160;
        src39 <= 16'hfe59;
        src40 <= 16'h23b6;
        src41 <= 16'h196a;
        src42 <= 16'h2756;
        src43 <= 16'h7662;
        src44 <= 16'h66a6;
        src45 <= 16'h490f;
        src46 <= 16'heed5;
        src47 <= 16'h1705;
        src48 <= 16'hf654;
        src49 <= 16'h677b;
        src50 <= 16'h701d;
        src51 <= 16'ha55a;
        src52 <= 16'he548;
        src53 <= 16'h74ee;
        src54 <= 16'h621f;
        src55 <= 16'hcc5;
        src56 <= 16'hfeaf;
        src57 <= 16'h57a8;
        src58 <= 16'h8597;
        src59 <= 16'h5732;
        src60 <= 16'h2782;
        src61 <= 16'hef52;
        src62 <= 16'he221;
        src63 <= 16'ha4f8;
        src64 <= 16'h6340;
        src65 <= 16'hc5c2;
        src66 <= 16'h6ca9;
        src67 <= 16'h217e;
        src68 <= 16'h6485;
        src69 <= 16'hdf36;
        src70 <= 16'h8aca;
        src71 <= 16'h477d;
        src72 <= 16'h99fe;
        src73 <= 16'h8a6f;
        src74 <= 16'h7c6c;
        src75 <= 16'ha0c0;
        src76 <= 16'hb7e7;
        src77 <= 16'h98dd;
        src78 <= 16'hc2eb;
        src79 <= 16'hf8de;
        src80 <= 16'h78ee;
        src81 <= 16'hce68;
        src82 <= 16'h8182;
        src83 <= 16'hb7c2;
        src84 <= 16'h4476;
        src85 <= 16'h5f65;
        src86 <= 16'h97b;
        src87 <= 16'h454c;
        src88 <= 16'he81f;
        src89 <= 16'hba6f;
        src90 <= 16'he181;
        src91 <= 16'h38e1;
        src92 <= 16'h44e9;
        src93 <= 16'h6e81;
        src94 <= 16'ha440;
        src95 <= 16'hace8;
        src96 <= 16'h64a;
        src97 <= 16'h16f2;
        src98 <= 16'hdac9;
        src99 <= 16'hd931;
        src100 <= 16'h5ceb;
        src101 <= 16'hdc49;
        src102 <= 16'h2129;
        src103 <= 16'h4e0f;
        src104 <= 16'heefb;
        src105 <= 16'h456d;
        src106 <= 16'hc85c;
        src107 <= 16'hce38;
        src108 <= 16'h82aa;
        src109 <= 16'h8a07;
        src110 <= 16'h9214;
        src111 <= 16'hc3ef;
        src112 <= 16'ha430;
        src113 <= 16'h3e6a;
        src114 <= 16'he539;
        src115 <= 16'h201f;
        src116 <= 16'h592f;
        src117 <= 16'h3b94;
        src118 <= 16'hb77f;
        src119 <= 16'hbd54;
        src120 <= 16'h3d1e;
        src121 <= 16'h1a69;
        src122 <= 16'h887a;
        src123 <= 16'h785f;
        src124 <= 16'h9793;
        src125 <= 16'h2303;
        src126 <= 16'h43d0;
        src127 <= 16'h438f;
        src128 <= 16'h1f6d;
        src129 <= 16'hd50;
        src130 <= 16'h8278;
        src131 <= 16'hbf27;
        src132 <= 16'h543c;
        src133 <= 16'hfc83;
        src134 <= 16'hbd37;
        src135 <= 16'h7453;
        src136 <= 16'h50f3;
        src137 <= 16'hb52e;
        src138 <= 16'hcfbe;
        src139 <= 16'hc7c7;
        src140 <= 16'h2e0a;
        src141 <= 16'hb88a;
        src142 <= 16'h60f4;
        src143 <= 16'h99d8;
        src144 <= 16'h5241;
        src145 <= 16'hdadc;
        src146 <= 16'h1a3;
        src147 <= 16'hf2a0;
        src148 <= 16'h78e3;
        src149 <= 16'h4410;
        src150 <= 16'hd695;
        src151 <= 16'ha21;
        src152 <= 16'ha6c7;
        src153 <= 16'h90e3;
        src154 <= 16'he853;
        src155 <= 16'ha26a;
        src156 <= 16'h9c22;
        src157 <= 16'h3894;
        src158 <= 16'h217e;
        src159 <= 16'h1e36;
        src160 <= 16'h7853;
        src161 <= 16'h290c;
        exp <= 24'h529171;
        #1
        src0 <= 16'haac6;
        src1 <= 16'he82b;
        src2 <= 16'hdf;
        src3 <= 16'hf75f;
        src4 <= 16'h3c79;
        src5 <= 16'h6092;
        src6 <= 16'ha0ba;
        src7 <= 16'h824e;
        src8 <= 16'hcb25;
        src9 <= 16'h9692;
        src10 <= 16'hcc71;
        src11 <= 16'hac72;
        src12 <= 16'h15bd;
        src13 <= 16'hf8c1;
        src14 <= 16'h8641;
        src15 <= 16'hcbf9;
        src16 <= 16'hf9da;
        src17 <= 16'h5d3a;
        src18 <= 16'h95a7;
        src19 <= 16'h8850;
        src20 <= 16'hc1c1;
        src21 <= 16'h7a1a;
        src22 <= 16'h43b1;
        src23 <= 16'h7f12;
        src24 <= 16'h1455;
        src25 <= 16'h74a0;
        src26 <= 16'he959;
        src27 <= 16'hd436;
        src28 <= 16'hb6cf;
        src29 <= 16'hefe9;
        src30 <= 16'h21b8;
        src31 <= 16'h9a94;
        src32 <= 16'h505d;
        src33 <= 16'hae47;
        src34 <= 16'ha976;
        src35 <= 16'h2ce3;
        src36 <= 16'hac70;
        src37 <= 16'h35d8;
        src38 <= 16'hdbc7;
        src39 <= 16'hed56;
        src40 <= 16'hef8d;
        src41 <= 16'hd500;
        src42 <= 16'h372c;
        src43 <= 16'h4202;
        src44 <= 16'hf81;
        src45 <= 16'hd397;
        src46 <= 16'h2bda;
        src47 <= 16'hce09;
        src48 <= 16'h61f3;
        src49 <= 16'h1a95;
        src50 <= 16'h588c;
        src51 <= 16'h6eb8;
        src52 <= 16'h63a5;
        src53 <= 16'h6fc7;
        src54 <= 16'h297f;
        src55 <= 16'h9911;
        src56 <= 16'h5e30;
        src57 <= 16'h93f4;
        src58 <= 16'h73d;
        src59 <= 16'h2f9f;
        src60 <= 16'h934e;
        src61 <= 16'h3d79;
        src62 <= 16'hee60;
        src63 <= 16'ha64f;
        src64 <= 16'ha44a;
        src65 <= 16'h8a2e;
        src66 <= 16'h5298;
        src67 <= 16'h19cd;
        src68 <= 16'h37ad;
        src69 <= 16'h4d46;
        src70 <= 16'hc96;
        src71 <= 16'h6837;
        src72 <= 16'hadfe;
        src73 <= 16'h9858;
        src74 <= 16'hda17;
        src75 <= 16'h1ff3;
        src76 <= 16'hebcb;
        src77 <= 16'h2253;
        src78 <= 16'hde64;
        src79 <= 16'h5361;
        src80 <= 16'h491f;
        src81 <= 16'h382a;
        src82 <= 16'hd8f6;
        src83 <= 16'hafe1;
        src84 <= 16'hf76e;
        src85 <= 16'he464;
        src86 <= 16'h9465;
        src87 <= 16'h5997;
        src88 <= 16'ha2e;
        src89 <= 16'he520;
        src90 <= 16'h4ccc;
        src91 <= 16'hfe38;
        src92 <= 16'h2723;
        src93 <= 16'h578c;
        src94 <= 16'h2dc4;
        src95 <= 16'ha012;
        src96 <= 16'h91fd;
        src97 <= 16'he059;
        src98 <= 16'h90b7;
        src99 <= 16'hdc28;
        src100 <= 16'hd545;
        src101 <= 16'h7838;
        src102 <= 16'hed40;
        src103 <= 16'h2937;
        src104 <= 16'h6e1a;
        src105 <= 16'h3118;
        src106 <= 16'h35e4;
        src107 <= 16'h6158;
        src108 <= 16'h115d;
        src109 <= 16'h165;
        src110 <= 16'ha8a9;
        src111 <= 16'h52ec;
        src112 <= 16'hceb6;
        src113 <= 16'hbc0c;
        src114 <= 16'hf6e0;
        src115 <= 16'hd7de;
        src116 <= 16'h787a;
        src117 <= 16'hde14;
        src118 <= 16'h6360;
        src119 <= 16'h3f49;
        src120 <= 16'h865f;
        src121 <= 16'h1ffa;
        src122 <= 16'h40f;
        src123 <= 16'hf0cc;
        src124 <= 16'h259f;
        src125 <= 16'h99d3;
        src126 <= 16'h7d23;
        src127 <= 16'hcef;
        src128 <= 16'h929c;
        src129 <= 16'hd40e;
        src130 <= 16'h9840;
        src131 <= 16'h30ed;
        src132 <= 16'h49b3;
        src133 <= 16'ha0f1;
        src134 <= 16'h5fc3;
        src135 <= 16'hf8f;
        src136 <= 16'hfef7;
        src137 <= 16'hc3af;
        src138 <= 16'hd94e;
        src139 <= 16'hce7f;
        src140 <= 16'h23ad;
        src141 <= 16'h36eb;
        src142 <= 16'he859;
        src143 <= 16'h7dec;
        src144 <= 16'hbce4;
        src145 <= 16'h208a;
        src146 <= 16'hd423;
        src147 <= 16'hc094;
        src148 <= 16'h3a3d;
        src149 <= 16'h158f;
        src150 <= 16'h8bf4;
        src151 <= 16'h2f29;
        src152 <= 16'h1216;
        src153 <= 16'he2bd;
        src154 <= 16'hb8b3;
        src155 <= 16'h5221;
        src156 <= 16'hf168;
        src157 <= 16'h2211;
        src158 <= 16'h608a;
        src159 <= 16'hec9a;
        src160 <= 16'h2998;
        src161 <= 16'h4bf;
        exp <= 24'h5196e3;
        #1
        src0 <= 16'hc368;
        src1 <= 16'hd2d8;
        src2 <= 16'h5b46;
        src3 <= 16'h99e5;
        src4 <= 16'h3255;
        src5 <= 16'h7fea;
        src6 <= 16'h5ad;
        src7 <= 16'h4470;
        src8 <= 16'hbe89;
        src9 <= 16'hcf3f;
        src10 <= 16'haf2b;
        src11 <= 16'h464b;
        src12 <= 16'h80f0;
        src13 <= 16'h9653;
        src14 <= 16'he5f0;
        src15 <= 16'hcd3b;
        src16 <= 16'hd899;
        src17 <= 16'h6482;
        src18 <= 16'h647f;
        src19 <= 16'h2e07;
        src20 <= 16'h7c9f;
        src21 <= 16'h9844;
        src22 <= 16'h616e;
        src23 <= 16'h8d;
        src24 <= 16'h7743;
        src25 <= 16'h6fcd;
        src26 <= 16'h5038;
        src27 <= 16'h6b4;
        src28 <= 16'hd483;
        src29 <= 16'hc7a7;
        src30 <= 16'h989f;
        src31 <= 16'h5331;
        src32 <= 16'haff4;
        src33 <= 16'hf194;
        src34 <= 16'h277f;
        src35 <= 16'h44;
        src36 <= 16'hd1a4;
        src37 <= 16'he3fb;
        src38 <= 16'h338d;
        src39 <= 16'haa1d;
        src40 <= 16'h582;
        src41 <= 16'he058;
        src42 <= 16'h89a8;
        src43 <= 16'hf404;
        src44 <= 16'h5742;
        src45 <= 16'hc810;
        src46 <= 16'hf640;
        src47 <= 16'h721a;
        src48 <= 16'h1168;
        src49 <= 16'h59da;
        src50 <= 16'h73ed;
        src51 <= 16'ha385;
        src52 <= 16'h115e;
        src53 <= 16'h53be;
        src54 <= 16'hbe3f;
        src55 <= 16'h49a0;
        src56 <= 16'hc609;
        src57 <= 16'h8f89;
        src58 <= 16'h436d;
        src59 <= 16'h6d70;
        src60 <= 16'h37f6;
        src61 <= 16'h5758;
        src62 <= 16'h6485;
        src63 <= 16'h1caa;
        src64 <= 16'h7f89;
        src65 <= 16'h9f71;
        src66 <= 16'h317e;
        src67 <= 16'h762c;
        src68 <= 16'hcb8b;
        src69 <= 16'h9998;
        src70 <= 16'h6905;
        src71 <= 16'h1c09;
        src72 <= 16'hd218;
        src73 <= 16'hc839;
        src74 <= 16'h8f97;
        src75 <= 16'hf16;
        src76 <= 16'h12b7;
        src77 <= 16'h986c;
        src78 <= 16'h5316;
        src79 <= 16'hb13e;
        src80 <= 16'h5554;
        src81 <= 16'hc091;
        src82 <= 16'hcb2f;
        src83 <= 16'h1a25;
        src84 <= 16'h3b5e;
        src85 <= 16'hca30;
        src86 <= 16'hfe88;
        src87 <= 16'hc5ad;
        src88 <= 16'h70a7;
        src89 <= 16'h14d3;
        src90 <= 16'h8c4d;
        src91 <= 16'h7d6f;
        src92 <= 16'h2693;
        src93 <= 16'h8e51;
        src94 <= 16'h2ace;
        src95 <= 16'hb5f7;
        src96 <= 16'h3e94;
        src97 <= 16'h4361;
        src98 <= 16'ha38a;
        src99 <= 16'h143;
        src100 <= 16'h60d6;
        src101 <= 16'hc54e;
        src102 <= 16'h5977;
        src103 <= 16'hb144;
        src104 <= 16'h146f;
        src105 <= 16'h6635;
        src106 <= 16'h7449;
        src107 <= 16'h2dad;
        src108 <= 16'hc7f7;
        src109 <= 16'h5715;
        src110 <= 16'h7621;
        src111 <= 16'h465c;
        src112 <= 16'hb1c3;
        src113 <= 16'hbb24;
        src114 <= 16'h369;
        src115 <= 16'h8152;
        src116 <= 16'hceda;
        src117 <= 16'h650b;
        src118 <= 16'hc92c;
        src119 <= 16'h523d;
        src120 <= 16'hd23;
        src121 <= 16'haca7;
        src122 <= 16'h8acf;
        src123 <= 16'hd112;
        src124 <= 16'hbc90;
        src125 <= 16'hb2a5;
        src126 <= 16'h2e1d;
        src127 <= 16'h71e7;
        src128 <= 16'hc079;
        src129 <= 16'ha067;
        src130 <= 16'h4feb;
        src131 <= 16'hc199;
        src132 <= 16'h25ec;
        src133 <= 16'h8316;
        src134 <= 16'he67f;
        src135 <= 16'h6b71;
        src136 <= 16'hc3e8;
        src137 <= 16'hde3;
        src138 <= 16'h756;
        src139 <= 16'hc2b9;
        src140 <= 16'h3b89;
        src141 <= 16'hd86e;
        src142 <= 16'hbf9c;
        src143 <= 16'h53d7;
        src144 <= 16'hbb24;
        src145 <= 16'h2dcc;
        src146 <= 16'hfc0;
        src147 <= 16'h8fe8;
        src148 <= 16'h6feb;
        src149 <= 16'h6f6f;
        src150 <= 16'h6e69;
        src151 <= 16'h806d;
        src152 <= 16'h6326;
        src153 <= 16'h9938;
        src154 <= 16'hbc60;
        src155 <= 16'h92dd;
        src156 <= 16'he413;
        src157 <= 16'h2578;
        src158 <= 16'h7858;
        src159 <= 16'h8697;
        src160 <= 16'he000;
        src161 <= 16'ha487;
        exp <= 24'h4ec904;
        #1
        src0 <= 16'hc80a;
        src1 <= 16'h864f;
        src2 <= 16'h6488;
        src3 <= 16'hb24c;
        src4 <= 16'he0b8;
        src5 <= 16'he550;
        src6 <= 16'ha5a7;
        src7 <= 16'h7644;
        src8 <= 16'hcd6;
        src9 <= 16'he9a7;
        src10 <= 16'hb95b;
        src11 <= 16'h457f;
        src12 <= 16'hc09f;
        src13 <= 16'h1ebe;
        src14 <= 16'h29b2;
        src15 <= 16'hdfc3;
        src16 <= 16'hef5b;
        src17 <= 16'h6a32;
        src18 <= 16'hc658;
        src19 <= 16'h26da;
        src20 <= 16'hd687;
        src21 <= 16'heaf0;
        src22 <= 16'h395b;
        src23 <= 16'h2f3f;
        src24 <= 16'hb31f;
        src25 <= 16'hfd5a;
        src26 <= 16'h60e6;
        src27 <= 16'h5d3d;
        src28 <= 16'h7a29;
        src29 <= 16'h9ca;
        src30 <= 16'he4e8;
        src31 <= 16'he69d;
        src32 <= 16'he6f1;
        src33 <= 16'h744;
        src34 <= 16'hde84;
        src35 <= 16'h1886;
        src36 <= 16'h205c;
        src37 <= 16'hec57;
        src38 <= 16'hc8c7;
        src39 <= 16'ha2fe;
        src40 <= 16'ha0f6;
        src41 <= 16'h529c;
        src42 <= 16'ha89d;
        src43 <= 16'h7616;
        src44 <= 16'h187f;
        src45 <= 16'h21e0;
        src46 <= 16'h76d2;
        src47 <= 16'hb346;
        src48 <= 16'h44a9;
        src49 <= 16'hc31e;
        src50 <= 16'h5dcd;
        src51 <= 16'h6bb4;
        src52 <= 16'h2faa;
        src53 <= 16'hd084;
        src54 <= 16'h9915;
        src55 <= 16'h6493;
        src56 <= 16'h567c;
        src57 <= 16'h5eb8;
        src58 <= 16'h8a27;
        src59 <= 16'h87e9;
        src60 <= 16'h26d6;
        src61 <= 16'h365f;
        src62 <= 16'h6012;
        src63 <= 16'h758b;
        src64 <= 16'h5548;
        src65 <= 16'hbac5;
        src66 <= 16'h8a4b;
        src67 <= 16'h8b;
        src68 <= 16'h1977;
        src69 <= 16'h579c;
        src70 <= 16'h6ac;
        src71 <= 16'hfe1d;
        src72 <= 16'h5007;
        src73 <= 16'h74d7;
        src74 <= 16'h4274;
        src75 <= 16'h4d25;
        src76 <= 16'h403a;
        src77 <= 16'h3704;
        src78 <= 16'h3e25;
        src79 <= 16'h6c3c;
        src80 <= 16'hd74b;
        src81 <= 16'hbcec;
        src82 <= 16'h49af;
        src83 <= 16'hc856;
        src84 <= 16'hb061;
        src85 <= 16'h4cc6;
        src86 <= 16'h7f04;
        src87 <= 16'ha580;
        src88 <= 16'hc60;
        src89 <= 16'hcae6;
        src90 <= 16'h7ac9;
        src91 <= 16'h718b;
        src92 <= 16'hda7d;
        src93 <= 16'h3e15;
        src94 <= 16'h30d0;
        src95 <= 16'h8d55;
        src96 <= 16'h5e5a;
        src97 <= 16'h471a;
        src98 <= 16'hf7a9;
        src99 <= 16'h1b7d;
        src100 <= 16'h3cb8;
        src101 <= 16'h9317;
        src102 <= 16'hb724;
        src103 <= 16'h3a33;
        src104 <= 16'h3863;
        src105 <= 16'hdab0;
        src106 <= 16'h1e2b;
        src107 <= 16'ha2c0;
        src108 <= 16'h72b6;
        src109 <= 16'h7b8e;
        src110 <= 16'h8697;
        src111 <= 16'h1e96;
        src112 <= 16'hdfc7;
        src113 <= 16'h523a;
        src114 <= 16'h203e;
        src115 <= 16'hff24;
        src116 <= 16'hc5db;
        src117 <= 16'he504;
        src118 <= 16'h183c;
        src119 <= 16'ha92d;
        src120 <= 16'h9bea;
        src121 <= 16'h4604;
        src122 <= 16'h7d1f;
        src123 <= 16'h1da3;
        src124 <= 16'h7976;
        src125 <= 16'h154;
        src126 <= 16'h3028;
        src127 <= 16'h8cb8;
        src128 <= 16'hc272;
        src129 <= 16'h185f;
        src130 <= 16'he114;
        src131 <= 16'he97b;
        src132 <= 16'hb4e5;
        src133 <= 16'hda25;
        src134 <= 16'h8f1a;
        src135 <= 16'h8125;
        src136 <= 16'h68be;
        src137 <= 16'h16c0;
        src138 <= 16'h5b34;
        src139 <= 16'h729d;
        src140 <= 16'ha27d;
        src141 <= 16'hf1c6;
        src142 <= 16'h9705;
        src143 <= 16'h9987;
        src144 <= 16'h9cbd;
        src145 <= 16'hf1b7;
        src146 <= 16'hce36;
        src147 <= 16'h87c4;
        src148 <= 16'hf322;
        src149 <= 16'h9cfa;
        src150 <= 16'hdaf7;
        src151 <= 16'h8b70;
        src152 <= 16'he076;
        src153 <= 16'h26fa;
        src154 <= 16'hc8b0;
        src155 <= 16'h1b54;
        src156 <= 16'hf73;
        src157 <= 16'h62bc;
        src158 <= 16'h5513;
        src159 <= 16'h3461;
        src160 <= 16'h8af7;
        src161 <= 16'h5774;
        exp <= 24'h50294f;
        #1
        src0 <= 16'h2eb0;
        src1 <= 16'h996c;
        src2 <= 16'h3cbd;
        src3 <= 16'h89e3;
        src4 <= 16'h76e8;
        src5 <= 16'he9d;
        src6 <= 16'h1ec;
        src7 <= 16'h96a9;
        src8 <= 16'hc4b;
        src9 <= 16'hbf1d;
        src10 <= 16'hb972;
        src11 <= 16'h488f;
        src12 <= 16'h93eb;
        src13 <= 16'h80e;
        src14 <= 16'ha6a3;
        src15 <= 16'h7d20;
        src16 <= 16'hd313;
        src17 <= 16'hf130;
        src18 <= 16'h84cf;
        src19 <= 16'h7556;
        src20 <= 16'h8840;
        src21 <= 16'hb9a9;
        src22 <= 16'h8ae0;
        src23 <= 16'h28ba;
        src24 <= 16'he9d;
        src25 <= 16'h58ab;
        src26 <= 16'h2824;
        src27 <= 16'h2e9b;
        src28 <= 16'h53fc;
        src29 <= 16'h1a67;
        src30 <= 16'hb016;
        src31 <= 16'h73f5;
        src32 <= 16'hfd44;
        src33 <= 16'hf92b;
        src34 <= 16'h542f;
        src35 <= 16'hd9b1;
        src36 <= 16'hdd1d;
        src37 <= 16'h356b;
        src38 <= 16'h6336;
        src39 <= 16'hdf64;
        src40 <= 16'h8482;
        src41 <= 16'hb174;
        src42 <= 16'h5b53;
        src43 <= 16'hc960;
        src44 <= 16'hef63;
        src45 <= 16'h303a;
        src46 <= 16'h4d3c;
        src47 <= 16'h8fbd;
        src48 <= 16'h1964;
        src49 <= 16'hfd29;
        src50 <= 16'hbf53;
        src51 <= 16'h7e07;
        src52 <= 16'h1bcf;
        src53 <= 16'h3c0f;
        src54 <= 16'h5aa2;
        src55 <= 16'he637;
        src56 <= 16'h460b;
        src57 <= 16'h60bc;
        src58 <= 16'h1207;
        src59 <= 16'h9f6c;
        src60 <= 16'hee98;
        src61 <= 16'h9d16;
        src62 <= 16'h31a1;
        src63 <= 16'h2843;
        src64 <= 16'h66dd;
        src65 <= 16'hea2f;
        src66 <= 16'h1534;
        src67 <= 16'hedfa;
        src68 <= 16'h8756;
        src69 <= 16'h1f31;
        src70 <= 16'ha5a4;
        src71 <= 16'hdf8c;
        src72 <= 16'h7c59;
        src73 <= 16'h9a5a;
        src74 <= 16'h5523;
        src75 <= 16'hf2d5;
        src76 <= 16'h782e;
        src77 <= 16'hf8e4;
        src78 <= 16'h77fa;
        src79 <= 16'h48f0;
        src80 <= 16'h8f5d;
        src81 <= 16'hbc5f;
        src82 <= 16'he77f;
        src83 <= 16'hf3cb;
        src84 <= 16'h776f;
        src85 <= 16'hb914;
        src86 <= 16'hf487;
        src87 <= 16'h4d64;
        src88 <= 16'h3cd4;
        src89 <= 16'h8db4;
        src90 <= 16'h1e6c;
        src91 <= 16'hf53f;
        src92 <= 16'hb8a0;
        src93 <= 16'h4067;
        src94 <= 16'h6acd;
        src95 <= 16'h33ac;
        src96 <= 16'hc4d0;
        src97 <= 16'hfea3;
        src98 <= 16'h8323;
        src99 <= 16'hb37b;
        src100 <= 16'h46d;
        src101 <= 16'hdedd;
        src102 <= 16'h96d;
        src103 <= 16'he3fe;
        src104 <= 16'hbb4e;
        src105 <= 16'h7a5a;
        src106 <= 16'h4da0;
        src107 <= 16'he853;
        src108 <= 16'hf43b;
        src109 <= 16'hb67f;
        src110 <= 16'h8109;
        src111 <= 16'h1705;
        src112 <= 16'h3cff;
        src113 <= 16'habff;
        src114 <= 16'h3f90;
        src115 <= 16'hdcc7;
        src116 <= 16'h77b4;
        src117 <= 16'hde5f;
        src118 <= 16'h561d;
        src119 <= 16'h5725;
        src120 <= 16'hf35;
        src121 <= 16'he20d;
        src122 <= 16'hde62;
        src123 <= 16'he2e6;
        src124 <= 16'h4237;
        src125 <= 16'h6fc4;
        src126 <= 16'h6279;
        src127 <= 16'hc792;
        src128 <= 16'hf5af;
        src129 <= 16'h702a;
        src130 <= 16'h21a5;
        src131 <= 16'h6ae6;
        src132 <= 16'h10ee;
        src133 <= 16'hb61d;
        src134 <= 16'hc9d1;
        src135 <= 16'h937;
        src136 <= 16'he8bc;
        src137 <= 16'hf73c;
        src138 <= 16'h525b;
        src139 <= 16'hbfc7;
        src140 <= 16'h1298;
        src141 <= 16'h7bd;
        src142 <= 16'hba41;
        src143 <= 16'h70eb;
        src144 <= 16'h35d1;
        src145 <= 16'hde04;
        src146 <= 16'hce97;
        src147 <= 16'hebe;
        src148 <= 16'h4a3;
        src149 <= 16'h6576;
        src150 <= 16'hfcc5;
        src151 <= 16'hc21a;
        src152 <= 16'h952b;
        src153 <= 16'hc07b;
        src154 <= 16'h474c;
        src155 <= 16'h3e0d;
        src156 <= 16'h579;
        src157 <= 16'hb2a5;
        src158 <= 16'hd1eb;
        src159 <= 16'h35ca;
        src160 <= 16'h826f;
        src161 <= 16'h62ab;
        exp <= 24'h52c7b7;
        #1
        src0 <= 16'h1038;
        src1 <= 16'h7534;
        src2 <= 16'h500f;
        src3 <= 16'hbafe;
        src4 <= 16'h56c4;
        src5 <= 16'h491c;
        src6 <= 16'h73a3;
        src7 <= 16'hf432;
        src8 <= 16'hf0b9;
        src9 <= 16'h3a06;
        src10 <= 16'h3217;
        src11 <= 16'hf93e;
        src12 <= 16'had62;
        src13 <= 16'h7ad3;
        src14 <= 16'h5e92;
        src15 <= 16'hd660;
        src16 <= 16'h1685;
        src17 <= 16'he38a;
        src18 <= 16'ha296;
        src19 <= 16'h2fd9;
        src20 <= 16'h2ae7;
        src21 <= 16'h8b9c;
        src22 <= 16'h21fe;
        src23 <= 16'he2cd;
        src24 <= 16'h3d36;
        src25 <= 16'h9f12;
        src26 <= 16'h609c;
        src27 <= 16'h5758;
        src28 <= 16'h919;
        src29 <= 16'hbcd0;
        src30 <= 16'h5d11;
        src31 <= 16'h5a9;
        src32 <= 16'h2da7;
        src33 <= 16'ha220;
        src34 <= 16'h5014;
        src35 <= 16'h952c;
        src36 <= 16'h93c6;
        src37 <= 16'h5af1;
        src38 <= 16'h6663;
        src39 <= 16'hf868;
        src40 <= 16'h4751;
        src41 <= 16'he11b;
        src42 <= 16'hb0f1;
        src43 <= 16'h67e3;
        src44 <= 16'hf870;
        src45 <= 16'h8239;
        src46 <= 16'h2d41;
        src47 <= 16'hecba;
        src48 <= 16'hb2cc;
        src49 <= 16'had59;
        src50 <= 16'hfb46;
        src51 <= 16'h681c;
        src52 <= 16'h37b6;
        src53 <= 16'h8057;
        src54 <= 16'h689b;
        src55 <= 16'hd5e2;
        src56 <= 16'ha0cf;
        src57 <= 16'h42ee;
        src58 <= 16'hf73a;
        src59 <= 16'hd3dd;
        src60 <= 16'hcd76;
        src61 <= 16'h8d15;
        src62 <= 16'h2947;
        src63 <= 16'h6e1a;
        src64 <= 16'he739;
        src65 <= 16'h9585;
        src66 <= 16'ha17;
        src67 <= 16'hc569;
        src68 <= 16'hafb1;
        src69 <= 16'h5a11;
        src70 <= 16'h71cb;
        src71 <= 16'hb9;
        src72 <= 16'h7e64;
        src73 <= 16'ha035;
        src74 <= 16'h5648;
        src75 <= 16'h9a6c;
        src76 <= 16'hc873;
        src77 <= 16'hb5d8;
        src78 <= 16'h7ab9;
        src79 <= 16'h2eff;
        src80 <= 16'hd6c;
        src81 <= 16'h4bcc;
        src82 <= 16'hdbb1;
        src83 <= 16'h84ba;
        src84 <= 16'h27b3;
        src85 <= 16'hc950;
        src86 <= 16'h1f88;
        src87 <= 16'hd476;
        src88 <= 16'hb181;
        src89 <= 16'h65e9;
        src90 <= 16'h80fe;
        src91 <= 16'hd550;
        src92 <= 16'hd238;
        src93 <= 16'h427f;
        src94 <= 16'h16a9;
        src95 <= 16'h262b;
        src96 <= 16'hf283;
        src97 <= 16'hc5b1;
        src98 <= 16'h553e;
        src99 <= 16'h921e;
        src100 <= 16'h5fbc;
        src101 <= 16'h3eae;
        src102 <= 16'h15d7;
        src103 <= 16'h5daa;
        src104 <= 16'h9c34;
        src105 <= 16'h22fc;
        src106 <= 16'he76c;
        src107 <= 16'h708;
        src108 <= 16'hf816;
        src109 <= 16'h111f;
        src110 <= 16'hc031;
        src111 <= 16'hdb91;
        src112 <= 16'h4a4c;
        src113 <= 16'ha9ba;
        src114 <= 16'h1f47;
        src115 <= 16'hf04;
        src116 <= 16'hf0cc;
        src117 <= 16'ha04;
        src118 <= 16'h5a0a;
        src119 <= 16'hc24d;
        src120 <= 16'h5a05;
        src121 <= 16'h95af;
        src122 <= 16'h6151;
        src123 <= 16'h9f7a;
        src124 <= 16'h9c5c;
        src125 <= 16'h7654;
        src126 <= 16'hb832;
        src127 <= 16'hf154;
        src128 <= 16'h6e00;
        src129 <= 16'hddbe;
        src130 <= 16'ha39;
        src131 <= 16'h9e46;
        src132 <= 16'h9ecf;
        src133 <= 16'h8eb4;
        src134 <= 16'h3c00;
        src135 <= 16'h5c87;
        src136 <= 16'h6c2;
        src137 <= 16'ha614;
        src138 <= 16'h81b3;
        src139 <= 16'h78b7;
        src140 <= 16'hbbc3;
        src141 <= 16'h42a3;
        src142 <= 16'h9629;
        src143 <= 16'hf995;
        src144 <= 16'hd623;
        src145 <= 16'h11d1;
        src146 <= 16'h64c;
        src147 <= 16'h5e73;
        src148 <= 16'h6183;
        src149 <= 16'h249f;
        src150 <= 16'hd73e;
        src151 <= 16'hb2ed;
        src152 <= 16'h2d11;
        src153 <= 16'h39;
        src154 <= 16'hb6d;
        src155 <= 16'ha4a9;
        src156 <= 16'h341c;
        src157 <= 16'h68e5;
        src158 <= 16'hfe11;
        src159 <= 16'hf41;
        src160 <= 16'hc04a;
        src161 <= 16'h3be2;
        exp <= 24'h4edbda;
        #1
        src0 <= 16'h508;
        src1 <= 16'h2df5;
        src2 <= 16'h6979;
        src3 <= 16'h7f95;
        src4 <= 16'hdbfd;
        src5 <= 16'h626b;
        src6 <= 16'haad0;
        src7 <= 16'h1b3d;
        src8 <= 16'h7beb;
        src9 <= 16'h7356;
        src10 <= 16'he3d2;
        src11 <= 16'hc7bb;
        src12 <= 16'h4ad5;
        src13 <= 16'he5ff;
        src14 <= 16'h5f5c;
        src15 <= 16'h36b4;
        src16 <= 16'h7832;
        src17 <= 16'hbaeb;
        src18 <= 16'hfd8;
        src19 <= 16'h9344;
        src20 <= 16'h21b9;
        src21 <= 16'h53c4;
        src22 <= 16'h5514;
        src23 <= 16'h17ed;
        src24 <= 16'h9970;
        src25 <= 16'h8559;
        src26 <= 16'hca62;
        src27 <= 16'h8938;
        src28 <= 16'hada4;
        src29 <= 16'h51d9;
        src30 <= 16'h83e5;
        src31 <= 16'h83aa;
        src32 <= 16'h5333;
        src33 <= 16'h3011;
        src34 <= 16'h9be9;
        src35 <= 16'h41e5;
        src36 <= 16'hb76a;
        src37 <= 16'h3189;
        src38 <= 16'ha058;
        src39 <= 16'h527d;
        src40 <= 16'h9ae6;
        src41 <= 16'hb0a;
        src42 <= 16'he5fb;
        src43 <= 16'h3595;
        src44 <= 16'h3072;
        src45 <= 16'h2a3e;
        src46 <= 16'h825e;
        src47 <= 16'h1a80;
        src48 <= 16'hed32;
        src49 <= 16'hfb26;
        src50 <= 16'hf734;
        src51 <= 16'hcdec;
        src52 <= 16'h5998;
        src53 <= 16'hb91c;
        src54 <= 16'h208;
        src55 <= 16'h89d6;
        src56 <= 16'h22a7;
        src57 <= 16'h8b6d;
        src58 <= 16'h3f39;
        src59 <= 16'h60e3;
        src60 <= 16'hb5fe;
        src61 <= 16'ha4ad;
        src62 <= 16'he50;
        src63 <= 16'h44be;
        src64 <= 16'h4f7c;
        src65 <= 16'h86fa;
        src66 <= 16'h395d;
        src67 <= 16'h1c44;
        src68 <= 16'hce0;
        src69 <= 16'hedc7;
        src70 <= 16'h7a0f;
        src71 <= 16'h1597;
        src72 <= 16'ha478;
        src73 <= 16'hc292;
        src74 <= 16'hcd4f;
        src75 <= 16'h8f1f;
        src76 <= 16'h9393;
        src77 <= 16'h4143;
        src78 <= 16'haf8b;
        src79 <= 16'h86cf;
        src80 <= 16'he5ac;
        src81 <= 16'h2581;
        src82 <= 16'h99cd;
        src83 <= 16'hbf9d;
        src84 <= 16'h7708;
        src85 <= 16'h4ccc;
        src86 <= 16'hfdac;
        src87 <= 16'hb1ae;
        src88 <= 16'h328e;
        src89 <= 16'h47ac;
        src90 <= 16'he8f5;
        src91 <= 16'hb592;
        src92 <= 16'hb0d;
        src93 <= 16'h3ad4;
        src94 <= 16'hf01c;
        src95 <= 16'he2ac;
        src96 <= 16'hc7e5;
        src97 <= 16'h6db5;
        src98 <= 16'h5976;
        src99 <= 16'h89cd;
        src100 <= 16'h2723;
        src101 <= 16'h75d1;
        src102 <= 16'ha31d;
        src103 <= 16'h719c;
        src104 <= 16'h335;
        src105 <= 16'hc503;
        src106 <= 16'h2768;
        src107 <= 16'habeb;
        src108 <= 16'h6959;
        src109 <= 16'hc638;
        src110 <= 16'hc3e2;
        src111 <= 16'h5e54;
        src112 <= 16'ha4c6;
        src113 <= 16'h8966;
        src114 <= 16'haec1;
        src115 <= 16'hea8b;
        src116 <= 16'he718;
        src117 <= 16'h1cd8;
        src118 <= 16'ha059;
        src119 <= 16'h3bf9;
        src120 <= 16'h544d;
        src121 <= 16'h311b;
        src122 <= 16'h13ca;
        src123 <= 16'hf5d6;
        src124 <= 16'hf78d;
        src125 <= 16'h8152;
        src126 <= 16'hb0b5;
        src127 <= 16'hf945;
        src128 <= 16'h8e2d;
        src129 <= 16'hfe1b;
        src130 <= 16'he902;
        src131 <= 16'h4f7b;
        src132 <= 16'h40fa;
        src133 <= 16'h98d9;
        src134 <= 16'hc450;
        src135 <= 16'h5073;
        src136 <= 16'h1f1c;
        src137 <= 16'h3ed8;
        src138 <= 16'h856e;
        src139 <= 16'h8b2f;
        src140 <= 16'hcf67;
        src141 <= 16'h14f7;
        src142 <= 16'h4836;
        src143 <= 16'h8ff2;
        src144 <= 16'h4d7a;
        src145 <= 16'h12e5;
        src146 <= 16'h8ef5;
        src147 <= 16'h7c6d;
        src148 <= 16'he29c;
        src149 <= 16'hb96d;
        src150 <= 16'h2c2c;
        src151 <= 16'h4ba3;
        src152 <= 16'h7959;
        src153 <= 16'h3606;
        src154 <= 16'h4ad3;
        src155 <= 16'h9fbf;
        src156 <= 16'hbdf6;
        src157 <= 16'h7730;
        src158 <= 16'h9283;
        src159 <= 16'h21d;
        src160 <= 16'h97d;
        src161 <= 16'h8d3c;
        exp <= 24'h4dea60;
        #1
        src0 <= 16'h99b1;
        src1 <= 16'h4454;
        src2 <= 16'h827e;
        src3 <= 16'h745e;
        src4 <= 16'h36c9;
        src5 <= 16'h8799;
        src6 <= 16'h11ca;
        src7 <= 16'h20fd;
        src8 <= 16'hec84;
        src9 <= 16'h452f;
        src10 <= 16'h9bc3;
        src11 <= 16'h23c0;
        src12 <= 16'h37d;
        src13 <= 16'hd8c8;
        src14 <= 16'he9b;
        src15 <= 16'h2b23;
        src16 <= 16'h5ce0;
        src17 <= 16'hf5b2;
        src18 <= 16'h4ed7;
        src19 <= 16'h7874;
        src20 <= 16'h86d9;
        src21 <= 16'h11c8;
        src22 <= 16'hf51e;
        src23 <= 16'hbfa2;
        src24 <= 16'h3db0;
        src25 <= 16'h3faa;
        src26 <= 16'hf4ed;
        src27 <= 16'ha72b;
        src28 <= 16'h99b;
        src29 <= 16'h7d41;
        src30 <= 16'h5c1f;
        src31 <= 16'h109f;
        src32 <= 16'h3a0a;
        src33 <= 16'he206;
        src34 <= 16'h36df;
        src35 <= 16'h65bd;
        src36 <= 16'h64d5;
        src37 <= 16'h2cb3;
        src38 <= 16'hb88f;
        src39 <= 16'hb8d8;
        src40 <= 16'ha762;
        src41 <= 16'h63ea;
        src42 <= 16'h695d;
        src43 <= 16'hbec8;
        src44 <= 16'h2335;
        src45 <= 16'h5219;
        src46 <= 16'h2054;
        src47 <= 16'h578;
        src48 <= 16'hb644;
        src49 <= 16'h4388;
        src50 <= 16'h21f6;
        src51 <= 16'h7da5;
        src52 <= 16'h3e01;
        src53 <= 16'he464;
        src54 <= 16'h4f9;
        src55 <= 16'h19e6;
        src56 <= 16'h9d58;
        src57 <= 16'h8c6a;
        src58 <= 16'hef60;
        src59 <= 16'ha37;
        src60 <= 16'h3c08;
        src61 <= 16'hd4e;
        src62 <= 16'h22d0;
        src63 <= 16'ha936;
        src64 <= 16'h291a;
        src65 <= 16'h1d11;
        src66 <= 16'hd83d;
        src67 <= 16'h56a5;
        src68 <= 16'h6cc4;
        src69 <= 16'hbba9;
        src70 <= 16'hbab9;
        src71 <= 16'h556;
        src72 <= 16'h5136;
        src73 <= 16'h4b9b;
        src74 <= 16'h78cd;
        src75 <= 16'h5193;
        src76 <= 16'h3525;
        src77 <= 16'h9a4e;
        src78 <= 16'h6795;
        src79 <= 16'he22b;
        src80 <= 16'h3260;
        src81 <= 16'ha402;
        src82 <= 16'hcdf9;
        src83 <= 16'hcd9f;
        src84 <= 16'h9ec5;
        src85 <= 16'hcbf7;
        src86 <= 16'h6a4f;
        src87 <= 16'hed4b;
        src88 <= 16'h5f9f;
        src89 <= 16'h858a;
        src90 <= 16'hdff6;
        src91 <= 16'h381e;
        src92 <= 16'h6a26;
        src93 <= 16'h6a77;
        src94 <= 16'hf5f2;
        src95 <= 16'hcfe0;
        src96 <= 16'h987e;
        src97 <= 16'hf60;
        src98 <= 16'haaba;
        src99 <= 16'ha097;
        src100 <= 16'h2ccf;
        src101 <= 16'hfdde;
        src102 <= 16'hb561;
        src103 <= 16'he65;
        src104 <= 16'h6bea;
        src105 <= 16'h51be;
        src106 <= 16'h9c8c;
        src107 <= 16'h6c42;
        src108 <= 16'hce86;
        src109 <= 16'hf870;
        src110 <= 16'hb0b8;
        src111 <= 16'hd9b3;
        src112 <= 16'h8e51;
        src113 <= 16'he230;
        src114 <= 16'h536;
        src115 <= 16'h8b39;
        src116 <= 16'he699;
        src117 <= 16'hfd2d;
        src118 <= 16'hd011;
        src119 <= 16'h7c69;
        src120 <= 16'h2a08;
        src121 <= 16'hfb83;
        src122 <= 16'h4207;
        src123 <= 16'h8e0;
        src124 <= 16'h4690;
        src125 <= 16'hb67b;
        src126 <= 16'hdf4d;
        src127 <= 16'he3a5;
        src128 <= 16'hc6c6;
        src129 <= 16'hadd4;
        src130 <= 16'hfd17;
        src131 <= 16'h1c6;
        src132 <= 16'h3002;
        src133 <= 16'hdc49;
        src134 <= 16'h665b;
        src135 <= 16'h9f7c;
        src136 <= 16'h8734;
        src137 <= 16'h51fc;
        src138 <= 16'h5733;
        src139 <= 16'hb43a;
        src140 <= 16'h23b6;
        src141 <= 16'h16e5;
        src142 <= 16'h5355;
        src143 <= 16'hef48;
        src144 <= 16'h16cb;
        src145 <= 16'hba51;
        src146 <= 16'hf798;
        src147 <= 16'h329;
        src148 <= 16'h27e1;
        src149 <= 16'h990;
        src150 <= 16'h7a5d;
        src151 <= 16'h9523;
        src152 <= 16'hea3e;
        src153 <= 16'h302c;
        src154 <= 16'h871a;
        src155 <= 16'h9371;
        src156 <= 16'h85e6;
        src157 <= 16'h87b4;
        src158 <= 16'h5c53;
        src159 <= 16'h9f4f;
        src160 <= 16'h2b6a;
        src161 <= 16'he27b;
        exp <= 24'h4d2466;
        #1
        src0 <= 16'h89dd;
        src1 <= 16'h5d07;
        src2 <= 16'h27d1;
        src3 <= 16'h881;
        src4 <= 16'h7c32;
        src5 <= 16'h9c3e;
        src6 <= 16'ha782;
        src7 <= 16'h3f51;
        src8 <= 16'he10d;
        src9 <= 16'ha0a9;
        src10 <= 16'hcf4e;
        src11 <= 16'ha945;
        src12 <= 16'hac52;
        src13 <= 16'h79e3;
        src14 <= 16'h4a8f;
        src15 <= 16'ha08a;
        src16 <= 16'h4d8c;
        src17 <= 16'h3ca2;
        src18 <= 16'ha2a8;
        src19 <= 16'hbc75;
        src20 <= 16'h1aa9;
        src21 <= 16'hef36;
        src22 <= 16'hbe38;
        src23 <= 16'h917c;
        src24 <= 16'h1bb5;
        src25 <= 16'hfbb4;
        src26 <= 16'h4108;
        src27 <= 16'hd8a8;
        src28 <= 16'h232e;
        src29 <= 16'h3ce4;
        src30 <= 16'ha2af;
        src31 <= 16'h6f77;
        src32 <= 16'hca93;
        src33 <= 16'h6fe2;
        src34 <= 16'hafad;
        src35 <= 16'h6782;
        src36 <= 16'h3f31;
        src37 <= 16'h7ea5;
        src38 <= 16'h1fe0;
        src39 <= 16'h2442;
        src40 <= 16'h8ce9;
        src41 <= 16'h14ac;
        src42 <= 16'hb93b;
        src43 <= 16'hd7e5;
        src44 <= 16'h694c;
        src45 <= 16'h5597;
        src46 <= 16'h2ae1;
        src47 <= 16'h1a8b;
        src48 <= 16'h95ca;
        src49 <= 16'haa43;
        src50 <= 16'h5781;
        src51 <= 16'h72cd;
        src52 <= 16'h3d1e;
        src53 <= 16'h71b7;
        src54 <= 16'he6d0;
        src55 <= 16'h727a;
        src56 <= 16'hc6db;
        src57 <= 16'h3f92;
        src58 <= 16'h2ea9;
        src59 <= 16'hd02;
        src60 <= 16'h7739;
        src61 <= 16'h35e4;
        src62 <= 16'h50b6;
        src63 <= 16'hb71f;
        src64 <= 16'h2b04;
        src65 <= 16'ha8b7;
        src66 <= 16'hf1a5;
        src67 <= 16'h2031;
        src68 <= 16'h660f;
        src69 <= 16'haccd;
        src70 <= 16'h4271;
        src71 <= 16'h159c;
        src72 <= 16'h104c;
        src73 <= 16'hed2;
        src74 <= 16'h3d11;
        src75 <= 16'h6418;
        src76 <= 16'h90ca;
        src77 <= 16'h9053;
        src78 <= 16'h61c9;
        src79 <= 16'h630d;
        src80 <= 16'hcd63;
        src81 <= 16'h7222;
        src82 <= 16'h67d0;
        src83 <= 16'hd653;
        src84 <= 16'hf667;
        src85 <= 16'h3157;
        src86 <= 16'hdd49;
        src87 <= 16'h982;
        src88 <= 16'h11e9;
        src89 <= 16'h6588;
        src90 <= 16'h4ef0;
        src91 <= 16'h4161;
        src92 <= 16'h73c2;
        src93 <= 16'hde21;
        src94 <= 16'h7df5;
        src95 <= 16'h1524;
        src96 <= 16'h6f40;
        src97 <= 16'hc17d;
        src98 <= 16'h273b;
        src99 <= 16'hc548;
        src100 <= 16'h93e4;
        src101 <= 16'h7bbd;
        src102 <= 16'h749f;
        src103 <= 16'h3469;
        src104 <= 16'h86df;
        src105 <= 16'he7db;
        src106 <= 16'hba6e;
        src107 <= 16'h58c9;
        src108 <= 16'h6c5c;
        src109 <= 16'h6ee2;
        src110 <= 16'hf0;
        src111 <= 16'h44cc;
        src112 <= 16'h2e2f;
        src113 <= 16'hbcc2;
        src114 <= 16'h3cfc;
        src115 <= 16'h62e9;
        src116 <= 16'h2ea6;
        src117 <= 16'hac6c;
        src118 <= 16'hcdcb;
        src119 <= 16'h46a0;
        src120 <= 16'h89d4;
        src121 <= 16'hc75c;
        src122 <= 16'hf12c;
        src123 <= 16'hac18;
        src124 <= 16'hb1a0;
        src125 <= 16'hd430;
        src126 <= 16'h7c5c;
        src127 <= 16'h871c;
        src128 <= 16'hf208;
        src129 <= 16'h25;
        src130 <= 16'h68ce;
        src131 <= 16'hed86;
        src132 <= 16'h74f4;
        src133 <= 16'h8088;
        src134 <= 16'h6d38;
        src135 <= 16'hbae0;
        src136 <= 16'hce;
        src137 <= 16'hb60c;
        src138 <= 16'h891b;
        src139 <= 16'he003;
        src140 <= 16'h719b;
        src141 <= 16'h50c5;
        src142 <= 16'h23fe;
        src143 <= 16'ha5b1;
        src144 <= 16'h2058;
        src145 <= 16'h46d1;
        src146 <= 16'h8a60;
        src147 <= 16'h5569;
        src148 <= 16'h70fc;
        src149 <= 16'hb5a8;
        src150 <= 16'h90da;
        src151 <= 16'hab9d;
        src152 <= 16'h9581;
        src153 <= 16'hcd4e;
        src154 <= 16'h881;
        src155 <= 16'h2c49;
        src156 <= 16'h89e;
        src157 <= 16'h1b83;
        src158 <= 16'h6b93;
        src159 <= 16'h6634;
        src160 <= 16'he10b;
        src161 <= 16'h67e6;
        exp <= 24'h4b0984;
        #1
        src0 <= 16'h435b;
        src1 <= 16'h2e6b;
        src2 <= 16'h450;
        src3 <= 16'ha857;
        src4 <= 16'h4bb3;
        src5 <= 16'h7de6;
        src6 <= 16'h7c1b;
        src7 <= 16'he96f;
        src8 <= 16'hebbf;
        src9 <= 16'ha2a1;
        src10 <= 16'ha599;
        src11 <= 16'h53c4;
        src12 <= 16'hb307;
        src13 <= 16'h3e28;
        src14 <= 16'h3d1b;
        src15 <= 16'h42be;
        src16 <= 16'hd8;
        src17 <= 16'he1d7;
        src18 <= 16'hf338;
        src19 <= 16'hf3bd;
        src20 <= 16'h830f;
        src21 <= 16'h59be;
        src22 <= 16'h9e2b;
        src23 <= 16'hcacb;
        src24 <= 16'h88e6;
        src25 <= 16'hc395;
        src26 <= 16'hf97;
        src27 <= 16'hafa8;
        src28 <= 16'hec12;
        src29 <= 16'h6049;
        src30 <= 16'hcd51;
        src31 <= 16'h76ce;
        src32 <= 16'h2f31;
        src33 <= 16'ha546;
        src34 <= 16'h3413;
        src35 <= 16'he5a9;
        src36 <= 16'h694f;
        src37 <= 16'h1e9;
        src38 <= 16'ha298;
        src39 <= 16'h2660;
        src40 <= 16'hc00;
        src41 <= 16'hd806;
        src42 <= 16'h97de;
        src43 <= 16'hdc0e;
        src44 <= 16'hdd70;
        src45 <= 16'h1946;
        src46 <= 16'hba14;
        src47 <= 16'h9060;
        src48 <= 16'h1398;
        src49 <= 16'h9658;
        src50 <= 16'h89e7;
        src51 <= 16'h4239;
        src52 <= 16'he7d6;
        src53 <= 16'hda1b;
        src54 <= 16'h5a4a;
        src55 <= 16'hc886;
        src56 <= 16'h5886;
        src57 <= 16'h2344;
        src58 <= 16'h6916;
        src59 <= 16'h26cd;
        src60 <= 16'hf9f;
        src61 <= 16'h3b5e;
        src62 <= 16'h7507;
        src63 <= 16'h9e53;
        src64 <= 16'h140e;
        src65 <= 16'h2b7e;
        src66 <= 16'ha360;
        src67 <= 16'h6b0a;
        src68 <= 16'hb41;
        src69 <= 16'h194c;
        src70 <= 16'hc622;
        src71 <= 16'h632a;
        src72 <= 16'h9195;
        src73 <= 16'h170a;
        src74 <= 16'hc2d8;
        src75 <= 16'hc05f;
        src76 <= 16'h5a3d;
        src77 <= 16'h8089;
        src78 <= 16'hc431;
        src79 <= 16'hc0f2;
        src80 <= 16'h92d4;
        src81 <= 16'haaa6;
        src82 <= 16'h3243;
        src83 <= 16'hc4ea;
        src84 <= 16'h3ed5;
        src85 <= 16'h5609;
        src86 <= 16'h87bb;
        src87 <= 16'h30d5;
        src88 <= 16'hff9;
        src89 <= 16'h6388;
        src90 <= 16'h3cc1;
        src91 <= 16'h88c2;
        src92 <= 16'hc334;
        src93 <= 16'h6947;
        src94 <= 16'h65d9;
        src95 <= 16'he3e6;
        src96 <= 16'hc193;
        src97 <= 16'hd615;
        src98 <= 16'h7eda;
        src99 <= 16'h8fc2;
        src100 <= 16'hab55;
        src101 <= 16'h67a4;
        src102 <= 16'hca01;
        src103 <= 16'h18c0;
        src104 <= 16'ha777;
        src105 <= 16'hcdb9;
        src106 <= 16'hb06;
        src107 <= 16'hbfde;
        src108 <= 16'h5b38;
        src109 <= 16'hb22c;
        src110 <= 16'h6a01;
        src111 <= 16'hc127;
        src112 <= 16'h4bb2;
        src113 <= 16'hebe8;
        src114 <= 16'h12df;
        src115 <= 16'h4c1b;
        src116 <= 16'heaf4;
        src117 <= 16'h1b0c;
        src118 <= 16'h6dea;
        src119 <= 16'h297c;
        src120 <= 16'hd4d2;
        src121 <= 16'h1513;
        src122 <= 16'hcb02;
        src123 <= 16'ha8b0;
        src124 <= 16'h8c03;
        src125 <= 16'h675;
        src126 <= 16'h3413;
        src127 <= 16'h3672;
        src128 <= 16'hef13;
        src129 <= 16'h8aee;
        src130 <= 16'h4648;
        src131 <= 16'he40a;
        src132 <= 16'h63ee;
        src133 <= 16'h638d;
        src134 <= 16'h862c;
        src135 <= 16'h51e1;
        src136 <= 16'h4409;
        src137 <= 16'h534a;
        src138 <= 16'hb166;
        src139 <= 16'h9f89;
        src140 <= 16'h3135;
        src141 <= 16'h3992;
        src142 <= 16'h2ad6;
        src143 <= 16'hecf5;
        src144 <= 16'he037;
        src145 <= 16'h9a3c;
        src146 <= 16'hf45c;
        src147 <= 16'h73ae;
        src148 <= 16'hceed;
        src149 <= 16'hdada;
        src150 <= 16'h274e;
        src151 <= 16'h3b12;
        src152 <= 16'hd265;
        src153 <= 16'h9749;
        src154 <= 16'hd40b;
        src155 <= 16'hb43a;
        src156 <= 16'he1e6;
        src157 <= 16'h8648;
        src158 <= 16'h5147;
        src159 <= 16'h35a4;
        src160 <= 16'h20a3;
        src161 <= 16'he944;
        exp <= 24'h4ff697;
        #1
        src0 <= 16'h368d;
        src1 <= 16'hb1ae;
        src2 <= 16'h3358;
        src3 <= 16'h37d3;
        src4 <= 16'h58c4;
        src5 <= 16'h54d9;
        src6 <= 16'h7ff7;
        src7 <= 16'h2c7a;
        src8 <= 16'hd8b4;
        src9 <= 16'hb5a9;
        src10 <= 16'h4935;
        src11 <= 16'h9e4d;
        src12 <= 16'h44aa;
        src13 <= 16'h2273;
        src14 <= 16'h5b0b;
        src15 <= 16'hb288;
        src16 <= 16'hee7f;
        src17 <= 16'hf9ec;
        src18 <= 16'had00;
        src19 <= 16'h6e31;
        src20 <= 16'h9917;
        src21 <= 16'h4f0a;
        src22 <= 16'hf59f;
        src23 <= 16'hed12;
        src24 <= 16'hfc84;
        src25 <= 16'h7782;
        src26 <= 16'h11c4;
        src27 <= 16'h98ac;
        src28 <= 16'h6f42;
        src29 <= 16'h4ab7;
        src30 <= 16'h7ff;
        src31 <= 16'h6b36;
        src32 <= 16'h8795;
        src33 <= 16'h35ad;
        src34 <= 16'ha945;
        src35 <= 16'haa9f;
        src36 <= 16'h9e9e;
        src37 <= 16'h41c5;
        src38 <= 16'ha8f7;
        src39 <= 16'h3aac;
        src40 <= 16'h9dce;
        src41 <= 16'h3480;
        src42 <= 16'hda15;
        src43 <= 16'h9502;
        src44 <= 16'h7d16;
        src45 <= 16'he23b;
        src46 <= 16'h76e8;
        src47 <= 16'hf9f0;
        src48 <= 16'hbc78;
        src49 <= 16'h7807;
        src50 <= 16'h2a34;
        src51 <= 16'h23f7;
        src52 <= 16'hd507;
        src53 <= 16'hfe61;
        src54 <= 16'hdbe8;
        src55 <= 16'h984d;
        src56 <= 16'h899a;
        src57 <= 16'h72a4;
        src58 <= 16'h6205;
        src59 <= 16'h708d;
        src60 <= 16'h5541;
        src61 <= 16'h501a;
        src62 <= 16'h7034;
        src63 <= 16'hf766;
        src64 <= 16'h5c60;
        src65 <= 16'hd467;
        src66 <= 16'h7cca;
        src67 <= 16'hf634;
        src68 <= 16'h3d2;
        src69 <= 16'h18ec;
        src70 <= 16'h1a93;
        src71 <= 16'h19ec;
        src72 <= 16'h68f8;
        src73 <= 16'hb5ff;
        src74 <= 16'hfde1;
        src75 <= 16'hf58;
        src76 <= 16'hab6e;
        src77 <= 16'h1356;
        src78 <= 16'h16ca;
        src79 <= 16'hf0c7;
        src80 <= 16'h79f7;
        src81 <= 16'h7ea2;
        src82 <= 16'hdf1b;
        src83 <= 16'h1fc1;
        src84 <= 16'hdfac;
        src85 <= 16'hb42a;
        src86 <= 16'h10e6;
        src87 <= 16'h8999;
        src88 <= 16'ha2d2;
        src89 <= 16'haa85;
        src90 <= 16'h3487;
        src91 <= 16'hdb7;
        src92 <= 16'hdc07;
        src93 <= 16'h6458;
        src94 <= 16'h69e2;
        src95 <= 16'h164d;
        src96 <= 16'h9222;
        src97 <= 16'hc8a7;
        src98 <= 16'hdf6c;
        src99 <= 16'he52f;
        src100 <= 16'h2216;
        src101 <= 16'hdb33;
        src102 <= 16'hfbd5;
        src103 <= 16'hba89;
        src104 <= 16'h1de5;
        src105 <= 16'hc90b;
        src106 <= 16'h657e;
        src107 <= 16'h3a78;
        src108 <= 16'hacf0;
        src109 <= 16'h675d;
        src110 <= 16'h36b6;
        src111 <= 16'hfafa;
        src112 <= 16'hca71;
        src113 <= 16'h88ba;
        src114 <= 16'hd263;
        src115 <= 16'hdfe8;
        src116 <= 16'h6c88;
        src117 <= 16'h5053;
        src118 <= 16'h1cab;
        src119 <= 16'h9826;
        src120 <= 16'hf1c3;
        src121 <= 16'h281f;
        src122 <= 16'h4866;
        src123 <= 16'hfea0;
        src124 <= 16'h361d;
        src125 <= 16'h2a3e;
        src126 <= 16'h8b57;
        src127 <= 16'h51f8;
        src128 <= 16'h7fe0;
        src129 <= 16'h5136;
        src130 <= 16'hf012;
        src131 <= 16'h366d;
        src132 <= 16'h6f42;
        src133 <= 16'h25fc;
        src134 <= 16'h7b2a;
        src135 <= 16'h7ac8;
        src136 <= 16'h8e9;
        src137 <= 16'hef98;
        src138 <= 16'hdece;
        src139 <= 16'h67ce;
        src140 <= 16'hd051;
        src141 <= 16'h964a;
        src142 <= 16'h643d;
        src143 <= 16'h3b77;
        src144 <= 16'h4eb1;
        src145 <= 16'hb316;
        src146 <= 16'h9b79;
        src147 <= 16'hbe58;
        src148 <= 16'hb14;
        src149 <= 16'hf0cb;
        src150 <= 16'h9fa7;
        src151 <= 16'hd67d;
        src152 <= 16'h3b8c;
        src153 <= 16'h3a18;
        src154 <= 16'h50a0;
        src155 <= 16'h1dbf;
        src156 <= 16'hace7;
        src157 <= 16'h7b09;
        src158 <= 16'hf55a;
        src159 <= 16'heb2d;
        src160 <= 16'h41d0;
        src161 <= 16'h7933;
        exp <= 24'h528f3a;
        #1
        src0 <= 16'h62c6;
        src1 <= 16'h6155;
        src2 <= 16'hc65c;
        src3 <= 16'h2785;
        src4 <= 16'hdea;
        src5 <= 16'h337a;
        src6 <= 16'h89d7;
        src7 <= 16'h79a0;
        src8 <= 16'hd12e;
        src9 <= 16'had96;
        src10 <= 16'h2b48;
        src11 <= 16'h7e6b;
        src12 <= 16'he63a;
        src13 <= 16'hbe51;
        src14 <= 16'h1b15;
        src15 <= 16'hb400;
        src16 <= 16'h95fc;
        src17 <= 16'ha4ea;
        src18 <= 16'hc597;
        src19 <= 16'hdfcf;
        src20 <= 16'h7e5c;
        src21 <= 16'h5219;
        src22 <= 16'ha769;
        src23 <= 16'hd513;
        src24 <= 16'h3be1;
        src25 <= 16'h78ec;
        src26 <= 16'h1d30;
        src27 <= 16'h5a9c;
        src28 <= 16'hbc48;
        src29 <= 16'h1fb1;
        src30 <= 16'h4ee;
        src31 <= 16'hdc67;
        src32 <= 16'h9a92;
        src33 <= 16'h156f;
        src34 <= 16'hcfda;
        src35 <= 16'h8f7;
        src36 <= 16'he068;
        src37 <= 16'hac97;
        src38 <= 16'heda6;
        src39 <= 16'h85a3;
        src40 <= 16'hd0d5;
        src41 <= 16'hb96f;
        src42 <= 16'hcea4;
        src43 <= 16'h8762;
        src44 <= 16'hac1f;
        src45 <= 16'h9f89;
        src46 <= 16'h2590;
        src47 <= 16'hcbc7;
        src48 <= 16'hcbf3;
        src49 <= 16'h80bf;
        src50 <= 16'h6b1c;
        src51 <= 16'h8343;
        src52 <= 16'h547b;
        src53 <= 16'hd1b5;
        src54 <= 16'h42a3;
        src55 <= 16'h9e1c;
        src56 <= 16'hffbd;
        src57 <= 16'h2946;
        src58 <= 16'h6230;
        src59 <= 16'hca1e;
        src60 <= 16'h79eb;
        src61 <= 16'h4a0a;
        src62 <= 16'hea91;
        src63 <= 16'h59d0;
        src64 <= 16'h5237;
        src65 <= 16'hedc6;
        src66 <= 16'h3264;
        src67 <= 16'h1c26;
        src68 <= 16'h67e9;
        src69 <= 16'h96c6;
        src70 <= 16'h95b9;
        src71 <= 16'hd387;
        src72 <= 16'h3c04;
        src73 <= 16'hab30;
        src74 <= 16'h22f9;
        src75 <= 16'h1dcf;
        src76 <= 16'h3c53;
        src77 <= 16'ha8b6;
        src78 <= 16'h674c;
        src79 <= 16'h329c;
        src80 <= 16'h8a78;
        src81 <= 16'h3998;
        src82 <= 16'h8819;
        src83 <= 16'h5668;
        src84 <= 16'h91aa;
        src85 <= 16'hfa1b;
        src86 <= 16'h4812;
        src87 <= 16'h3c42;
        src88 <= 16'hae7e;
        src89 <= 16'hdda1;
        src90 <= 16'h91e5;
        src91 <= 16'h6c5f;
        src92 <= 16'hd99d;
        src93 <= 16'hc921;
        src94 <= 16'h8e22;
        src95 <= 16'h669c;
        src96 <= 16'h267f;
        src97 <= 16'hae38;
        src98 <= 16'hab29;
        src99 <= 16'h2da5;
        src100 <= 16'h9a26;
        src101 <= 16'hf47f;
        src102 <= 16'hc807;
        src103 <= 16'h99e2;
        src104 <= 16'h29a7;
        src105 <= 16'he016;
        src106 <= 16'hb27a;
        src107 <= 16'h945f;
        src108 <= 16'hccde;
        src109 <= 16'hbb3b;
        src110 <= 16'h2c14;
        src111 <= 16'h78e2;
        src112 <= 16'h18e2;
        src113 <= 16'h9222;
        src114 <= 16'hddd0;
        src115 <= 16'hb4b1;
        src116 <= 16'h378d;
        src117 <= 16'h765d;
        src118 <= 16'h9396;
        src119 <= 16'hee7b;
        src120 <= 16'ha286;
        src121 <= 16'hdeda;
        src122 <= 16'ha185;
        src123 <= 16'h7349;
        src124 <= 16'hd566;
        src125 <= 16'h8d1a;
        src126 <= 16'hd48c;
        src127 <= 16'h40c6;
        src128 <= 16'he5f6;
        src129 <= 16'hd410;
        src130 <= 16'h50a4;
        src131 <= 16'h4472;
        src132 <= 16'h3050;
        src133 <= 16'h3fd7;
        src134 <= 16'h19d1;
        src135 <= 16'hd085;
        src136 <= 16'h77df;
        src137 <= 16'h311;
        src138 <= 16'h7b1d;
        src139 <= 16'h2b72;
        src140 <= 16'hd848;
        src141 <= 16'ha6e0;
        src142 <= 16'h58;
        src143 <= 16'h7c36;
        src144 <= 16'h168d;
        src145 <= 16'hb1f1;
        src146 <= 16'hbf57;
        src147 <= 16'hb627;
        src148 <= 16'hb131;
        src149 <= 16'h16bc;
        src150 <= 16'h2134;
        src151 <= 16'h9e3a;
        src152 <= 16'hbeb9;
        src153 <= 16'h56bb;
        src154 <= 16'h3997;
        src155 <= 16'h6bf0;
        src156 <= 16'h95aa;
        src157 <= 16'h3d55;
        src158 <= 16'hf30d;
        src159 <= 16'h75f3;
        src160 <= 16'hdd89;
        src161 <= 16'h8685;
        exp <= 24'h53e06d;
        #1
        src0 <= 16'h564c;
        src1 <= 16'hf114;
        src2 <= 16'hbb4;
        src3 <= 16'hafa2;
        src4 <= 16'h7f66;
        src5 <= 16'h2ce0;
        src6 <= 16'hdd86;
        src7 <= 16'h2319;
        src8 <= 16'h3122;
        src9 <= 16'h163c;
        src10 <= 16'hdb3a;
        src11 <= 16'h3b39;
        src12 <= 16'h2099;
        src13 <= 16'h74ef;
        src14 <= 16'hc7c1;
        src15 <= 16'h646b;
        src16 <= 16'hb546;
        src17 <= 16'he940;
        src18 <= 16'h5e6;
        src19 <= 16'hb1a;
        src20 <= 16'hd3b3;
        src21 <= 16'h6eb3;
        src22 <= 16'he313;
        src23 <= 16'ha455;
        src24 <= 16'hc982;
        src25 <= 16'h37a6;
        src26 <= 16'h89bb;
        src27 <= 16'h97b7;
        src28 <= 16'h93f9;
        src29 <= 16'h8dfb;
        src30 <= 16'hb0b6;
        src31 <= 16'h2da5;
        src32 <= 16'h6208;
        src33 <= 16'h896d;
        src34 <= 16'h5f95;
        src35 <= 16'heef5;
        src36 <= 16'he16;
        src37 <= 16'h9075;
        src38 <= 16'h2064;
        src39 <= 16'hcfa6;
        src40 <= 16'h40cc;
        src41 <= 16'h2596;
        src42 <= 16'h9eb0;
        src43 <= 16'hb61b;
        src44 <= 16'h5c1;
        src45 <= 16'h4d5c;
        src46 <= 16'h300d;
        src47 <= 16'h2c7b;
        src48 <= 16'h2f58;
        src49 <= 16'h2c87;
        src50 <= 16'h636a;
        src51 <= 16'h4c84;
        src52 <= 16'hd014;
        src53 <= 16'h195c;
        src54 <= 16'h2b75;
        src55 <= 16'ha5ea;
        src56 <= 16'h9386;
        src57 <= 16'h5aa7;
        src58 <= 16'h2fe2;
        src59 <= 16'hc2d2;
        src60 <= 16'h46b9;
        src61 <= 16'h95d9;
        src62 <= 16'h9d88;
        src63 <= 16'h5173;
        src64 <= 16'hf76d;
        src65 <= 16'hf590;
        src66 <= 16'h8fd0;
        src67 <= 16'h24a1;
        src68 <= 16'ha237;
        src69 <= 16'hefc7;
        src70 <= 16'h565c;
        src71 <= 16'hef22;
        src72 <= 16'h6487;
        src73 <= 16'hef6f;
        src74 <= 16'h50b9;
        src75 <= 16'h67a0;
        src76 <= 16'h13bc;
        src77 <= 16'hefa5;
        src78 <= 16'h982d;
        src79 <= 16'h2154;
        src80 <= 16'hfee3;
        src81 <= 16'hdc0d;
        src82 <= 16'h23b4;
        src83 <= 16'hddc3;
        src84 <= 16'he3e7;
        src85 <= 16'hb0a0;
        src86 <= 16'h5acf;
        src87 <= 16'h63e4;
        src88 <= 16'h831b;
        src89 <= 16'hd24b;
        src90 <= 16'h7e7a;
        src91 <= 16'h214c;
        src92 <= 16'h9d90;
        src93 <= 16'h87ae;
        src94 <= 16'h75fa;
        src95 <= 16'hb0e8;
        src96 <= 16'hf951;
        src97 <= 16'hbf54;
        src98 <= 16'hed0f;
        src99 <= 16'hbea8;
        src100 <= 16'hae11;
        src101 <= 16'hbd25;
        src102 <= 16'hf10a;
        src103 <= 16'h7f43;
        src104 <= 16'h3fb0;
        src105 <= 16'h2b67;
        src106 <= 16'hdb6b;
        src107 <= 16'h540f;
        src108 <= 16'hc1ed;
        src109 <= 16'h1085;
        src110 <= 16'h2f80;
        src111 <= 16'h9dab;
        src112 <= 16'hff4f;
        src113 <= 16'h544b;
        src114 <= 16'h3c46;
        src115 <= 16'h8fef;
        src116 <= 16'h53bb;
        src117 <= 16'h1020;
        src118 <= 16'h6b82;
        src119 <= 16'ha947;
        src120 <= 16'h9195;
        src121 <= 16'h79fe;
        src122 <= 16'hc408;
        src123 <= 16'he4d6;
        src124 <= 16'haef0;
        src125 <= 16'hf938;
        src126 <= 16'h1a91;
        src127 <= 16'h3617;
        src128 <= 16'heb15;
        src129 <= 16'h4b66;
        src130 <= 16'h56ee;
        src131 <= 16'hd2f;
        src132 <= 16'h4107;
        src133 <= 16'h27e8;
        src134 <= 16'h5c11;
        src135 <= 16'hed5;
        src136 <= 16'h45df;
        src137 <= 16'hf23f;
        src138 <= 16'h3ace;
        src139 <= 16'h969e;
        src140 <= 16'hbce7;
        src141 <= 16'h848a;
        src142 <= 16'h990e;
        src143 <= 16'hbf26;
        src144 <= 16'hb772;
        src145 <= 16'he430;
        src146 <= 16'h1fe0;
        src147 <= 16'h8eba;
        src148 <= 16'h5c6d;
        src149 <= 16'hea03;
        src150 <= 16'h9807;
        src151 <= 16'h1364;
        src152 <= 16'hcd6a;
        src153 <= 16'h729d;
        src154 <= 16'h77a4;
        src155 <= 16'h81af;
        src156 <= 16'h19df;
        src157 <= 16'h4a04;
        src158 <= 16'hedb9;
        src159 <= 16'hbd28;
        src160 <= 16'hc978;
        src161 <= 16'h9464;
        exp <= 24'h517843;
        #1
        src0 <= 16'h148;
        src1 <= 16'hb99d;
        src2 <= 16'h2ca7;
        src3 <= 16'hb2ce;
        src4 <= 16'hf5be;
        src5 <= 16'h5c1d;
        src6 <= 16'h3366;
        src7 <= 16'hf43b;
        src8 <= 16'h6528;
        src9 <= 16'hf5c3;
        src10 <= 16'h1cbc;
        src11 <= 16'hbc72;
        src12 <= 16'h96a0;
        src13 <= 16'h8029;
        src14 <= 16'haba3;
        src15 <= 16'hc1d0;
        src16 <= 16'h3a8f;
        src17 <= 16'hae38;
        src18 <= 16'h151;
        src19 <= 16'h1375;
        src20 <= 16'hde2c;
        src21 <= 16'h1c77;
        src22 <= 16'hae85;
        src23 <= 16'h1355;
        src24 <= 16'hb83a;
        src25 <= 16'h4f3e;
        src26 <= 16'hc993;
        src27 <= 16'h7334;
        src28 <= 16'h57ae;
        src29 <= 16'hf45c;
        src30 <= 16'h938c;
        src31 <= 16'hfbd8;
        src32 <= 16'h7c1c;
        src33 <= 16'h1281;
        src34 <= 16'h75d0;
        src35 <= 16'h28fd;
        src36 <= 16'hb91;
        src37 <= 16'h1389;
        src38 <= 16'hb06d;
        src39 <= 16'h3276;
        src40 <= 16'h281f;
        src41 <= 16'h2d34;
        src42 <= 16'h6d4f;
        src43 <= 16'hd898;
        src44 <= 16'h5e23;
        src45 <= 16'h7053;
        src46 <= 16'h17ef;
        src47 <= 16'h9bf9;
        src48 <= 16'h4448;
        src49 <= 16'h6cfe;
        src50 <= 16'hbde1;
        src51 <= 16'h1b5f;
        src52 <= 16'hb0c;
        src53 <= 16'h5933;
        src54 <= 16'h772d;
        src55 <= 16'hef0b;
        src56 <= 16'h8a40;
        src57 <= 16'h570;
        src58 <= 16'h689b;
        src59 <= 16'h5803;
        src60 <= 16'hf2eb;
        src61 <= 16'h304b;
        src62 <= 16'h382a;
        src63 <= 16'h696c;
        src64 <= 16'h6fe9;
        src65 <= 16'h6ccf;
        src66 <= 16'h5b79;
        src67 <= 16'hc2c3;
        src68 <= 16'h24f0;
        src69 <= 16'h99e1;
        src70 <= 16'h2827;
        src71 <= 16'h1d55;
        src72 <= 16'h4fc7;
        src73 <= 16'h8cc9;
        src74 <= 16'h9aa0;
        src75 <= 16'he9ca;
        src76 <= 16'haa28;
        src77 <= 16'h90d2;
        src78 <= 16'hd5bb;
        src79 <= 16'heff8;
        src80 <= 16'hce86;
        src81 <= 16'h1ba9;
        src82 <= 16'h6ce2;
        src83 <= 16'h35ee;
        src84 <= 16'h8cdd;
        src85 <= 16'h450;
        src86 <= 16'h882;
        src87 <= 16'h197;
        src88 <= 16'h69c9;
        src89 <= 16'h5ecc;
        src90 <= 16'h8ffc;
        src91 <= 16'hae63;
        src92 <= 16'h6637;
        src93 <= 16'hebe8;
        src94 <= 16'h520d;
        src95 <= 16'hd4b1;
        src96 <= 16'hae9b;
        src97 <= 16'h82be;
        src98 <= 16'h7b52;
        src99 <= 16'h7893;
        src100 <= 16'h4b6e;
        src101 <= 16'h2303;
        src102 <= 16'h1fd8;
        src103 <= 16'hff6;
        src104 <= 16'h773e;
        src105 <= 16'h8af1;
        src106 <= 16'ha894;
        src107 <= 16'h203d;
        src108 <= 16'h2eb5;
        src109 <= 16'h891e;
        src110 <= 16'hcd3d;
        src111 <= 16'h25a0;
        src112 <= 16'ha789;
        src113 <= 16'h7e8b;
        src114 <= 16'h65e5;
        src115 <= 16'h3990;
        src116 <= 16'ha49c;
        src117 <= 16'h7c95;
        src118 <= 16'h53f7;
        src119 <= 16'ha5c4;
        src120 <= 16'he26a;
        src121 <= 16'ha1cf;
        src122 <= 16'h7760;
        src123 <= 16'h3e43;
        src124 <= 16'h305f;
        src125 <= 16'h6d17;
        src126 <= 16'ha0bd;
        src127 <= 16'hac83;
        src128 <= 16'hec4b;
        src129 <= 16'hc8c8;
        src130 <= 16'h2402;
        src131 <= 16'ha41b;
        src132 <= 16'hb63f;
        src133 <= 16'hda9d;
        src134 <= 16'hd235;
        src135 <= 16'h386c;
        src136 <= 16'h57d0;
        src137 <= 16'hc3e5;
        src138 <= 16'h961a;
        src139 <= 16'h8673;
        src140 <= 16'h4598;
        src141 <= 16'h8be7;
        src142 <= 16'h1841;
        src143 <= 16'he9a4;
        src144 <= 16'h7378;
        src145 <= 16'hf5c4;
        src146 <= 16'h78e0;
        src147 <= 16'he340;
        src148 <= 16'h695;
        src149 <= 16'h51f4;
        src150 <= 16'h5a8c;
        src151 <= 16'h6e33;
        src152 <= 16'h6318;
        src153 <= 16'h2594;
        src154 <= 16'h50f5;
        src155 <= 16'h74f2;
        src156 <= 16'h1e9d;
        src157 <= 16'hff7c;
        src158 <= 16'hf2b5;
        src159 <= 16'h2d8e;
        src160 <= 16'habd5;
        src161 <= 16'hf4ac;
        exp <= 24'h4bdc91;
        #1
        src0 <= 16'h51de;
        src1 <= 16'h761a;
        src2 <= 16'h9acf;
        src3 <= 16'h304c;
        src4 <= 16'ha18f;
        src5 <= 16'h1dbf;
        src6 <= 16'h4281;
        src7 <= 16'h93e6;
        src8 <= 16'h776a;
        src9 <= 16'h2344;
        src10 <= 16'hf579;
        src11 <= 16'h4d07;
        src12 <= 16'hb19c;
        src13 <= 16'h21c8;
        src14 <= 16'h79c5;
        src15 <= 16'h6805;
        src16 <= 16'h3cc5;
        src17 <= 16'hbade;
        src18 <= 16'h9a5b;
        src19 <= 16'hb419;
        src20 <= 16'h82e;
        src21 <= 16'ha967;
        src22 <= 16'hf0dd;
        src23 <= 16'hb1ad;
        src24 <= 16'hd53b;
        src25 <= 16'hebd3;
        src26 <= 16'hfed2;
        src27 <= 16'heacc;
        src28 <= 16'hd6b6;
        src29 <= 16'hdf72;
        src30 <= 16'h5e8e;
        src31 <= 16'h6649;
        src32 <= 16'hb28f;
        src33 <= 16'h364f;
        src34 <= 16'hea53;
        src35 <= 16'ha11e;
        src36 <= 16'hd3a8;
        src37 <= 16'he84f;
        src38 <= 16'h1752;
        src39 <= 16'h81e;
        src40 <= 16'hd479;
        src41 <= 16'hc074;
        src42 <= 16'h302c;
        src43 <= 16'hb7f5;
        src44 <= 16'h8bc8;
        src45 <= 16'h8d77;
        src46 <= 16'h196;
        src47 <= 16'h1595;
        src48 <= 16'ha067;
        src49 <= 16'hcf57;
        src50 <= 16'hd870;
        src51 <= 16'h50ed;
        src52 <= 16'h4a68;
        src53 <= 16'h4e5f;
        src54 <= 16'h4ae7;
        src55 <= 16'h3a29;
        src56 <= 16'hd2a3;
        src57 <= 16'h1e05;
        src58 <= 16'haa94;
        src59 <= 16'h8ed4;
        src60 <= 16'h4a50;
        src61 <= 16'h86c0;
        src62 <= 16'h1c68;
        src63 <= 16'h9784;
        src64 <= 16'h1e01;
        src65 <= 16'hdeac;
        src66 <= 16'hce7e;
        src67 <= 16'h8882;
        src68 <= 16'h6e82;
        src69 <= 16'h8ecf;
        src70 <= 16'h2f34;
        src71 <= 16'h8c3;
        src72 <= 16'h4da9;
        src73 <= 16'h8c7f;
        src74 <= 16'h91c1;
        src75 <= 16'hadaa;
        src76 <= 16'hce04;
        src77 <= 16'he6db;
        src78 <= 16'h2ec;
        src79 <= 16'h7edb;
        src80 <= 16'hdf56;
        src81 <= 16'h28cf;
        src82 <= 16'h9afd;
        src83 <= 16'hda0c;
        src84 <= 16'h177d;
        src85 <= 16'hbe67;
        src86 <= 16'hb6bc;
        src87 <= 16'h8f52;
        src88 <= 16'ha7f5;
        src89 <= 16'h5e94;
        src90 <= 16'h22eb;
        src91 <= 16'hbe99;
        src92 <= 16'hb205;
        src93 <= 16'h35e1;
        src94 <= 16'hc102;
        src95 <= 16'h729a;
        src96 <= 16'h15a8;
        src97 <= 16'h3918;
        src98 <= 16'hcdb4;
        src99 <= 16'ha01b;
        src100 <= 16'hb5af;
        src101 <= 16'h1e9e;
        src102 <= 16'h8088;
        src103 <= 16'h544a;
        src104 <= 16'h9f88;
        src105 <= 16'h6c95;
        src106 <= 16'hf7c9;
        src107 <= 16'ha3cd;
        src108 <= 16'ha2a0;
        src109 <= 16'h8d72;
        src110 <= 16'hd053;
        src111 <= 16'h8619;
        src112 <= 16'h72f5;
        src113 <= 16'hd5ab;
        src114 <= 16'h5f9b;
        src115 <= 16'h3bdc;
        src116 <= 16'h7aa;
        src117 <= 16'h2835;
        src118 <= 16'hc635;
        src119 <= 16'hb448;
        src120 <= 16'hfa97;
        src121 <= 16'h1651;
        src122 <= 16'haa39;
        src123 <= 16'hdd84;
        src124 <= 16'h909f;
        src125 <= 16'h8335;
        src126 <= 16'hb710;
        src127 <= 16'h2e65;
        src128 <= 16'hefe;
        src129 <= 16'h3294;
        src130 <= 16'h4fb0;
        src131 <= 16'h16ac;
        src132 <= 16'hfb0f;
        src133 <= 16'h26c7;
        src134 <= 16'h744f;
        src135 <= 16'h6eff;
        src136 <= 16'hadfa;
        src137 <= 16'h714c;
        src138 <= 16'hb771;
        src139 <= 16'h469a;
        src140 <= 16'hff33;
        src141 <= 16'h2c4e;
        src142 <= 16'h8748;
        src143 <= 16'h561e;
        src144 <= 16'h6947;
        src145 <= 16'h69e0;
        src146 <= 16'h226e;
        src147 <= 16'h4a7d;
        src148 <= 16'he356;
        src149 <= 16'h99ef;
        src150 <= 16'h7ec0;
        src151 <= 16'h88ba;
        src152 <= 16'h3ff3;
        src153 <= 16'hd5b;
        src154 <= 16'h3c6e;
        src155 <= 16'hc1c2;
        src156 <= 16'h1fb5;
        src157 <= 16'h78a5;
        src158 <= 16'h96f4;
        src159 <= 16'hb5c6;
        src160 <= 16'h1a96;
        src161 <= 16'h7d5b;
        exp <= 24'h5068ec;
        #1
        src0 <= 16'h2935;
        src1 <= 16'ha3c2;
        src2 <= 16'hd30e;
        src3 <= 16'h394c;
        src4 <= 16'he386;
        src5 <= 16'h786c;
        src6 <= 16'h5e5c;
        src7 <= 16'h3855;
        src8 <= 16'h4483;
        src9 <= 16'h817c;
        src10 <= 16'hbea2;
        src11 <= 16'h7527;
        src12 <= 16'h348f;
        src13 <= 16'hb862;
        src14 <= 16'h28a7;
        src15 <= 16'h9c45;
        src16 <= 16'he53b;
        src17 <= 16'ha89c;
        src18 <= 16'hd974;
        src19 <= 16'h965f;
        src20 <= 16'hfaaf;
        src21 <= 16'h6eed;
        src22 <= 16'hf140;
        src23 <= 16'hdf6e;
        src24 <= 16'hed91;
        src25 <= 16'h73;
        src26 <= 16'h5e94;
        src27 <= 16'hca6b;
        src28 <= 16'h348;
        src29 <= 16'h6977;
        src30 <= 16'h498e;
        src31 <= 16'h6b70;
        src32 <= 16'h7726;
        src33 <= 16'he84f;
        src34 <= 16'hb001;
        src35 <= 16'h4c01;
        src36 <= 16'h6122;
        src37 <= 16'h5e9a;
        src38 <= 16'h43a1;
        src39 <= 16'h1815;
        src40 <= 16'hb26a;
        src41 <= 16'h2ca6;
        src42 <= 16'h6e6;
        src43 <= 16'h4f71;
        src44 <= 16'h6b7c;
        src45 <= 16'h1795;
        src46 <= 16'he125;
        src47 <= 16'h37af;
        src48 <= 16'h773f;
        src49 <= 16'h3c04;
        src50 <= 16'hc118;
        src51 <= 16'h63c8;
        src52 <= 16'h757;
        src53 <= 16'h9a0e;
        src54 <= 16'h16bb;
        src55 <= 16'ha71c;
        src56 <= 16'he40d;
        src57 <= 16'h7adb;
        src58 <= 16'h28f8;
        src59 <= 16'h1f50;
        src60 <= 16'h28b5;
        src61 <= 16'hcf84;
        src62 <= 16'h29a1;
        src63 <= 16'ha015;
        src64 <= 16'hea8;
        src65 <= 16'hdff0;
        src66 <= 16'h7aa2;
        src67 <= 16'hbef;
        src68 <= 16'hcd60;
        src69 <= 16'h97e9;
        src70 <= 16'h9efa;
        src71 <= 16'hdf92;
        src72 <= 16'h25cb;
        src73 <= 16'haaa1;
        src74 <= 16'hd0c8;
        src75 <= 16'ha04;
        src76 <= 16'h1b3a;
        src77 <= 16'h6ce5;
        src78 <= 16'h61bb;
        src79 <= 16'h704d;
        src80 <= 16'hdf28;
        src81 <= 16'haf5a;
        src82 <= 16'h2e2a;
        src83 <= 16'h9dbf;
        src84 <= 16'h8396;
        src85 <= 16'hec57;
        src86 <= 16'hdaae;
        src87 <= 16'h4c88;
        src88 <= 16'h2177;
        src89 <= 16'hd6fa;
        src90 <= 16'haabe;
        src91 <= 16'h36d7;
        src92 <= 16'h3227;
        src93 <= 16'h4a0b;
        src94 <= 16'hc611;
        src95 <= 16'h9049;
        src96 <= 16'h96e5;
        src97 <= 16'hf14;
        src98 <= 16'hd888;
        src99 <= 16'hf967;
        src100 <= 16'hb42f;
        src101 <= 16'hbdca;
        src102 <= 16'hcdbf;
        src103 <= 16'h802c;
        src104 <= 16'h93a8;
        src105 <= 16'hbd7e;
        src106 <= 16'hecfa;
        src107 <= 16'h2032;
        src108 <= 16'hf927;
        src109 <= 16'h57ca;
        src110 <= 16'h4b0f;
        src111 <= 16'h7a33;
        src112 <= 16'hf2c4;
        src113 <= 16'h8394;
        src114 <= 16'h303c;
        src115 <= 16'h8867;
        src116 <= 16'hddcd;
        src117 <= 16'h8767;
        src118 <= 16'h77e9;
        src119 <= 16'hdbee;
        src120 <= 16'h89e5;
        src121 <= 16'h478a;
        src122 <= 16'h1ec7;
        src123 <= 16'h701;
        src124 <= 16'h2a32;
        src125 <= 16'h9908;
        src126 <= 16'hb786;
        src127 <= 16'h297c;
        src128 <= 16'hd5dc;
        src129 <= 16'h6f11;
        src130 <= 16'h1db1;
        src131 <= 16'hd203;
        src132 <= 16'hdcf2;
        src133 <= 16'h12a0;
        src134 <= 16'hae3b;
        src135 <= 16'h1388;
        src136 <= 16'h32c5;
        src137 <= 16'h4ba2;
        src138 <= 16'h44b0;
        src139 <= 16'h4761;
        src140 <= 16'h34e0;
        src141 <= 16'hc126;
        src142 <= 16'h8be2;
        src143 <= 16'h8e7e;
        src144 <= 16'hbc85;
        src145 <= 16'h9193;
        src146 <= 16'ha6d5;
        src147 <= 16'hca98;
        src148 <= 16'h908f;
        src149 <= 16'hde6b;
        src150 <= 16'h6475;
        src151 <= 16'h4bee;
        src152 <= 16'hdda;
        src153 <= 16'h68e0;
        src154 <= 16'h4693;
        src155 <= 16'h817c;
        src156 <= 16'h7304;
        src157 <= 16'he11f;
        src158 <= 16'h811;
        src159 <= 16'h61c1;
        src160 <= 16'h1fa0;
        src161 <= 16'h8142;
        exp <= 24'h4e7a9d;
        #1
        src0 <= 16'h719e;
        src1 <= 16'h93bb;
        src2 <= 16'h93cd;
        src3 <= 16'h13ad;
        src4 <= 16'h17c;
        src5 <= 16'h4569;
        src6 <= 16'hb463;
        src7 <= 16'he473;
        src8 <= 16'h30fb;
        src9 <= 16'hffa3;
        src10 <= 16'hc48f;
        src11 <= 16'h1388;
        src12 <= 16'h8b30;
        src13 <= 16'h738d;
        src14 <= 16'he602;
        src15 <= 16'he464;
        src16 <= 16'h526;
        src17 <= 16'h7eae;
        src18 <= 16'hfaeb;
        src19 <= 16'h28ea;
        src20 <= 16'h6cad;
        src21 <= 16'h7890;
        src22 <= 16'h59bd;
        src23 <= 16'h71d8;
        src24 <= 16'h2734;
        src25 <= 16'hdb91;
        src26 <= 16'hb1ad;
        src27 <= 16'h402;
        src28 <= 16'h1836;
        src29 <= 16'hdd98;
        src30 <= 16'h72e8;
        src31 <= 16'hc55b;
        src32 <= 16'hb4db;
        src33 <= 16'h46b5;
        src34 <= 16'ha5b5;
        src35 <= 16'h4911;
        src36 <= 16'h8c98;
        src37 <= 16'ha6d6;
        src38 <= 16'hd01d;
        src39 <= 16'h7821;
        src40 <= 16'h5513;
        src41 <= 16'hc849;
        src42 <= 16'h532a;
        src43 <= 16'h2022;
        src44 <= 16'h5659;
        src45 <= 16'h8df;
        src46 <= 16'h9b40;
        src47 <= 16'hb7d8;
        src48 <= 16'h33b8;
        src49 <= 16'h36ed;
        src50 <= 16'hce2;
        src51 <= 16'h2306;
        src52 <= 16'h33f9;
        src53 <= 16'h6c4e;
        src54 <= 16'he7b1;
        src55 <= 16'hfa2d;
        src56 <= 16'h289d;
        src57 <= 16'h5403;
        src58 <= 16'h5e14;
        src59 <= 16'h182b;
        src60 <= 16'h5860;
        src61 <= 16'he425;
        src62 <= 16'h5395;
        src63 <= 16'hfe73;
        src64 <= 16'h8af9;
        src65 <= 16'h477d;
        src66 <= 16'h9043;
        src67 <= 16'h467b;
        src68 <= 16'hc1b0;
        src69 <= 16'hf716;
        src70 <= 16'h8cc8;
        src71 <= 16'h88a3;
        src72 <= 16'h1353;
        src73 <= 16'hd1a2;
        src74 <= 16'h2d1a;
        src75 <= 16'hc740;
        src76 <= 16'h1fff;
        src77 <= 16'h25c6;
        src78 <= 16'hc1da;
        src79 <= 16'h92e6;
        src80 <= 16'he9a5;
        src81 <= 16'he8c;
        src82 <= 16'h4527;
        src83 <= 16'hcb8;
        src84 <= 16'h483f;
        src85 <= 16'hbdd;
        src86 <= 16'hdaf0;
        src87 <= 16'h4875;
        src88 <= 16'h7773;
        src89 <= 16'h7ced;
        src90 <= 16'h6508;
        src91 <= 16'h8c28;
        src92 <= 16'h177b;
        src93 <= 16'hbfb0;
        src94 <= 16'hd00a;
        src95 <= 16'h4442;
        src96 <= 16'h6db8;
        src97 <= 16'ha668;
        src98 <= 16'heea1;
        src99 <= 16'hc386;
        src100 <= 16'h9f5;
        src101 <= 16'h3a49;
        src102 <= 16'h3137;
        src103 <= 16'hec1a;
        src104 <= 16'h1570;
        src105 <= 16'h519e;
        src106 <= 16'hbc3f;
        src107 <= 16'hc093;
        src108 <= 16'hf926;
        src109 <= 16'hcbb0;
        src110 <= 16'h7dea;
        src111 <= 16'h45dc;
        src112 <= 16'hb9d;
        src113 <= 16'h851;
        src114 <= 16'h884;
        src115 <= 16'h677c;
        src116 <= 16'hf7a3;
        src117 <= 16'h9b1a;
        src118 <= 16'hc470;
        src119 <= 16'hab8;
        src120 <= 16'h9cb2;
        src121 <= 16'h43d8;
        src122 <= 16'h6103;
        src123 <= 16'h87a2;
        src124 <= 16'hc240;
        src125 <= 16'h7a3e;
        src126 <= 16'h349c;
        src127 <= 16'ha160;
        src128 <= 16'h814c;
        src129 <= 16'h2bd2;
        src130 <= 16'h9829;
        src131 <= 16'h9cc0;
        src132 <= 16'hed13;
        src133 <= 16'haa3b;
        src134 <= 16'hb795;
        src135 <= 16'h88d7;
        src136 <= 16'h323c;
        src137 <= 16'ha354;
        src138 <= 16'h7008;
        src139 <= 16'h8fdf;
        src140 <= 16'he23;
        src141 <= 16'h7416;
        src142 <= 16'h1db7;
        src143 <= 16'h9548;
        src144 <= 16'h4e7a;
        src145 <= 16'h23e;
        src146 <= 16'h2994;
        src147 <= 16'hc92e;
        src148 <= 16'h496b;
        src149 <= 16'hbb8b;
        src150 <= 16'hafcd;
        src151 <= 16'h6f5;
        src152 <= 16'h42c1;
        src153 <= 16'h95c5;
        src154 <= 16'h8c7d;
        src155 <= 16'h809f;
        src156 <= 16'he8f4;
        src157 <= 16'h8ff0;
        src158 <= 16'hb5de;
        src159 <= 16'h8cc6;
        src160 <= 16'h6ec4;
        src161 <= 16'h286;
        exp <= 24'h4b8e33;
        #1
        src0 <= 16'h1e35;
        src1 <= 16'h568e;
        src2 <= 16'hd207;
        src3 <= 16'h1d17;
        src4 <= 16'h5741;
        src5 <= 16'hb1cc;
        src6 <= 16'h897d;
        src7 <= 16'hcf0f;
        src8 <= 16'h4e99;
        src9 <= 16'h55d;
        src10 <= 16'h9cc4;
        src11 <= 16'h8041;
        src12 <= 16'ha02c;
        src13 <= 16'h37a0;
        src14 <= 16'hb5eb;
        src15 <= 16'hd3c8;
        src16 <= 16'h5d9f;
        src17 <= 16'hb558;
        src18 <= 16'h3f0a;
        src19 <= 16'h574;
        src20 <= 16'h5756;
        src21 <= 16'h6f24;
        src22 <= 16'h3ad7;
        src23 <= 16'hd8f;
        src24 <= 16'h92ae;
        src25 <= 16'h6717;
        src26 <= 16'h19f9;
        src27 <= 16'h8161;
        src28 <= 16'h5873;
        src29 <= 16'h63a0;
        src30 <= 16'h67e9;
        src31 <= 16'hbeb4;
        src32 <= 16'h81ed;
        src33 <= 16'h8a13;
        src34 <= 16'hd1f1;
        src35 <= 16'h65f0;
        src36 <= 16'hd7a0;
        src37 <= 16'h539c;
        src38 <= 16'h5723;
        src39 <= 16'h1150;
        src40 <= 16'h249;
        src41 <= 16'hc4ab;
        src42 <= 16'hcc38;
        src43 <= 16'h691a;
        src44 <= 16'h3821;
        src45 <= 16'h6200;
        src46 <= 16'haa16;
        src47 <= 16'h38;
        src48 <= 16'h89a9;
        src49 <= 16'h4bfe;
        src50 <= 16'hc944;
        src51 <= 16'h3aa7;
        src52 <= 16'h780c;
        src53 <= 16'h9f2e;
        src54 <= 16'h9e8d;
        src55 <= 16'hfa07;
        src56 <= 16'hd2c0;
        src57 <= 16'he153;
        src58 <= 16'h90a7;
        src59 <= 16'h677a;
        src60 <= 16'hb987;
        src61 <= 16'hca7f;
        src62 <= 16'ha937;
        src63 <= 16'hd443;
        src64 <= 16'hca92;
        src65 <= 16'h4be;
        src66 <= 16'hc07b;
        src67 <= 16'h2fed;
        src68 <= 16'h4846;
        src69 <= 16'h3eab;
        src70 <= 16'h741e;
        src71 <= 16'h2298;
        src72 <= 16'h40e0;
        src73 <= 16'h3375;
        src74 <= 16'h61f0;
        src75 <= 16'h7a2a;
        src76 <= 16'hbb97;
        src77 <= 16'hfc74;
        src78 <= 16'h2d1a;
        src79 <= 16'h8843;
        src80 <= 16'h4f55;
        src81 <= 16'h2448;
        src82 <= 16'h57c3;
        src83 <= 16'h4a09;
        src84 <= 16'h3428;
        src85 <= 16'h2971;
        src86 <= 16'h84d9;
        src87 <= 16'he86;
        src88 <= 16'hadf9;
        src89 <= 16'h2c9e;
        src90 <= 16'h3e0d;
        src91 <= 16'had56;
        src92 <= 16'h3afe;
        src93 <= 16'h2a40;
        src94 <= 16'haac7;
        src95 <= 16'hf4b4;
        src96 <= 16'h9fce;
        src97 <= 16'h371d;
        src98 <= 16'h191;
        src99 <= 16'h2f8a;
        src100 <= 16'h31d2;
        src101 <= 16'hc559;
        src102 <= 16'h405c;
        src103 <= 16'h3073;
        src104 <= 16'h26c7;
        src105 <= 16'hb920;
        src106 <= 16'hf9a1;
        src107 <= 16'heaa2;
        src108 <= 16'h188e;
        src109 <= 16'hbb9a;
        src110 <= 16'h5ece;
        src111 <= 16'h4b93;
        src112 <= 16'h95ba;
        src113 <= 16'h5232;
        src114 <= 16'hc30a;
        src115 <= 16'h81f4;
        src116 <= 16'h30fb;
        src117 <= 16'heb2c;
        src118 <= 16'hcc66;
        src119 <= 16'h7077;
        src120 <= 16'h73c1;
        src121 <= 16'ha7de;
        src122 <= 16'h886b;
        src123 <= 16'h2c4c;
        src124 <= 16'h3cb9;
        src125 <= 16'h46d9;
        src126 <= 16'h3c2a;
        src127 <= 16'hefc9;
        src128 <= 16'h6c3c;
        src129 <= 16'h4d14;
        src130 <= 16'h7d58;
        src131 <= 16'he690;
        src132 <= 16'he572;
        src133 <= 16'hdc51;
        src134 <= 16'ha477;
        src135 <= 16'h8eb1;
        src136 <= 16'h8e9f;
        src137 <= 16'hbd9f;
        src138 <= 16'h6e1b;
        src139 <= 16'h9146;
        src140 <= 16'h81da;
        src141 <= 16'hb781;
        src142 <= 16'h8c3;
        src143 <= 16'h9979;
        src144 <= 16'hb536;
        src145 <= 16'h4a04;
        src146 <= 16'h2a34;
        src147 <= 16'h3c77;
        src148 <= 16'h5471;
        src149 <= 16'h5617;
        src150 <= 16'h454f;
        src151 <= 16'h6a9c;
        src152 <= 16'h5e3f;
        src153 <= 16'h5558;
        src154 <= 16'hd479;
        src155 <= 16'h1608;
        src156 <= 16'h256;
        src157 <= 16'h95aa;
        src158 <= 16'h6c17;
        src159 <= 16'h4dcc;
        src160 <= 16'hd3e0;
        src161 <= 16'hc7bc;
        exp <= 24'h4a6f7f;
        #1
        src0 <= 16'he480;
        src1 <= 16'h4a03;
        src2 <= 16'ha123;
        src3 <= 16'ha0c4;
        src4 <= 16'he129;
        src5 <= 16'h7f14;
        src6 <= 16'ha684;
        src7 <= 16'h1eda;
        src8 <= 16'h3f4a;
        src9 <= 16'h9f4d;
        src10 <= 16'ha365;
        src11 <= 16'h33c5;
        src12 <= 16'h50ea;
        src13 <= 16'h3ab4;
        src14 <= 16'h4dfa;
        src15 <= 16'heb22;
        src16 <= 16'h8b6;
        src17 <= 16'h6772;
        src18 <= 16'h7e60;
        src19 <= 16'h6669;
        src20 <= 16'h2385;
        src21 <= 16'h8ee6;
        src22 <= 16'h7020;
        src23 <= 16'ha916;
        src24 <= 16'h5c31;
        src25 <= 16'he79b;
        src26 <= 16'h4ba8;
        src27 <= 16'h3bc;
        src28 <= 16'h23eb;
        src29 <= 16'h28b2;
        src30 <= 16'h62f5;
        src31 <= 16'hcd90;
        src32 <= 16'h2d52;
        src33 <= 16'h7a89;
        src34 <= 16'hcee9;
        src35 <= 16'h2bd2;
        src36 <= 16'hefe9;
        src37 <= 16'h75da;
        src38 <= 16'hba27;
        src39 <= 16'he5e9;
        src40 <= 16'hea60;
        src41 <= 16'hceb;
        src42 <= 16'h4982;
        src43 <= 16'h57ef;
        src44 <= 16'h28dc;
        src45 <= 16'h5218;
        src46 <= 16'h41d;
        src47 <= 16'hd7a1;
        src48 <= 16'hf163;
        src49 <= 16'ha791;
        src50 <= 16'h5e64;
        src51 <= 16'hc4e1;
        src52 <= 16'h7f25;
        src53 <= 16'h6925;
        src54 <= 16'ha578;
        src55 <= 16'he6c8;
        src56 <= 16'hd9ca;
        src57 <= 16'h13f7;
        src58 <= 16'h1c7b;
        src59 <= 16'he0ca;
        src60 <= 16'heac7;
        src61 <= 16'hab91;
        src62 <= 16'ha316;
        src63 <= 16'h3e12;
        src64 <= 16'h8772;
        src65 <= 16'he6ee;
        src66 <= 16'h4e4a;
        src67 <= 16'h7083;
        src68 <= 16'h6987;
        src69 <= 16'h7b1b;
        src70 <= 16'h20c5;
        src71 <= 16'ha3bd;
        src72 <= 16'he862;
        src73 <= 16'h788a;
        src74 <= 16'hb872;
        src75 <= 16'h6679;
        src76 <= 16'hd004;
        src77 <= 16'h5e2f;
        src78 <= 16'hdfe;
        src79 <= 16'h3998;
        src80 <= 16'h2f56;
        src81 <= 16'h20b2;
        src82 <= 16'h2a5e;
        src83 <= 16'h59d8;
        src84 <= 16'h8c5d;
        src85 <= 16'h25d4;
        src86 <= 16'hf817;
        src87 <= 16'h7b9f;
        src88 <= 16'h2431;
        src89 <= 16'hc051;
        src90 <= 16'he965;
        src91 <= 16'hb2a2;
        src92 <= 16'h973;
        src93 <= 16'h1d58;
        src94 <= 16'h2c2;
        src95 <= 16'hc418;
        src96 <= 16'hdc0d;
        src97 <= 16'hecb0;
        src98 <= 16'h8aa5;
        src99 <= 16'h83f9;
        src100 <= 16'h82d2;
        src101 <= 16'h6226;
        src102 <= 16'h9b23;
        src103 <= 16'heb74;
        src104 <= 16'h158e;
        src105 <= 16'h21a;
        src106 <= 16'hf014;
        src107 <= 16'h5446;
        src108 <= 16'hd81b;
        src109 <= 16'h6904;
        src110 <= 16'hda7c;
        src111 <= 16'hefe0;
        src112 <= 16'h66ec;
        src113 <= 16'he64;
        src114 <= 16'h5e95;
        src115 <= 16'h4d50;
        src116 <= 16'hb6ec;
        src117 <= 16'hecae;
        src118 <= 16'h5f57;
        src119 <= 16'h6c5c;
        src120 <= 16'h8eca;
        src121 <= 16'h785a;
        src122 <= 16'h89b4;
        src123 <= 16'h8fed;
        src124 <= 16'h9432;
        src125 <= 16'h24b4;
        src126 <= 16'he51e;
        src127 <= 16'h8e9b;
        src128 <= 16'h879b;
        src129 <= 16'hf750;
        src130 <= 16'h3d7b;
        src131 <= 16'hae26;
        src132 <= 16'h3008;
        src133 <= 16'h9da8;
        src134 <= 16'he86e;
        src135 <= 16'h15a8;
        src136 <= 16'h8898;
        src137 <= 16'hd8c;
        src138 <= 16'hf8ad;
        src139 <= 16'h1bae;
        src140 <= 16'h42c0;
        src141 <= 16'h6ae0;
        src142 <= 16'h2693;
        src143 <= 16'h6da3;
        src144 <= 16'ha70e;
        src145 <= 16'hdb77;
        src146 <= 16'h150e;
        src147 <= 16'hff19;
        src148 <= 16'hdc71;
        src149 <= 16'h635a;
        src150 <= 16'he382;
        src151 <= 16'hd576;
        src152 <= 16'hfdc6;
        src153 <= 16'h2263;
        src154 <= 16'h3a83;
        src155 <= 16'h5867;
        src156 <= 16'hf9b9;
        src157 <= 16'hbdb7;
        src158 <= 16'h6bc7;
        src159 <= 16'hf6e5;
        src160 <= 16'h7199;
        src161 <= 16'h85f5;
        exp <= 24'h519fe8;
        #1
        src0 <= 16'heed7;
        src1 <= 16'h5d93;
        src2 <= 16'hed72;
        src3 <= 16'h6400;
        src4 <= 16'h8121;
        src5 <= 16'h8fbb;
        src6 <= 16'hdd9c;
        src7 <= 16'h6c3;
        src8 <= 16'h63f6;
        src9 <= 16'h4536;
        src10 <= 16'hc83c;
        src11 <= 16'h2ecc;
        src12 <= 16'hd6c8;
        src13 <= 16'h2a81;
        src14 <= 16'hec0d;
        src15 <= 16'hff90;
        src16 <= 16'h7721;
        src17 <= 16'h11b2;
        src18 <= 16'h84f2;
        src19 <= 16'hba41;
        src20 <= 16'hc874;
        src21 <= 16'hbd16;
        src22 <= 16'hca67;
        src23 <= 16'h3c9f;
        src24 <= 16'h86a8;
        src25 <= 16'h20d8;
        src26 <= 16'h331;
        src27 <= 16'h84b2;
        src28 <= 16'h3be3;
        src29 <= 16'h6fed;
        src30 <= 16'hf576;
        src31 <= 16'h1510;
        src32 <= 16'h45dc;
        src33 <= 16'hbd60;
        src34 <= 16'h2c9a;
        src35 <= 16'h1996;
        src36 <= 16'hd73c;
        src37 <= 16'hb843;
        src38 <= 16'he0e3;
        src39 <= 16'hda88;
        src40 <= 16'h3964;
        src41 <= 16'ha702;
        src42 <= 16'h5b86;
        src43 <= 16'h56b;
        src44 <= 16'hf539;
        src45 <= 16'hcbd5;
        src46 <= 16'h5005;
        src47 <= 16'hce0a;
        src48 <= 16'hdb3f;
        src49 <= 16'h8a77;
        src50 <= 16'h9ff1;
        src51 <= 16'h76a8;
        src52 <= 16'h2e1b;
        src53 <= 16'hd7ce;
        src54 <= 16'h2fc0;
        src55 <= 16'h9368;
        src56 <= 16'h9f27;
        src57 <= 16'h4689;
        src58 <= 16'h29fd;
        src59 <= 16'h9cce;
        src60 <= 16'ha2ce;
        src61 <= 16'hb6ae;
        src62 <= 16'heda0;
        src63 <= 16'h80c9;
        src64 <= 16'h6975;
        src65 <= 16'ha240;
        src66 <= 16'h44de;
        src67 <= 16'hda8b;
        src68 <= 16'hc5ee;
        src69 <= 16'h6805;
        src70 <= 16'ha992;
        src71 <= 16'hd40a;
        src72 <= 16'hedc0;
        src73 <= 16'h7e1;
        src74 <= 16'h5beb;
        src75 <= 16'he699;
        src76 <= 16'hba2a;
        src77 <= 16'h3a5d;
        src78 <= 16'h22e1;
        src79 <= 16'hf031;
        src80 <= 16'h1b18;
        src81 <= 16'hffe1;
        src82 <= 16'hbb51;
        src83 <= 16'hfb42;
        src84 <= 16'h80f5;
        src85 <= 16'he374;
        src86 <= 16'hff72;
        src87 <= 16'hc8a1;
        src88 <= 16'hb32e;
        src89 <= 16'h1cc8;
        src90 <= 16'hab35;
        src91 <= 16'he0e6;
        src92 <= 16'h12ac;
        src93 <= 16'h7ca1;
        src94 <= 16'hbd1c;
        src95 <= 16'hd9da;
        src96 <= 16'h8a4a;
        src97 <= 16'h13b5;
        src98 <= 16'h6dc5;
        src99 <= 16'h9109;
        src100 <= 16'hd5c2;
        src101 <= 16'hbf42;
        src102 <= 16'h16a8;
        src103 <= 16'hf9ad;
        src104 <= 16'hb285;
        src105 <= 16'h79c0;
        src106 <= 16'h6cd6;
        src107 <= 16'hfe32;
        src108 <= 16'h1316;
        src109 <= 16'h29eb;
        src110 <= 16'h1f2;
        src111 <= 16'h8d2c;
        src112 <= 16'he7b9;
        src113 <= 16'h698e;
        src114 <= 16'h31f6;
        src115 <= 16'hbc30;
        src116 <= 16'hc73e;
        src117 <= 16'h5784;
        src118 <= 16'hc2df;
        src119 <= 16'hfccd;
        src120 <= 16'hc81d;
        src121 <= 16'h26f9;
        src122 <= 16'ha90f;
        src123 <= 16'h668;
        src124 <= 16'h1223;
        src125 <= 16'h5e4e;
        src126 <= 16'h3743;
        src127 <= 16'hbe3;
        src128 <= 16'h28;
        src129 <= 16'h6e8c;
        src130 <= 16'hf3b1;
        src131 <= 16'h38f6;
        src132 <= 16'hd773;
        src133 <= 16'hdaf0;
        src134 <= 16'hb21b;
        src135 <= 16'h390a;
        src136 <= 16'hedc;
        src137 <= 16'hd60;
        src138 <= 16'h5a69;
        src139 <= 16'h9fd2;
        src140 <= 16'h2507;
        src141 <= 16'h2acd;
        src142 <= 16'h16c7;
        src143 <= 16'h6708;
        src144 <= 16'hfb96;
        src145 <= 16'ha6e4;
        src146 <= 16'h6666;
        src147 <= 16'hab9d;
        src148 <= 16'h8baa;
        src149 <= 16'hd072;
        src150 <= 16'h4007;
        src151 <= 16'hec8d;
        src152 <= 16'hbae8;
        src153 <= 16'ha07;
        src154 <= 16'h67ba;
        src155 <= 16'h8f2a;
        src156 <= 16'h77e2;
        src157 <= 16'h6dd7;
        src158 <= 16'h7d56;
        src159 <= 16'h2b10;
        src160 <= 16'hb6e9;
        src161 <= 16'haca;
        exp <= 24'h53db31;
        #1
        src0 <= 16'h2123;
        src1 <= 16'h953c;
        src2 <= 16'h5147;
        src3 <= 16'h6802;
        src4 <= 16'had71;
        src5 <= 16'h6025;
        src6 <= 16'hb608;
        src7 <= 16'he590;
        src8 <= 16'hb386;
        src9 <= 16'h64cf;
        src10 <= 16'hbcb8;
        src11 <= 16'h42ff;
        src12 <= 16'h2c3d;
        src13 <= 16'he2ed;
        src14 <= 16'h7a68;
        src15 <= 16'h4f65;
        src16 <= 16'hc1b7;
        src17 <= 16'h10fb;
        src18 <= 16'hed4e;
        src19 <= 16'h784e;
        src20 <= 16'hefa;
        src21 <= 16'hd77b;
        src22 <= 16'h6294;
        src23 <= 16'h43d7;
        src24 <= 16'h402f;
        src25 <= 16'hddd7;
        src26 <= 16'hda0c;
        src27 <= 16'h7690;
        src28 <= 16'h1d35;
        src29 <= 16'hf8fe;
        src30 <= 16'h7864;
        src31 <= 16'h925c;
        src32 <= 16'hc511;
        src33 <= 16'h120a;
        src34 <= 16'hdccc;
        src35 <= 16'hb7f7;
        src36 <= 16'h1947;
        src37 <= 16'h175e;
        src38 <= 16'h9f07;
        src39 <= 16'h2f45;
        src40 <= 16'h4b70;
        src41 <= 16'h1ccb;
        src42 <= 16'h3580;
        src43 <= 16'h47f7;
        src44 <= 16'h4ad5;
        src45 <= 16'hcc3d;
        src46 <= 16'he4b6;
        src47 <= 16'h784;
        src48 <= 16'h699;
        src49 <= 16'h1d3c;
        src50 <= 16'h6187;
        src51 <= 16'h793c;
        src52 <= 16'h5108;
        src53 <= 16'h2e95;
        src54 <= 16'h7607;
        src55 <= 16'h3c60;
        src56 <= 16'ha2ea;
        src57 <= 16'h9bff;
        src58 <= 16'h3e69;
        src59 <= 16'hbe8e;
        src60 <= 16'h187c;
        src61 <= 16'hcbfe;
        src62 <= 16'h1553;
        src63 <= 16'h33c1;
        src64 <= 16'h2d20;
        src65 <= 16'h80a4;
        src66 <= 16'h9b76;
        src67 <= 16'hc15;
        src68 <= 16'h6654;
        src69 <= 16'h5c8e;
        src70 <= 16'h547c;
        src71 <= 16'he5d7;
        src72 <= 16'h355;
        src73 <= 16'h25e2;
        src74 <= 16'hd357;
        src75 <= 16'h85e1;
        src76 <= 16'h2c1;
        src77 <= 16'h495a;
        src78 <= 16'h7ed2;
        src79 <= 16'h14a7;
        src80 <= 16'h987;
        src81 <= 16'hfbeb;
        src82 <= 16'h8a45;
        src83 <= 16'h8492;
        src84 <= 16'h21c5;
        src85 <= 16'hd698;
        src86 <= 16'h7e16;
        src87 <= 16'hed7d;
        src88 <= 16'hf0b8;
        src89 <= 16'h9b08;
        src90 <= 16'he638;
        src91 <= 16'h68e5;
        src92 <= 16'ha69c;
        src93 <= 16'h9e1f;
        src94 <= 16'h87a1;
        src95 <= 16'h69ef;
        src96 <= 16'hc2d1;
        src97 <= 16'hf349;
        src98 <= 16'ha64a;
        src99 <= 16'hcea5;
        src100 <= 16'h78b3;
        src101 <= 16'h5474;
        src102 <= 16'h6c79;
        src103 <= 16'h5d75;
        src104 <= 16'hb6e7;
        src105 <= 16'hdff9;
        src106 <= 16'h3408;
        src107 <= 16'ha841;
        src108 <= 16'hab3b;
        src109 <= 16'h5f93;
        src110 <= 16'h25d6;
        src111 <= 16'h14ec;
        src112 <= 16'h2974;
        src113 <= 16'h29a2;
        src114 <= 16'hda96;
        src115 <= 16'hd9ae;
        src116 <= 16'hd190;
        src117 <= 16'h5a83;
        src118 <= 16'hcaf8;
        src119 <= 16'h1427;
        src120 <= 16'h8ea6;
        src121 <= 16'h1298;
        src122 <= 16'h5b8e;
        src123 <= 16'hd7ee;
        src124 <= 16'hd4b8;
        src125 <= 16'hc5ba;
        src126 <= 16'h70aa;
        src127 <= 16'h1d34;
        src128 <= 16'h16df;
        src129 <= 16'h7bc6;
        src130 <= 16'h7bab;
        src131 <= 16'h47d;
        src132 <= 16'hac2;
        src133 <= 16'h4b4c;
        src134 <= 16'he143;
        src135 <= 16'h87b9;
        src136 <= 16'h1db3;
        src137 <= 16'h1f3a;
        src138 <= 16'h771c;
        src139 <= 16'h935b;
        src140 <= 16'h8ee4;
        src141 <= 16'hfcee;
        src142 <= 16'h7a;
        src143 <= 16'hbed2;
        src144 <= 16'hb617;
        src145 <= 16'h4657;
        src146 <= 16'h5c13;
        src147 <= 16'hbf5;
        src148 <= 16'h8a68;
        src149 <= 16'h3e9f;
        src150 <= 16'he2d0;
        src151 <= 16'hacd9;
        src152 <= 16'h55b0;
        src153 <= 16'hfc52;
        src154 <= 16'he95a;
        src155 <= 16'he4bf;
        src156 <= 16'ha97e;
        src157 <= 16'h29be;
        src158 <= 16'h31d8;
        src159 <= 16'h249b;
        src160 <= 16'hf492;
        src161 <= 16'h52e7;
        exp <= 24'h4bc78a;
        #1
        src0 <= 16'h38bf;
        src1 <= 16'h560c;
        src2 <= 16'he326;
        src3 <= 16'h1cc2;
        src4 <= 16'hb89d;
        src5 <= 16'h3629;
        src6 <= 16'hff9c;
        src7 <= 16'h79a1;
        src8 <= 16'ha5d;
        src9 <= 16'ha039;
        src10 <= 16'he7dd;
        src11 <= 16'h9ae5;
        src12 <= 16'h49b2;
        src13 <= 16'hd6ae;
        src14 <= 16'h6b47;
        src15 <= 16'h272d;
        src16 <= 16'h4369;
        src17 <= 16'h5a2a;
        src18 <= 16'hc0ff;
        src19 <= 16'h7017;
        src20 <= 16'h917c;
        src21 <= 16'h907d;
        src22 <= 16'h903d;
        src23 <= 16'h23cc;
        src24 <= 16'hb83f;
        src25 <= 16'hcc69;
        src26 <= 16'h1350;
        src27 <= 16'h792f;
        src28 <= 16'he2b4;
        src29 <= 16'hbf2e;
        src30 <= 16'h10e0;
        src31 <= 16'h8109;
        src32 <= 16'he640;
        src33 <= 16'h1b39;
        src34 <= 16'h4c43;
        src35 <= 16'h1fa8;
        src36 <= 16'h5a2c;
        src37 <= 16'h81d7;
        src38 <= 16'h16fa;
        src39 <= 16'h8873;
        src40 <= 16'h359c;
        src41 <= 16'h2514;
        src42 <= 16'h6ce7;
        src43 <= 16'h7b80;
        src44 <= 16'h89de;
        src45 <= 16'ha952;
        src46 <= 16'h1046;
        src47 <= 16'h1774;
        src48 <= 16'h5f84;
        src49 <= 16'h395b;
        src50 <= 16'hca34;
        src51 <= 16'h25f8;
        src52 <= 16'h52ab;
        src53 <= 16'h2372;
        src54 <= 16'had8f;
        src55 <= 16'h9ec6;
        src56 <= 16'h60bd;
        src57 <= 16'h92f4;
        src58 <= 16'h422e;
        src59 <= 16'hf368;
        src60 <= 16'h705f;
        src61 <= 16'h1e89;
        src62 <= 16'h168e;
        src63 <= 16'h4cd8;
        src64 <= 16'haa06;
        src65 <= 16'hd486;
        src66 <= 16'h6298;
        src67 <= 16'hcafd;
        src68 <= 16'h9a9c;
        src69 <= 16'h9142;
        src70 <= 16'hac41;
        src71 <= 16'ha8d5;
        src72 <= 16'h26c3;
        src73 <= 16'had79;
        src74 <= 16'h3d5c;
        src75 <= 16'hb11b;
        src76 <= 16'h9fb1;
        src77 <= 16'hb240;
        src78 <= 16'h95b1;
        src79 <= 16'h69f6;
        src80 <= 16'hb3a1;
        src81 <= 16'ha1af;
        src82 <= 16'hb4be;
        src83 <= 16'h8ed7;
        src84 <= 16'hc3f3;
        src85 <= 16'h7258;
        src86 <= 16'h6b28;
        src87 <= 16'hed79;
        src88 <= 16'hc2db;
        src89 <= 16'h6051;
        src90 <= 16'hd772;
        src91 <= 16'h9436;
        src92 <= 16'h5ffd;
        src93 <= 16'h4e88;
        src94 <= 16'hf786;
        src95 <= 16'h9dee;
        src96 <= 16'h84d2;
        src97 <= 16'h7813;
        src98 <= 16'h7d95;
        src99 <= 16'h62a2;
        src100 <= 16'hbe28;
        src101 <= 16'h9c32;
        src102 <= 16'hb970;
        src103 <= 16'h1fe8;
        src104 <= 16'h7720;
        src105 <= 16'h9b18;
        src106 <= 16'h53ad;
        src107 <= 16'hccf7;
        src108 <= 16'hec9d;
        src109 <= 16'h8700;
        src110 <= 16'h9ba2;
        src111 <= 16'h74e6;
        src112 <= 16'h4849;
        src113 <= 16'h86a4;
        src114 <= 16'h9700;
        src115 <= 16'h25f3;
        src116 <= 16'he878;
        src117 <= 16'haff9;
        src118 <= 16'hc566;
        src119 <= 16'hed0a;
        src120 <= 16'h664e;
        src121 <= 16'h9abd;
        src122 <= 16'he724;
        src123 <= 16'ha495;
        src124 <= 16'hca40;
        src125 <= 16'h4030;
        src126 <= 16'hbc9e;
        src127 <= 16'h76ae;
        src128 <= 16'h2936;
        src129 <= 16'h70af;
        src130 <= 16'hca18;
        src131 <= 16'hfd58;
        src132 <= 16'h2400;
        src133 <= 16'hf144;
        src134 <= 16'h404e;
        src135 <= 16'h2146;
        src136 <= 16'h2df0;
        src137 <= 16'h7260;
        src138 <= 16'h24ac;
        src139 <= 16'hd7f8;
        src140 <= 16'h1670;
        src141 <= 16'hb486;
        src142 <= 16'h6429;
        src143 <= 16'h6d92;
        src144 <= 16'h3bf1;
        src145 <= 16'h41e0;
        src146 <= 16'h3e3b;
        src147 <= 16'hecae;
        src148 <= 16'h45f3;
        src149 <= 16'hf02f;
        src150 <= 16'h9f0;
        src151 <= 16'h7607;
        src152 <= 16'hc895;
        src153 <= 16'h29f2;
        src154 <= 16'hbcde;
        src155 <= 16'h4d2a;
        src156 <= 16'hc19f;
        src157 <= 16'h3751;
        src158 <= 16'hef70;
        src159 <= 16'h17ce;
        src160 <= 16'h1d86;
        src161 <= 16'h88eb;
        exp <= 24'h506747;
        #1
        src0 <= 16'hfa39;
        src1 <= 16'h7f7c;
        src2 <= 16'h9e3c;
        src3 <= 16'h6098;
        src4 <= 16'hb6b1;
        src5 <= 16'hc964;
        src6 <= 16'h1534;
        src7 <= 16'hb7ee;
        src8 <= 16'hb6fe;
        src9 <= 16'h7586;
        src10 <= 16'h1f08;
        src11 <= 16'hffe9;
        src12 <= 16'h2c9c;
        src13 <= 16'h5d0a;
        src14 <= 16'he5f6;
        src15 <= 16'hce2a;
        src16 <= 16'h13bf;
        src17 <= 16'ha80d;
        src18 <= 16'h62c3;
        src19 <= 16'h4de9;
        src20 <= 16'hcc36;
        src21 <= 16'ha034;
        src22 <= 16'he682;
        src23 <= 16'hc5cc;
        src24 <= 16'hd8ad;
        src25 <= 16'ha01e;
        src26 <= 16'h67f5;
        src27 <= 16'h41c7;
        src28 <= 16'h5404;
        src29 <= 16'h5293;
        src30 <= 16'h9f2b;
        src31 <= 16'h4066;
        src32 <= 16'h9607;
        src33 <= 16'hd23e;
        src34 <= 16'hfd20;
        src35 <= 16'hb28e;
        src36 <= 16'hca21;
        src37 <= 16'had6e;
        src38 <= 16'h1c4d;
        src39 <= 16'hefee;
        src40 <= 16'h9277;
        src41 <= 16'hac2e;
        src42 <= 16'hbcd3;
        src43 <= 16'h878f;
        src44 <= 16'h1aa0;
        src45 <= 16'h5779;
        src46 <= 16'h7cec;
        src47 <= 16'hf142;
        src48 <= 16'h486e;
        src49 <= 16'h1b;
        src50 <= 16'h5715;
        src51 <= 16'h4a97;
        src52 <= 16'hc1ee;
        src53 <= 16'h31ed;
        src54 <= 16'hf377;
        src55 <= 16'hff63;
        src56 <= 16'hafe5;
        src57 <= 16'h1ebb;
        src58 <= 16'h4fc1;
        src59 <= 16'hf535;
        src60 <= 16'hb87e;
        src61 <= 16'hb084;
        src62 <= 16'h6409;
        src63 <= 16'h7a25;
        src64 <= 16'hf7f9;
        src65 <= 16'h7d91;
        src66 <= 16'he7;
        src67 <= 16'hd728;
        src68 <= 16'h1c21;
        src69 <= 16'hfd78;
        src70 <= 16'hfa6c;
        src71 <= 16'hadae;
        src72 <= 16'hb0ad;
        src73 <= 16'hda5b;
        src74 <= 16'h544;
        src75 <= 16'h6ea8;
        src76 <= 16'h44f6;
        src77 <= 16'h8cf6;
        src78 <= 16'h2fdd;
        src79 <= 16'h2c70;
        src80 <= 16'he82b;
        src81 <= 16'h25b;
        src82 <= 16'h7326;
        src83 <= 16'h9657;
        src84 <= 16'h16bc;
        src85 <= 16'h8277;
        src86 <= 16'hf26f;
        src87 <= 16'h6b8e;
        src88 <= 16'h2ea2;
        src89 <= 16'he6a2;
        src90 <= 16'h40ca;
        src91 <= 16'h7641;
        src92 <= 16'h6184;
        src93 <= 16'ha99c;
        src94 <= 16'h38;
        src95 <= 16'ha956;
        src96 <= 16'hcf;
        src97 <= 16'h9286;
        src98 <= 16'h7c68;
        src99 <= 16'h74b5;
        src100 <= 16'h48a8;
        src101 <= 16'h9147;
        src102 <= 16'h45eb;
        src103 <= 16'h91bc;
        src104 <= 16'hf020;
        src105 <= 16'he05d;
        src106 <= 16'h1686;
        src107 <= 16'h1020;
        src108 <= 16'h39d1;
        src109 <= 16'he8a9;
        src110 <= 16'h357b;
        src111 <= 16'h167e;
        src112 <= 16'h3b31;
        src113 <= 16'hb4c2;
        src114 <= 16'hcb0b;
        src115 <= 16'h362d;
        src116 <= 16'ha7e7;
        src117 <= 16'h6d89;
        src118 <= 16'h6b8d;
        src119 <= 16'h437f;
        src120 <= 16'h8140;
        src121 <= 16'hb606;
        src122 <= 16'h7851;
        src123 <= 16'h14d2;
        src124 <= 16'hba8d;
        src125 <= 16'hadef;
        src126 <= 16'h273a;
        src127 <= 16'h1e88;
        src128 <= 16'hf256;
        src129 <= 16'h49cc;
        src130 <= 16'h6d4c;
        src131 <= 16'h21b9;
        src132 <= 16'hc2a8;
        src133 <= 16'h702;
        src134 <= 16'h2d95;
        src135 <= 16'h58cc;
        src136 <= 16'hdf4a;
        src137 <= 16'h4f3b;
        src138 <= 16'h68e7;
        src139 <= 16'h5215;
        src140 <= 16'hb38c;
        src141 <= 16'hb8b2;
        src142 <= 16'hd6ee;
        src143 <= 16'hafcb;
        src144 <= 16'haa6c;
        src145 <= 16'hb605;
        src146 <= 16'h1971;
        src147 <= 16'h89d7;
        src148 <= 16'h820e;
        src149 <= 16'h192e;
        src150 <= 16'hd454;
        src151 <= 16'h75d7;
        src152 <= 16'h40dc;
        src153 <= 16'h7a7a;
        src154 <= 16'hc1ad;
        src155 <= 16'h6dd1;
        src156 <= 16'hf8c5;
        src157 <= 16'h5f7;
        src158 <= 16'h7eca;
        src159 <= 16'h10ae;
        src160 <= 16'h5bab;
        src161 <= 16'hc099;
        exp <= 24'h518a40;
        #1
        src0 <= 16'h7cb9;
        src1 <= 16'hc899;
        src2 <= 16'haadb;
        src3 <= 16'h2aba;
        src4 <= 16'hfbdf;
        src5 <= 16'hf586;
        src6 <= 16'h7450;
        src7 <= 16'h978b;
        src8 <= 16'ha1f;
        src9 <= 16'hf880;
        src10 <= 16'haefd;
        src11 <= 16'h94ff;
        src12 <= 16'h6af0;
        src13 <= 16'hcbdf;
        src14 <= 16'h6d5e;
        src15 <= 16'hdf67;
        src16 <= 16'h3462;
        src17 <= 16'h4601;
        src18 <= 16'h8355;
        src19 <= 16'h5295;
        src20 <= 16'hbff3;
        src21 <= 16'h9ade;
        src22 <= 16'hc3ae;
        src23 <= 16'h8635;
        src24 <= 16'h58a8;
        src25 <= 16'h40dc;
        src26 <= 16'h2334;
        src27 <= 16'h8126;
        src28 <= 16'hf4fc;
        src29 <= 16'h81f9;
        src30 <= 16'hefa7;
        src31 <= 16'hf59a;
        src32 <= 16'hafc;
        src33 <= 16'hbbc9;
        src34 <= 16'h73b9;
        src35 <= 16'h2005;
        src36 <= 16'h560e;
        src37 <= 16'h6528;
        src38 <= 16'hbbfc;
        src39 <= 16'h8b9b;
        src40 <= 16'h6af5;
        src41 <= 16'h6ed7;
        src42 <= 16'ha9a3;
        src43 <= 16'h85a0;
        src44 <= 16'h3e55;
        src45 <= 16'h8e10;
        src46 <= 16'ha5b1;
        src47 <= 16'ha329;
        src48 <= 16'h17ee;
        src49 <= 16'hb142;
        src50 <= 16'hab6b;
        src51 <= 16'h4779;
        src52 <= 16'h8f06;
        src53 <= 16'hd914;
        src54 <= 16'h3f1e;
        src55 <= 16'hb22b;
        src56 <= 16'h9ca;
        src57 <= 16'hc21b;
        src58 <= 16'h7065;
        src59 <= 16'hd13b;
        src60 <= 16'hd66b;
        src61 <= 16'hedeb;
        src62 <= 16'h3d91;
        src63 <= 16'hd8ea;
        src64 <= 16'ha040;
        src65 <= 16'h8421;
        src66 <= 16'h8087;
        src67 <= 16'h70c4;
        src68 <= 16'h6d4a;
        src69 <= 16'hf3bd;
        src70 <= 16'h561;
        src71 <= 16'h4361;
        src72 <= 16'h30ed;
        src73 <= 16'h5038;
        src74 <= 16'h78df;
        src75 <= 16'h22f0;
        src76 <= 16'h5443;
        src77 <= 16'hf78a;
        src78 <= 16'h9817;
        src79 <= 16'h4fe3;
        src80 <= 16'h930f;
        src81 <= 16'h5c05;
        src82 <= 16'hf64a;
        src83 <= 16'h4c66;
        src84 <= 16'hb122;
        src85 <= 16'hbfb3;
        src86 <= 16'hcb90;
        src87 <= 16'h416b;
        src88 <= 16'hd2a2;
        src89 <= 16'hff3b;
        src90 <= 16'hcb30;
        src91 <= 16'h3bde;
        src92 <= 16'hf098;
        src93 <= 16'hf766;
        src94 <= 16'h7c90;
        src95 <= 16'h4239;
        src96 <= 16'h1dd7;
        src97 <= 16'h13c1;
        src98 <= 16'hbe4c;
        src99 <= 16'hbbab;
        src100 <= 16'hfb59;
        src101 <= 16'h1baf;
        src102 <= 16'hc53;
        src103 <= 16'hac3f;
        src104 <= 16'h29ba;
        src105 <= 16'hd37;
        src106 <= 16'hf44;
        src107 <= 16'hcdbb;
        src108 <= 16'hb92e;
        src109 <= 16'hc6c4;
        src110 <= 16'hc348;
        src111 <= 16'hede7;
        src112 <= 16'hdc04;
        src113 <= 16'he03e;
        src114 <= 16'h2825;
        src115 <= 16'hbc95;
        src116 <= 16'hb693;
        src117 <= 16'h884e;
        src118 <= 16'hfc2f;
        src119 <= 16'h3032;
        src120 <= 16'he7b9;
        src121 <= 16'h1903;
        src122 <= 16'h56a6;
        src123 <= 16'h2424;
        src124 <= 16'h9389;
        src125 <= 16'h284;
        src126 <= 16'h7317;
        src127 <= 16'h1e5a;
        src128 <= 16'hce5e;
        src129 <= 16'h4426;
        src130 <= 16'h591;
        src131 <= 16'h59c1;
        src132 <= 16'h3be3;
        src133 <= 16'hd5e7;
        src134 <= 16'hf828;
        src135 <= 16'haac8;
        src136 <= 16'h5935;
        src137 <= 16'h3324;
        src138 <= 16'h60c6;
        src139 <= 16'h5a94;
        src140 <= 16'h7857;
        src141 <= 16'h9d5d;
        src142 <= 16'hb94f;
        src143 <= 16'h57cf;
        src144 <= 16'hbeb1;
        src145 <= 16'h17c8;
        src146 <= 16'hf6c3;
        src147 <= 16'h8079;
        src148 <= 16'h1c10;
        src149 <= 16'ha76c;
        src150 <= 16'h5dbd;
        src151 <= 16'ha1f0;
        src152 <= 16'h7cd3;
        src153 <= 16'h7872;
        src154 <= 16'h87ac;
        src155 <= 16'h8340;
        src156 <= 16'h6647;
        src157 <= 16'h7841;
        src158 <= 16'h4a26;
        src159 <= 16'hc16c;
        src160 <= 16'h6078;
        src161 <= 16'hf2a4;
        exp <= 24'h547d22;
        #1
        src0 <= 16'h7ccb;
        src1 <= 16'hc97e;
        src2 <= 16'ha93;
        src3 <= 16'h302;
        src4 <= 16'h674c;
        src5 <= 16'hfc0f;
        src6 <= 16'h83c3;
        src7 <= 16'h528a;
        src8 <= 16'h2846;
        src9 <= 16'h8ab;
        src10 <= 16'ha995;
        src11 <= 16'hcfde;
        src12 <= 16'h1ac7;
        src13 <= 16'h4825;
        src14 <= 16'h4d68;
        src15 <= 16'hea9d;
        src16 <= 16'h2674;
        src17 <= 16'h980f;
        src18 <= 16'h9eb2;
        src19 <= 16'h8308;
        src20 <= 16'h62af;
        src21 <= 16'h4889;
        src22 <= 16'hf050;
        src23 <= 16'h5fc4;
        src24 <= 16'h3402;
        src25 <= 16'he9d3;
        src26 <= 16'h334e;
        src27 <= 16'hf677;
        src28 <= 16'h55b4;
        src29 <= 16'he71f;
        src30 <= 16'haad7;
        src31 <= 16'h55bf;
        src32 <= 16'ha1fd;
        src33 <= 16'h7023;
        src34 <= 16'h5bf2;
        src35 <= 16'hdf2d;
        src36 <= 16'h5811;
        src37 <= 16'hf75;
        src38 <= 16'he745;
        src39 <= 16'hb857;
        src40 <= 16'h2c2d;
        src41 <= 16'he06c;
        src42 <= 16'h45b4;
        src43 <= 16'hec4a;
        src44 <= 16'h9c34;
        src45 <= 16'h90d;
        src46 <= 16'h722d;
        src47 <= 16'hbe4d;
        src48 <= 16'h413f;
        src49 <= 16'he255;
        src50 <= 16'h8332;
        src51 <= 16'h6da3;
        src52 <= 16'hbf3e;
        src53 <= 16'hb25b;
        src54 <= 16'h5619;
        src55 <= 16'h8c9e;
        src56 <= 16'hbaa8;
        src57 <= 16'h71f3;
        src58 <= 16'ha4de;
        src59 <= 16'h1099;
        src60 <= 16'hfc51;
        src61 <= 16'hbf38;
        src62 <= 16'h4eb6;
        src63 <= 16'hb8ff;
        src64 <= 16'h3a39;
        src65 <= 16'h47be;
        src66 <= 16'h3143;
        src67 <= 16'h4448;
        src68 <= 16'h34f5;
        src69 <= 16'hdd7a;
        src70 <= 16'h2db5;
        src71 <= 16'hfa8e;
        src72 <= 16'h1dba;
        src73 <= 16'ha83f;
        src74 <= 16'h98a4;
        src75 <= 16'hf280;
        src76 <= 16'hb5b4;
        src77 <= 16'haf3c;
        src78 <= 16'h497a;
        src79 <= 16'hcc41;
        src80 <= 16'hd604;
        src81 <= 16'heb73;
        src82 <= 16'ha796;
        src83 <= 16'h708b;
        src84 <= 16'hec46;
        src85 <= 16'h76a7;
        src86 <= 16'h70ca;
        src87 <= 16'he79d;
        src88 <= 16'h7035;
        src89 <= 16'h57e0;
        src90 <= 16'ha606;
        src91 <= 16'h778a;
        src92 <= 16'h9714;
        src93 <= 16'h35a7;
        src94 <= 16'h4695;
        src95 <= 16'h80af;
        src96 <= 16'h747;
        src97 <= 16'hec7c;
        src98 <= 16'h1850;
        src99 <= 16'h88b6;
        src100 <= 16'hb5aa;
        src101 <= 16'hca6c;
        src102 <= 16'h1e94;
        src103 <= 16'h34fd;
        src104 <= 16'h925c;
        src105 <= 16'hbc86;
        src106 <= 16'h90be;
        src107 <= 16'he461;
        src108 <= 16'h913e;
        src109 <= 16'hceb7;
        src110 <= 16'hb97e;
        src111 <= 16'h40b2;
        src112 <= 16'h5acb;
        src113 <= 16'h5261;
        src114 <= 16'hd3bb;
        src115 <= 16'h7df6;
        src116 <= 16'ha03;
        src117 <= 16'h43d7;
        src118 <= 16'h7a47;
        src119 <= 16'h6f60;
        src120 <= 16'h827d;
        src121 <= 16'hb8e8;
        src122 <= 16'h1053;
        src123 <= 16'hca2d;
        src124 <= 16'h1942;
        src125 <= 16'h42d6;
        src126 <= 16'h39de;
        src127 <= 16'h2657;
        src128 <= 16'hf92d;
        src129 <= 16'h95eb;
        src130 <= 16'h6788;
        src131 <= 16'h727b;
        src132 <= 16'hc666;
        src133 <= 16'h3839;
        src134 <= 16'hbf73;
        src135 <= 16'hec4d;
        src136 <= 16'he500;
        src137 <= 16'h9137;
        src138 <= 16'hbfc6;
        src139 <= 16'h58d6;
        src140 <= 16'ha6c8;
        src141 <= 16'h5177;
        src142 <= 16'h80ea;
        src143 <= 16'hce89;
        src144 <= 16'hd661;
        src145 <= 16'h905c;
        src146 <= 16'h3d6c;
        src147 <= 16'hff9b;
        src148 <= 16'h88c4;
        src149 <= 16'hd7d8;
        src150 <= 16'h2bbd;
        src151 <= 16'h63fe;
        src152 <= 16'hbedb;
        src153 <= 16'hdd61;
        src154 <= 16'hbe92;
        src155 <= 16'h9393;
        src156 <= 16'ha181;
        src157 <= 16'hc3b4;
        src158 <= 16'h2b06;
        src159 <= 16'h30c7;
        src160 <= 16'h6cf4;
        src161 <= 16'h7037;
        exp <= 24'h54507d;
        #1
        src0 <= 16'h297d;
        src1 <= 16'hf727;
        src2 <= 16'h6879;
        src3 <= 16'h2933;
        src4 <= 16'hdc7b;
        src5 <= 16'h43f5;
        src6 <= 16'h80d1;
        src7 <= 16'h7680;
        src8 <= 16'hbad6;
        src9 <= 16'h4a10;
        src10 <= 16'h539e;
        src11 <= 16'hb2b;
        src12 <= 16'h60e5;
        src13 <= 16'h508b;
        src14 <= 16'h5258;
        src15 <= 16'h6b17;
        src16 <= 16'hc242;
        src17 <= 16'h1a28;
        src18 <= 16'h33e9;
        src19 <= 16'ha9cf;
        src20 <= 16'he89f;
        src21 <= 16'hb15f;
        src22 <= 16'hfcd;
        src23 <= 16'h8f2c;
        src24 <= 16'h1450;
        src25 <= 16'h4e7f;
        src26 <= 16'h18bc;
        src27 <= 16'h317d;
        src28 <= 16'h4ef8;
        src29 <= 16'h52e7;
        src30 <= 16'h8cc1;
        src31 <= 16'hd79b;
        src32 <= 16'h9e17;
        src33 <= 16'h540e;
        src34 <= 16'h294;
        src35 <= 16'hff27;
        src36 <= 16'hc6ed;
        src37 <= 16'hd0b0;
        src38 <= 16'hc486;
        src39 <= 16'h7cb6;
        src40 <= 16'h23e2;
        src41 <= 16'h7e6d;
        src42 <= 16'hacb2;
        src43 <= 16'ha6bf;
        src44 <= 16'hdcfa;
        src45 <= 16'hda78;
        src46 <= 16'h3f30;
        src47 <= 16'h83d0;
        src48 <= 16'h12d8;
        src49 <= 16'hb151;
        src50 <= 16'h5b72;
        src51 <= 16'h516e;
        src52 <= 16'hf29;
        src53 <= 16'h1c23;
        src54 <= 16'h2bff;
        src55 <= 16'h730b;
        src56 <= 16'ha984;
        src57 <= 16'h40ae;
        src58 <= 16'hbfec;
        src59 <= 16'hb716;
        src60 <= 16'he34f;
        src61 <= 16'hdc2b;
        src62 <= 16'h84d1;
        src63 <= 16'h5d2c;
        src64 <= 16'hf28e;
        src65 <= 16'hcf1d;
        src66 <= 16'hf90c;
        src67 <= 16'h547d;
        src68 <= 16'h1c07;
        src69 <= 16'hcae1;
        src70 <= 16'hd739;
        src71 <= 16'h4983;
        src72 <= 16'h5c10;
        src73 <= 16'h821c;
        src74 <= 16'h513c;
        src75 <= 16'hcbd2;
        src76 <= 16'ha502;
        src77 <= 16'hb40c;
        src78 <= 16'h20fd;
        src79 <= 16'h73ce;
        src80 <= 16'hd9db;
        src81 <= 16'h4e32;
        src82 <= 16'hdb2;
        src83 <= 16'h31cb;
        src84 <= 16'h77b7;
        src85 <= 16'ha3b1;
        src86 <= 16'hdae9;
        src87 <= 16'hea3a;
        src88 <= 16'h30fb;
        src89 <= 16'h5214;
        src90 <= 16'h9f55;
        src91 <= 16'h4d55;
        src92 <= 16'h68a0;
        src93 <= 16'h6e6a;
        src94 <= 16'hd7de;
        src95 <= 16'h4947;
        src96 <= 16'hd780;
        src97 <= 16'hce65;
        src98 <= 16'hc313;
        src99 <= 16'h56e2;
        src100 <= 16'ha02d;
        src101 <= 16'h567f;
        src102 <= 16'haec0;
        src103 <= 16'h6897;
        src104 <= 16'h2675;
        src105 <= 16'hd7f0;
        src106 <= 16'h986f;
        src107 <= 16'hc480;
        src108 <= 16'h1ab2;
        src109 <= 16'haeb7;
        src110 <= 16'h2f8d;
        src111 <= 16'h2f34;
        src112 <= 16'h507a;
        src113 <= 16'h678e;
        src114 <= 16'h3ae3;
        src115 <= 16'h7299;
        src116 <= 16'ha86f;
        src117 <= 16'hc358;
        src118 <= 16'hb900;
        src119 <= 16'hd488;
        src120 <= 16'h39ca;
        src121 <= 16'h2122;
        src122 <= 16'hc22d;
        src123 <= 16'hb253;
        src124 <= 16'h7b91;
        src125 <= 16'h171d;
        src126 <= 16'hf80;
        src127 <= 16'h7e21;
        src128 <= 16'hd2f6;
        src129 <= 16'h46d1;
        src130 <= 16'hb695;
        src131 <= 16'hfa02;
        src132 <= 16'h318;
        src133 <= 16'haa95;
        src134 <= 16'h3f0e;
        src135 <= 16'h924;
        src136 <= 16'h57b1;
        src137 <= 16'hba00;
        src138 <= 16'h1902;
        src139 <= 16'h54c2;
        src140 <= 16'h3bd6;
        src141 <= 16'h8e5d;
        src142 <= 16'hfa34;
        src143 <= 16'h4f31;
        src144 <= 16'h4f0d;
        src145 <= 16'hd702;
        src146 <= 16'h7803;
        src147 <= 16'h698f;
        src148 <= 16'hdf68;
        src149 <= 16'h46f6;
        src150 <= 16'hd01b;
        src151 <= 16'hdfaf;
        src152 <= 16'he23f;
        src153 <= 16'h3a34;
        src154 <= 16'hf981;
        src155 <= 16'h1b7;
        src156 <= 16'he52d;
        src157 <= 16'h8993;
        src158 <= 16'hc72c;
        src159 <= 16'h1ce0;
        src160 <= 16'h38ef;
        src161 <= 16'h3519;
        exp <= 24'h4f1753;
        #1
        src0 <= 16'hf94;
        src1 <= 16'hb240;
        src2 <= 16'h9a77;
        src3 <= 16'hc1e4;
        src4 <= 16'he682;
        src5 <= 16'hd9f2;
        src6 <= 16'h88c2;
        src7 <= 16'h4f8a;
        src8 <= 16'hcf43;
        src9 <= 16'h26b9;
        src10 <= 16'hf50c;
        src11 <= 16'h8d33;
        src12 <= 16'h805c;
        src13 <= 16'h1b61;
        src14 <= 16'hef0;
        src15 <= 16'ha0cf;
        src16 <= 16'h92ea;
        src17 <= 16'h3f3e;
        src18 <= 16'hfa3d;
        src19 <= 16'h59ec;
        src20 <= 16'hda2b;
        src21 <= 16'h3669;
        src22 <= 16'hd76a;
        src23 <= 16'h3903;
        src24 <= 16'he632;
        src25 <= 16'hcf0a;
        src26 <= 16'hfbc3;
        src27 <= 16'hdfad;
        src28 <= 16'hd07a;
        src29 <= 16'he998;
        src30 <= 16'hfacf;
        src31 <= 16'h9d68;
        src32 <= 16'he6fb;
        src33 <= 16'h7e46;
        src34 <= 16'h38e2;
        src35 <= 16'h76b9;
        src36 <= 16'h2526;
        src37 <= 16'hfedf;
        src38 <= 16'h526c;
        src39 <= 16'hbd55;
        src40 <= 16'h186c;
        src41 <= 16'h590;
        src42 <= 16'h1eb8;
        src43 <= 16'h8ecb;
        src44 <= 16'h1566;
        src45 <= 16'h1bca;
        src46 <= 16'h17eb;
        src47 <= 16'h30c9;
        src48 <= 16'h40e6;
        src49 <= 16'h946e;
        src50 <= 16'h986;
        src51 <= 16'h7fd;
        src52 <= 16'h79c2;
        src53 <= 16'h42f9;
        src54 <= 16'h1021;
        src55 <= 16'hc84b;
        src56 <= 16'h2ebe;
        src57 <= 16'h1993;
        src58 <= 16'hb35d;
        src59 <= 16'hce64;
        src60 <= 16'h77d7;
        src61 <= 16'h3d57;
        src62 <= 16'hc7ae;
        src63 <= 16'h17ac;
        src64 <= 16'h1f21;
        src65 <= 16'h3804;
        src66 <= 16'hb28b;
        src67 <= 16'h6c75;
        src68 <= 16'h7576;
        src69 <= 16'ha634;
        src70 <= 16'hb4f4;
        src71 <= 16'hf1a3;
        src72 <= 16'hc173;
        src73 <= 16'hadc7;
        src74 <= 16'h9dcc;
        src75 <= 16'he4a6;
        src76 <= 16'h6851;
        src77 <= 16'h8c3;
        src78 <= 16'h51ff;
        src79 <= 16'h4548;
        src80 <= 16'hbb10;
        src81 <= 16'he12a;
        src82 <= 16'h65fc;
        src83 <= 16'hddd5;
        src84 <= 16'h3ee2;
        src85 <= 16'h67bf;
        src86 <= 16'h9772;
        src87 <= 16'ha02b;
        src88 <= 16'h587d;
        src89 <= 16'hbcbf;
        src90 <= 16'h5667;
        src91 <= 16'h5196;
        src92 <= 16'hc680;
        src93 <= 16'hb0df;
        src94 <= 16'h7d4f;
        src95 <= 16'h81f5;
        src96 <= 16'h716e;
        src97 <= 16'hb4e5;
        src98 <= 16'h6e3;
        src99 <= 16'hef11;
        src100 <= 16'hffe0;
        src101 <= 16'h16d3;
        src102 <= 16'h89fe;
        src103 <= 16'hd386;
        src104 <= 16'ha97;
        src105 <= 16'h9202;
        src106 <= 16'h4081;
        src107 <= 16'h5a26;
        src108 <= 16'hb7f5;
        src109 <= 16'h4cba;
        src110 <= 16'ha055;
        src111 <= 16'h32a7;
        src112 <= 16'h2f1b;
        src113 <= 16'h16c0;
        src114 <= 16'h1a0c;
        src115 <= 16'ha7eb;
        src116 <= 16'h4774;
        src117 <= 16'h8222;
        src118 <= 16'h9962;
        src119 <= 16'hae01;
        src120 <= 16'h44bb;
        src121 <= 16'hbcaf;
        src122 <= 16'h25b3;
        src123 <= 16'h956e;
        src124 <= 16'hb3d1;
        src125 <= 16'h9d03;
        src126 <= 16'h4890;
        src127 <= 16'ha7e9;
        src128 <= 16'h7c87;
        src129 <= 16'hcb55;
        src130 <= 16'hf774;
        src131 <= 16'h5e30;
        src132 <= 16'h82fe;
        src133 <= 16'h13fa;
        src134 <= 16'h629a;
        src135 <= 16'h12b1;
        src136 <= 16'hd66;
        src137 <= 16'hd6e;
        src138 <= 16'h2fe8;
        src139 <= 16'hc6af;
        src140 <= 16'h32f7;
        src141 <= 16'h3e1;
        src142 <= 16'hdf12;
        src143 <= 16'h4d6b;
        src144 <= 16'h1582;
        src145 <= 16'hfa82;
        src146 <= 16'hc9e9;
        src147 <= 16'hf433;
        src148 <= 16'h755;
        src149 <= 16'h327d;
        src150 <= 16'h7bd5;
        src151 <= 16'hbb63;
        src152 <= 16'h6f9f;
        src153 <= 16'hd5d3;
        src154 <= 16'he1af;
        src155 <= 16'hbcb4;
        src156 <= 16'h8256;
        src157 <= 16'hd12e;
        src158 <= 16'h252e;
        src159 <= 16'ha024;
        src160 <= 16'h1f16;
        src161 <= 16'hff67;
        exp <= 24'h4f60fd;
        #1
        src0 <= 16'ha89f;
        src1 <= 16'h4159;
        src2 <= 16'h7209;
        src3 <= 16'h67db;
        src4 <= 16'hb65;
        src5 <= 16'hc1ff;
        src6 <= 16'h1c43;
        src7 <= 16'h39e7;
        src8 <= 16'hcc39;
        src9 <= 16'h5884;
        src10 <= 16'h5bdc;
        src11 <= 16'h8b84;
        src12 <= 16'h1263;
        src13 <= 16'h5d2c;
        src14 <= 16'h15ec;
        src15 <= 16'h2f13;
        src16 <= 16'hc255;
        src17 <= 16'heec8;
        src18 <= 16'hcc36;
        src19 <= 16'h268b;
        src20 <= 16'hc057;
        src21 <= 16'h4aef;
        src22 <= 16'hce11;
        src23 <= 16'hb918;
        src24 <= 16'h5140;
        src25 <= 16'h9701;
        src26 <= 16'hf8cf;
        src27 <= 16'hf904;
        src28 <= 16'hded4;
        src29 <= 16'h582d;
        src30 <= 16'h5712;
        src31 <= 16'h4259;
        src32 <= 16'h98bc;
        src33 <= 16'h52a0;
        src34 <= 16'h9c0d;
        src35 <= 16'hd4ba;
        src36 <= 16'h249b;
        src37 <= 16'hb322;
        src38 <= 16'hf052;
        src39 <= 16'h2930;
        src40 <= 16'h8dea;
        src41 <= 16'h3565;
        src42 <= 16'h4802;
        src43 <= 16'hc68d;
        src44 <= 16'hd00f;
        src45 <= 16'h8a7f;
        src46 <= 16'h129c;
        src47 <= 16'h9e4a;
        src48 <= 16'h6b9c;
        src49 <= 16'h6f56;
        src50 <= 16'he084;
        src51 <= 16'hb3e1;
        src52 <= 16'hb765;
        src53 <= 16'h656e;
        src54 <= 16'h3f4c;
        src55 <= 16'h7277;
        src56 <= 16'h729d;
        src57 <= 16'hc02;
        src58 <= 16'h701f;
        src59 <= 16'he72;
        src60 <= 16'h2455;
        src61 <= 16'h1428;
        src62 <= 16'h4991;
        src63 <= 16'h53a4;
        src64 <= 16'h861c;
        src65 <= 16'h48e6;
        src66 <= 16'h797c;
        src67 <= 16'hafd3;
        src68 <= 16'h49d8;
        src69 <= 16'hfe0;
        src70 <= 16'h37f5;
        src71 <= 16'he626;
        src72 <= 16'he202;
        src73 <= 16'hba48;
        src74 <= 16'hd19a;
        src75 <= 16'he8e;
        src76 <= 16'hbd53;
        src77 <= 16'h24dd;
        src78 <= 16'hb5b0;
        src79 <= 16'hf48d;
        src80 <= 16'h5743;
        src81 <= 16'h5ab3;
        src82 <= 16'h7b47;
        src83 <= 16'h746d;
        src84 <= 16'hd71b;
        src85 <= 16'h6181;
        src86 <= 16'hfcf7;
        src87 <= 16'h4813;
        src88 <= 16'h1d6b;
        src89 <= 16'h5ed3;
        src90 <= 16'h782;
        src91 <= 16'h7b8d;
        src92 <= 16'h84a9;
        src93 <= 16'h13f7;
        src94 <= 16'h499;
        src95 <= 16'h930a;
        src96 <= 16'hf13d;
        src97 <= 16'h1d6f;
        src98 <= 16'he3f0;
        src99 <= 16'hfa66;
        src100 <= 16'h2ca1;
        src101 <= 16'h6aa0;
        src102 <= 16'hd99;
        src103 <= 16'hbfc1;
        src104 <= 16'hbace;
        src105 <= 16'h5663;
        src106 <= 16'h38b5;
        src107 <= 16'h7915;
        src108 <= 16'he6c4;
        src109 <= 16'hc972;
        src110 <= 16'hc8e9;
        src111 <= 16'h1e89;
        src112 <= 16'hd261;
        src113 <= 16'h6ef2;
        src114 <= 16'h4dc2;
        src115 <= 16'hfd8a;
        src116 <= 16'hd5c3;
        src117 <= 16'h4ab2;
        src118 <= 16'hdd28;
        src119 <= 16'hf539;
        src120 <= 16'h496a;
        src121 <= 16'h4da9;
        src122 <= 16'h15f7;
        src123 <= 16'h647d;
        src124 <= 16'h447f;
        src125 <= 16'h4c63;
        src126 <= 16'h6cf5;
        src127 <= 16'h3742;
        src128 <= 16'hb85d;
        src129 <= 16'hfa6e;
        src130 <= 16'ha71d;
        src131 <= 16'h7d6d;
        src132 <= 16'h8981;
        src133 <= 16'hb2dc;
        src134 <= 16'h665b;
        src135 <= 16'h186e;
        src136 <= 16'h90e0;
        src137 <= 16'hd1c7;
        src138 <= 16'hcbc3;
        src139 <= 16'h9f2a;
        src140 <= 16'h408;
        src141 <= 16'h5a1a;
        src142 <= 16'hc640;
        src143 <= 16'h9d96;
        src144 <= 16'h195f;
        src145 <= 16'h3e5;
        src146 <= 16'hfc72;
        src147 <= 16'hc42e;
        src148 <= 16'h8147;
        src149 <= 16'ha342;
        src150 <= 16'h493e;
        src151 <= 16'hfd50;
        src152 <= 16'h9ef7;
        src153 <= 16'h5612;
        src154 <= 16'h3960;
        src155 <= 16'h2b28;
        src156 <= 16'hccc4;
        src157 <= 16'h19ac;
        src158 <= 16'h9f18;
        src159 <= 16'h23cf;
        src160 <= 16'hf53c;
        src161 <= 16'hb995;
        exp <= 24'h4f1b58;
        #1
        src0 <= 16'h5dca;
        src1 <= 16'h543d;
        src2 <= 16'h3790;
        src3 <= 16'h7867;
        src4 <= 16'h6cb8;
        src5 <= 16'hdd30;
        src6 <= 16'h2e38;
        src7 <= 16'hb5c2;
        src8 <= 16'h4f85;
        src9 <= 16'hfd12;
        src10 <= 16'h1902;
        src11 <= 16'h4e40;
        src12 <= 16'hd8d3;
        src13 <= 16'h41af;
        src14 <= 16'hbe8f;
        src15 <= 16'hba22;
        src16 <= 16'hba43;
        src17 <= 16'hc30e;
        src18 <= 16'h8b05;
        src19 <= 16'hadf;
        src20 <= 16'hc198;
        src21 <= 16'h4021;
        src22 <= 16'h5388;
        src23 <= 16'h418;
        src24 <= 16'hb984;
        src25 <= 16'hdacb;
        src26 <= 16'ha9a9;
        src27 <= 16'h5693;
        src28 <= 16'h885f;
        src29 <= 16'he585;
        src30 <= 16'h7d6f;
        src31 <= 16'he188;
        src32 <= 16'h8501;
        src33 <= 16'hb05;
        src34 <= 16'ha5c6;
        src35 <= 16'h9262;
        src36 <= 16'h6d05;
        src37 <= 16'hc378;
        src38 <= 16'h4d20;
        src39 <= 16'hed8c;
        src40 <= 16'hd61a;
        src41 <= 16'h70be;
        src42 <= 16'hf69e;
        src43 <= 16'h3b05;
        src44 <= 16'h9754;
        src45 <= 16'ha557;
        src46 <= 16'h7bd5;
        src47 <= 16'h9906;
        src48 <= 16'hc48f;
        src49 <= 16'h9441;
        src50 <= 16'h6714;
        src51 <= 16'h1022;
        src52 <= 16'h2258;
        src53 <= 16'hafb9;
        src54 <= 16'haa0a;
        src55 <= 16'h3a4;
        src56 <= 16'h3257;
        src57 <= 16'h1521;
        src58 <= 16'h2c68;
        src59 <= 16'hce60;
        src60 <= 16'hbe18;
        src61 <= 16'he7f4;
        src62 <= 16'h66da;
        src63 <= 16'h18de;
        src64 <= 16'hd7fc;
        src65 <= 16'hc3d8;
        src66 <= 16'h120;
        src67 <= 16'hf478;
        src68 <= 16'h1196;
        src69 <= 16'h3f23;
        src70 <= 16'h3d59;
        src71 <= 16'h9a12;
        src72 <= 16'h45d9;
        src73 <= 16'h1115;
        src74 <= 16'h53ca;
        src75 <= 16'hea2c;
        src76 <= 16'h4d9;
        src77 <= 16'hbaf7;
        src78 <= 16'h1312;
        src79 <= 16'h2a38;
        src80 <= 16'h4a16;
        src81 <= 16'h4654;
        src82 <= 16'h9bbf;
        src83 <= 16'h5fb2;
        src84 <= 16'hc6c3;
        src85 <= 16'h88ef;
        src86 <= 16'hdcbb;
        src87 <= 16'h1f50;
        src88 <= 16'h183f;
        src89 <= 16'hdbb6;
        src90 <= 16'h8a00;
        src91 <= 16'h34ad;
        src92 <= 16'hc3ae;
        src93 <= 16'h957a;
        src94 <= 16'h611e;
        src95 <= 16'hb9da;
        src96 <= 16'h8ce6;
        src97 <= 16'hd3f3;
        src98 <= 16'ha769;
        src99 <= 16'hc8eb;
        src100 <= 16'hb011;
        src101 <= 16'h51f0;
        src102 <= 16'h401;
        src103 <= 16'h83fc;
        src104 <= 16'h9c41;
        src105 <= 16'h8f29;
        src106 <= 16'h15d;
        src107 <= 16'h370f;
        src108 <= 16'hb9bb;
        src109 <= 16'haf96;
        src110 <= 16'he203;
        src111 <= 16'hc35a;
        src112 <= 16'h4973;
        src113 <= 16'h850c;
        src114 <= 16'h460c;
        src115 <= 16'h68f6;
        src116 <= 16'h800d;
        src117 <= 16'h384d;
        src118 <= 16'hb138;
        src119 <= 16'h20f6;
        src120 <= 16'h6048;
        src121 <= 16'haf8;
        src122 <= 16'h8b86;
        src123 <= 16'hc6df;
        src124 <= 16'h60ce;
        src125 <= 16'h9022;
        src126 <= 16'h458;
        src127 <= 16'h6732;
        src128 <= 16'hb177;
        src129 <= 16'h5125;
        src130 <= 16'h30f5;
        src131 <= 16'h63bc;
        src132 <= 16'h5197;
        src133 <= 16'h998f;
        src134 <= 16'h4064;
        src135 <= 16'h15d8;
        src136 <= 16'he319;
        src137 <= 16'hf8a4;
        src138 <= 16'hae18;
        src139 <= 16'hdd9c;
        src140 <= 16'h7dc9;
        src141 <= 16'h241d;
        src142 <= 16'h92bb;
        src143 <= 16'he506;
        src144 <= 16'h9953;
        src145 <= 16'h2f3c;
        src146 <= 16'he5ee;
        src147 <= 16'h7edb;
        src148 <= 16'h8c78;
        src149 <= 16'h9b4;
        src150 <= 16'hde34;
        src151 <= 16'h585b;
        src152 <= 16'h3b3c;
        src153 <= 16'h96cb;
        src154 <= 16'h4ec6;
        src155 <= 16'hae0b;
        src156 <= 16'h7610;
        src157 <= 16'h8212;
        src158 <= 16'hd621;
        src159 <= 16'h1e1f;
        src160 <= 16'ha382;
        src161 <= 16'hce26;
        exp <= 24'h4f147c;
        #1
        src0 <= 16'h7e5a;
        src1 <= 16'hd275;
        src2 <= 16'h9f2;
        src3 <= 16'h3c72;
        src4 <= 16'hcffb;
        src5 <= 16'h63a0;
        src6 <= 16'h63f5;
        src7 <= 16'hc363;
        src8 <= 16'hc1bb;
        src9 <= 16'h7a0f;
        src10 <= 16'he8a4;
        src11 <= 16'hef8;
        src12 <= 16'h3178;
        src13 <= 16'hcaeb;
        src14 <= 16'h5ddc;
        src15 <= 16'hf597;
        src16 <= 16'h1f66;
        src17 <= 16'hd42a;
        src18 <= 16'hd235;
        src19 <= 16'h9c78;
        src20 <= 16'h1713;
        src21 <= 16'hf01e;
        src22 <= 16'ha85d;
        src23 <= 16'he89b;
        src24 <= 16'hf3d0;
        src25 <= 16'h963f;
        src26 <= 16'h3b7c;
        src27 <= 16'h50b;
        src28 <= 16'h12fe;
        src29 <= 16'h4c5e;
        src30 <= 16'h51ed;
        src31 <= 16'he5ef;
        src32 <= 16'he1c0;
        src33 <= 16'hcba9;
        src34 <= 16'h8494;
        src35 <= 16'h2e0d;
        src36 <= 16'h57ca;
        src37 <= 16'h8335;
        src38 <= 16'hd8f3;
        src39 <= 16'h4696;
        src40 <= 16'h322e;
        src41 <= 16'hfd07;
        src42 <= 16'h8a20;
        src43 <= 16'h551e;
        src44 <= 16'hca8;
        src45 <= 16'hb53;
        src46 <= 16'h4fc7;
        src47 <= 16'h6acc;
        src48 <= 16'hfa77;
        src49 <= 16'h6d01;
        src50 <= 16'hc951;
        src51 <= 16'h2218;
        src52 <= 16'h9f97;
        src53 <= 16'h9a68;
        src54 <= 16'h884a;
        src55 <= 16'h40c5;
        src56 <= 16'hee31;
        src57 <= 16'h4eec;
        src58 <= 16'h5e5b;
        src59 <= 16'h532c;
        src60 <= 16'h8aba;
        src61 <= 16'h5b2c;
        src62 <= 16'h612c;
        src63 <= 16'h7330;
        src64 <= 16'h4924;
        src65 <= 16'hc79f;
        src66 <= 16'h24de;
        src67 <= 16'he984;
        src68 <= 16'h4ecd;
        src69 <= 16'h3592;
        src70 <= 16'h519f;
        src71 <= 16'hba00;
        src72 <= 16'h23f1;
        src73 <= 16'hc93e;
        src74 <= 16'hcd27;
        src75 <= 16'he257;
        src76 <= 16'h1351;
        src77 <= 16'h2fa9;
        src78 <= 16'hb93c;
        src79 <= 16'he83;
        src80 <= 16'hb61a;
        src81 <= 16'h6713;
        src82 <= 16'h8f93;
        src83 <= 16'h5219;
        src84 <= 16'hf10;
        src85 <= 16'hc53f;
        src86 <= 16'h170a;
        src87 <= 16'h63cc;
        src88 <= 16'h63b9;
        src89 <= 16'h3144;
        src90 <= 16'h3535;
        src91 <= 16'h7407;
        src92 <= 16'hfe91;
        src93 <= 16'hcd5c;
        src94 <= 16'h7a72;
        src95 <= 16'he88a;
        src96 <= 16'h462e;
        src97 <= 16'hf784;
        src98 <= 16'h4c95;
        src99 <= 16'h64ef;
        src100 <= 16'hccb1;
        src101 <= 16'h79c1;
        src102 <= 16'h2966;
        src103 <= 16'hec99;
        src104 <= 16'ha0c7;
        src105 <= 16'hc5a8;
        src106 <= 16'he04;
        src107 <= 16'h9e9b;
        src108 <= 16'h1925;
        src109 <= 16'h7209;
        src110 <= 16'hd631;
        src111 <= 16'h465b;
        src112 <= 16'h5b52;
        src113 <= 16'h9702;
        src114 <= 16'h7db7;
        src115 <= 16'h8118;
        src116 <= 16'hce3f;
        src117 <= 16'hc733;
        src118 <= 16'ha1ae;
        src119 <= 16'h3d3d;
        src120 <= 16'hdb81;
        src121 <= 16'ha966;
        src122 <= 16'h7b57;
        src123 <= 16'h24f9;
        src124 <= 16'h77aa;
        src125 <= 16'h2c82;
        src126 <= 16'he6cb;
        src127 <= 16'h3972;
        src128 <= 16'h8036;
        src129 <= 16'ha894;
        src130 <= 16'h8f83;
        src131 <= 16'h894c;
        src132 <= 16'he7f2;
        src133 <= 16'hf2b7;
        src134 <= 16'h4aef;
        src135 <= 16'ha04d;
        src136 <= 16'h2bc0;
        src137 <= 16'hafa9;
        src138 <= 16'hb1f8;
        src139 <= 16'h8ace;
        src140 <= 16'ha03d;
        src141 <= 16'h7d90;
        src142 <= 16'hbdad;
        src143 <= 16'ha449;
        src144 <= 16'hf2e9;
        src145 <= 16'h8542;
        src146 <= 16'h9dc;
        src147 <= 16'hde07;
        src148 <= 16'hcdba;
        src149 <= 16'hdd1c;
        src150 <= 16'hf044;
        src151 <= 16'hfc4c;
        src152 <= 16'h8ce2;
        src153 <= 16'h6d7;
        src154 <= 16'h7ddb;
        src155 <= 16'h72e6;
        src156 <= 16'h7098;
        src157 <= 16'h7de3;
        src158 <= 16'hb17;
        src159 <= 16'h8a6c;
        src160 <= 16'hdbe9;
        src161 <= 16'hdc6;
        exp <= 24'h52fc41;
        #1
        src0 <= 16'h50b8;
        src1 <= 16'h5605;
        src2 <= 16'hb004;
        src3 <= 16'h8879;
        src4 <= 16'h4a67;
        src5 <= 16'h5061;
        src6 <= 16'hc5b5;
        src7 <= 16'h3acf;
        src8 <= 16'hf079;
        src9 <= 16'hf6ae;
        src10 <= 16'h8fea;
        src11 <= 16'hfb52;
        src12 <= 16'hfa85;
        src13 <= 16'h3a9d;
        src14 <= 16'h4b03;
        src15 <= 16'h1711;
        src16 <= 16'ha9ba;
        src17 <= 16'h16df;
        src18 <= 16'hca28;
        src19 <= 16'h97a2;
        src20 <= 16'h82ba;
        src21 <= 16'h3c69;
        src22 <= 16'h1e1b;
        src23 <= 16'hdd14;
        src24 <= 16'hb58a;
        src25 <= 16'hce4a;
        src26 <= 16'h3401;
        src27 <= 16'hce91;
        src28 <= 16'h7521;
        src29 <= 16'h449b;
        src30 <= 16'h66c;
        src31 <= 16'h6b3;
        src32 <= 16'ha592;
        src33 <= 16'h60e9;
        src34 <= 16'h9e73;
        src35 <= 16'h74e3;
        src36 <= 16'he863;
        src37 <= 16'had8e;
        src38 <= 16'h64bb;
        src39 <= 16'h990a;
        src40 <= 16'hd128;
        src41 <= 16'hd8bb;
        src42 <= 16'h25e3;
        src43 <= 16'h12dc;
        src44 <= 16'h5daa;
        src45 <= 16'h16c4;
        src46 <= 16'h29d6;
        src47 <= 16'h5553;
        src48 <= 16'he747;
        src49 <= 16'h36ec;
        src50 <= 16'hbbd3;
        src51 <= 16'h78de;
        src52 <= 16'hf243;
        src53 <= 16'hb439;
        src54 <= 16'hd9be;
        src55 <= 16'h3852;
        src56 <= 16'h3d14;
        src57 <= 16'hc4b2;
        src58 <= 16'h362;
        src59 <= 16'ha61b;
        src60 <= 16'h3a48;
        src61 <= 16'h4b8f;
        src62 <= 16'h3dd8;
        src63 <= 16'hbc2a;
        src64 <= 16'h1c2d;
        src65 <= 16'h697a;
        src66 <= 16'h1049;
        src67 <= 16'had6c;
        src68 <= 16'had6d;
        src69 <= 16'hb8cc;
        src70 <= 16'hffeb;
        src71 <= 16'h6158;
        src72 <= 16'h9d78;
        src73 <= 16'hceab;
        src74 <= 16'haf8;
        src75 <= 16'h2a4d;
        src76 <= 16'h50ca;
        src77 <= 16'h85bb;
        src78 <= 16'h5e8b;
        src79 <= 16'h6ef6;
        src80 <= 16'he29c;
        src81 <= 16'hce2d;
        src82 <= 16'h4610;
        src83 <= 16'h940;
        src84 <= 16'had0f;
        src85 <= 16'h7e13;
        src86 <= 16'h7ad3;
        src87 <= 16'he155;
        src88 <= 16'he536;
        src89 <= 16'he4d7;
        src90 <= 16'h100f;
        src91 <= 16'h92e5;
        src92 <= 16'h66e0;
        src93 <= 16'h6cd;
        src94 <= 16'h8e5d;
        src95 <= 16'h4380;
        src96 <= 16'h99ad;
        src97 <= 16'h7aa7;
        src98 <= 16'h54ce;
        src99 <= 16'hfc1b;
        src100 <= 16'h4a18;
        src101 <= 16'h71ae;
        src102 <= 16'hff6;
        src103 <= 16'h5812;
        src104 <= 16'hbf33;
        src105 <= 16'hb641;
        src106 <= 16'h8ab0;
        src107 <= 16'h2c9;
        src108 <= 16'h500b;
        src109 <= 16'hcdea;
        src110 <= 16'he45;
        src111 <= 16'h2076;
        src112 <= 16'h1f93;
        src113 <= 16'h941c;
        src114 <= 16'h50e4;
        src115 <= 16'hae45;
        src116 <= 16'ha0fd;
        src117 <= 16'h5467;
        src118 <= 16'h13c9;
        src119 <= 16'h6538;
        src120 <= 16'h6c30;
        src121 <= 16'hd086;
        src122 <= 16'h6b93;
        src123 <= 16'hd5f2;
        src124 <= 16'h5a5;
        src125 <= 16'h14a5;
        src126 <= 16'h6a92;
        src127 <= 16'hbe50;
        src128 <= 16'hbad;
        src129 <= 16'he0e4;
        src130 <= 16'h8276;
        src131 <= 16'h4717;
        src132 <= 16'h9919;
        src133 <= 16'h8567;
        src134 <= 16'hc223;
        src135 <= 16'h54be;
        src136 <= 16'h3a43;
        src137 <= 16'h84de;
        src138 <= 16'h1697;
        src139 <= 16'hfc36;
        src140 <= 16'hd871;
        src141 <= 16'h3f0b;
        src142 <= 16'hfedb;
        src143 <= 16'hf8e9;
        src144 <= 16'h22b6;
        src145 <= 16'h1d33;
        src146 <= 16'h36f5;
        src147 <= 16'h41c5;
        src148 <= 16'h546d;
        src149 <= 16'hd92;
        src150 <= 16'h90ad;
        src151 <= 16'h8e55;
        src152 <= 16'hbff4;
        src153 <= 16'h8e4f;
        src154 <= 16'hff26;
        src155 <= 16'h8fdd;
        src156 <= 16'hca12;
        src157 <= 16'hed3c;
        src158 <= 16'hb217;
        src159 <= 16'h6205;
        src160 <= 16'h2613;
        src161 <= 16'h5cda;
        exp <= 24'h4dd9cf;
        #1
        src0 <= 16'hd071;
        src1 <= 16'h63d9;
        src2 <= 16'h79e1;
        src3 <= 16'hed2c;
        src4 <= 16'h85a;
        src5 <= 16'h62de;
        src6 <= 16'hb48d;
        src7 <= 16'h2ade;
        src8 <= 16'h2b1e;
        src9 <= 16'h2660;
        src10 <= 16'h5842;
        src11 <= 16'h87f2;
        src12 <= 16'hba6e;
        src13 <= 16'h8490;
        src14 <= 16'h1826;
        src15 <= 16'ha79;
        src16 <= 16'hfb41;
        src17 <= 16'hb067;
        src18 <= 16'h9123;
        src19 <= 16'ha185;
        src20 <= 16'hf6ef;
        src21 <= 16'h11c2;
        src22 <= 16'he20b;
        src23 <= 16'h728f;
        src24 <= 16'ha869;
        src25 <= 16'h90fe;
        src26 <= 16'h2f16;
        src27 <= 16'h711d;
        src28 <= 16'h895c;
        src29 <= 16'h366f;
        src30 <= 16'h8485;
        src31 <= 16'h7d5d;
        src32 <= 16'hefcb;
        src33 <= 16'hc93e;
        src34 <= 16'h8eb1;
        src35 <= 16'h9d0c;
        src36 <= 16'haefb;
        src37 <= 16'haf5d;
        src38 <= 16'h5751;
        src39 <= 16'h9927;
        src40 <= 16'he81a;
        src41 <= 16'h7913;
        src42 <= 16'hbad2;
        src43 <= 16'h8ee2;
        src44 <= 16'h3200;
        src45 <= 16'h568a;
        src46 <= 16'h6869;
        src47 <= 16'h695f;
        src48 <= 16'h279;
        src49 <= 16'h7a20;
        src50 <= 16'h9b8c;
        src51 <= 16'h5e17;
        src52 <= 16'h3593;
        src53 <= 16'h24cf;
        src54 <= 16'h25a1;
        src55 <= 16'h47eb;
        src56 <= 16'h59cc;
        src57 <= 16'h3780;
        src58 <= 16'h401e;
        src59 <= 16'h9666;
        src60 <= 16'hbe32;
        src61 <= 16'hf2f5;
        src62 <= 16'hd503;
        src63 <= 16'hb834;
        src64 <= 16'h1c05;
        src65 <= 16'h2bcd;
        src66 <= 16'h6e03;
        src67 <= 16'h7727;
        src68 <= 16'h47d3;
        src69 <= 16'ha960;
        src70 <= 16'hbf12;
        src71 <= 16'h2f76;
        src72 <= 16'h43b6;
        src73 <= 16'hd883;
        src74 <= 16'hea19;
        src75 <= 16'h7705;
        src76 <= 16'hd795;
        src77 <= 16'h5bbd;
        src78 <= 16'h1b4;
        src79 <= 16'h282e;
        src80 <= 16'hd421;
        src81 <= 16'ha38e;
        src82 <= 16'h2d82;
        src83 <= 16'h368d;
        src84 <= 16'h592c;
        src85 <= 16'hf9c5;
        src86 <= 16'hd691;
        src87 <= 16'h11ac;
        src88 <= 16'h1e0a;
        src89 <= 16'h60d6;
        src90 <= 16'h8485;
        src91 <= 16'hb81c;
        src92 <= 16'h856d;
        src93 <= 16'h452;
        src94 <= 16'hb7f5;
        src95 <= 16'h22e0;
        src96 <= 16'h831f;
        src97 <= 16'h3efe;
        src98 <= 16'h34a7;
        src99 <= 16'hac6d;
        src100 <= 16'hb02;
        src101 <= 16'h7f69;
        src102 <= 16'h5d67;
        src103 <= 16'hfc48;
        src104 <= 16'h2fe0;
        src105 <= 16'hb8ea;
        src106 <= 16'hc4ee;
        src107 <= 16'hac0d;
        src108 <= 16'h71ec;
        src109 <= 16'h57f8;
        src110 <= 16'hc323;
        src111 <= 16'hcff2;
        src112 <= 16'haa1b;
        src113 <= 16'h88e9;
        src114 <= 16'hcd63;
        src115 <= 16'h6bcf;
        src116 <= 16'h9aa0;
        src117 <= 16'h60a9;
        src118 <= 16'haff2;
        src119 <= 16'h8929;
        src120 <= 16'h786d;
        src121 <= 16'h4ae9;
        src122 <= 16'he7e3;
        src123 <= 16'hc134;
        src124 <= 16'h79e9;
        src125 <= 16'h3d0a;
        src126 <= 16'hdc7e;
        src127 <= 16'hca58;
        src128 <= 16'h65e1;
        src129 <= 16'hcec8;
        src130 <= 16'h97f9;
        src131 <= 16'h5b7;
        src132 <= 16'h5541;
        src133 <= 16'hc5d0;
        src134 <= 16'h590e;
        src135 <= 16'h9e73;
        src136 <= 16'h5729;
        src137 <= 16'h3c7f;
        src138 <= 16'h5e5d;
        src139 <= 16'he087;
        src140 <= 16'ha08f;
        src141 <= 16'h8a29;
        src142 <= 16'hab4c;
        src143 <= 16'h3f09;
        src144 <= 16'hb632;
        src145 <= 16'he608;
        src146 <= 16'hb617;
        src147 <= 16'ha8f6;
        src148 <= 16'h926b;
        src149 <= 16'h270e;
        src150 <= 16'hb48d;
        src151 <= 16'h94c8;
        src152 <= 16'h2cd5;
        src153 <= 16'h25f1;
        src154 <= 16'hfd96;
        src155 <= 16'h7384;
        src156 <= 16'hc4e0;
        src157 <= 16'h2251;
        src158 <= 16'h5691;
        src159 <= 16'h253b;
        src160 <= 16'heb35;
        src161 <= 16'hbe6f;
        exp <= 24'h50cf82;
        #1
        src0 <= 16'h6374;
        src1 <= 16'h14bd;
        src2 <= 16'h4ea9;
        src3 <= 16'h2cd5;
        src4 <= 16'h9de2;
        src5 <= 16'h5daf;
        src6 <= 16'h7866;
        src7 <= 16'hefcb;
        src8 <= 16'h8b85;
        src9 <= 16'h9598;
        src10 <= 16'he5f3;
        src11 <= 16'h19a6;
        src12 <= 16'hd204;
        src13 <= 16'hb14c;
        src14 <= 16'h61b0;
        src15 <= 16'hdb7b;
        src16 <= 16'hb66c;
        src17 <= 16'h6e37;
        src18 <= 16'h2cd5;
        src19 <= 16'hf033;
        src20 <= 16'hbabb;
        src21 <= 16'hc62c;
        src22 <= 16'h7531;
        src23 <= 16'h3b26;
        src24 <= 16'h394c;
        src25 <= 16'hcb3a;
        src26 <= 16'h6cbf;
        src27 <= 16'hb7c2;
        src28 <= 16'h6da6;
        src29 <= 16'hdcd5;
        src30 <= 16'h3928;
        src31 <= 16'h2a98;
        src32 <= 16'hdeac;
        src33 <= 16'h3b1f;
        src34 <= 16'ha5bb;
        src35 <= 16'hf316;
        src36 <= 16'h829;
        src37 <= 16'h505;
        src38 <= 16'hd388;
        src39 <= 16'h5c16;
        src40 <= 16'h1e25;
        src41 <= 16'h1285;
        src42 <= 16'h4399;
        src43 <= 16'h949e;
        src44 <= 16'ha51a;
        src45 <= 16'h1a87;
        src46 <= 16'hba8c;
        src47 <= 16'h14fc;
        src48 <= 16'h2fc9;
        src49 <= 16'h3cc8;
        src50 <= 16'h4f66;
        src51 <= 16'hcef;
        src52 <= 16'h49c;
        src53 <= 16'hff6b;
        src54 <= 16'hf5c;
        src55 <= 16'he3eb;
        src56 <= 16'h8c3;
        src57 <= 16'hcd5a;
        src58 <= 16'ha85c;
        src59 <= 16'h26d3;
        src60 <= 16'hd9b6;
        src61 <= 16'h1a5b;
        src62 <= 16'h4e87;
        src63 <= 16'hba0b;
        src64 <= 16'hea1b;
        src65 <= 16'hdca7;
        src66 <= 16'hc84a;
        src67 <= 16'he713;
        src68 <= 16'h1181;
        src69 <= 16'h6e14;
        src70 <= 16'h27ea;
        src71 <= 16'h9f13;
        src72 <= 16'h567b;
        src73 <= 16'h8602;
        src74 <= 16'hf9cc;
        src75 <= 16'hb6a;
        src76 <= 16'h2308;
        src77 <= 16'hac4e;
        src78 <= 16'h99d1;
        src79 <= 16'h2d93;
        src80 <= 16'hb50f;
        src81 <= 16'h35a;
        src82 <= 16'hb636;
        src83 <= 16'h94f9;
        src84 <= 16'h9056;
        src85 <= 16'h1f72;
        src86 <= 16'h360f;
        src87 <= 16'he69f;
        src88 <= 16'hf641;
        src89 <= 16'h8ea1;
        src90 <= 16'h8d46;
        src91 <= 16'h747f;
        src92 <= 16'haa8d;
        src93 <= 16'hd7c6;
        src94 <= 16'h38e3;
        src95 <= 16'hd397;
        src96 <= 16'h7b4d;
        src97 <= 16'hf9c4;
        src98 <= 16'h4122;
        src99 <= 16'ha835;
        src100 <= 16'h4a0e;
        src101 <= 16'hd060;
        src102 <= 16'h4d45;
        src103 <= 16'h9b63;
        src104 <= 16'hc74d;
        src105 <= 16'h4534;
        src106 <= 16'hd5c4;
        src107 <= 16'hc308;
        src108 <= 16'hf289;
        src109 <= 16'h96a8;
        src110 <= 16'h3bcb;
        src111 <= 16'hf2b9;
        src112 <= 16'h6b50;
        src113 <= 16'hbc54;
        src114 <= 16'hc8d;
        src115 <= 16'h4379;
        src116 <= 16'hbe1;
        src117 <= 16'haf55;
        src118 <= 16'h97e3;
        src119 <= 16'h402b;
        src120 <= 16'h3ca5;
        src121 <= 16'hfb04;
        src122 <= 16'h3a6f;
        src123 <= 16'h3883;
        src124 <= 16'h28a4;
        src125 <= 16'hfae0;
        src126 <= 16'h489;
        src127 <= 16'h4bbf;
        src128 <= 16'h6905;
        src129 <= 16'h775b;
        src130 <= 16'h8761;
        src131 <= 16'h9d6c;
        src132 <= 16'hbd17;
        src133 <= 16'hea55;
        src134 <= 16'hefff;
        src135 <= 16'h6e3d;
        src136 <= 16'h54b4;
        src137 <= 16'h32b3;
        src138 <= 16'hf875;
        src139 <= 16'h46f;
        src140 <= 16'hb01a;
        src141 <= 16'h4ba;
        src142 <= 16'he3a3;
        src143 <= 16'hb5a;
        src144 <= 16'hcf81;
        src145 <= 16'h268a;
        src146 <= 16'h7399;
        src147 <= 16'h9ba4;
        src148 <= 16'he1f3;
        src149 <= 16'hb9ca;
        src150 <= 16'h2d6d;
        src151 <= 16'h9dee;
        src152 <= 16'hd4ab;
        src153 <= 16'habdb;
        src154 <= 16'ha282;
        src155 <= 16'h2c3e;
        src156 <= 16'hab9a;
        src157 <= 16'hd90b;
        src158 <= 16'h6dc3;
        src159 <= 16'h5610;
        src160 <= 16'h4d18;
        src161 <= 16'hf06f;
        exp <= 24'h50e36d;
        #1
        src0 <= 16'h8a56;
        src1 <= 16'he4e0;
        src2 <= 16'hfea4;
        src3 <= 16'ha8e6;
        src4 <= 16'h7891;
        src5 <= 16'h869a;
        src6 <= 16'he2bd;
        src7 <= 16'hc76d;
        src8 <= 16'h7fdc;
        src9 <= 16'h7514;
        src10 <= 16'hb63;
        src11 <= 16'hb843;
        src12 <= 16'hf60d;
        src13 <= 16'ha52e;
        src14 <= 16'h214f;
        src15 <= 16'hd897;
        src16 <= 16'h554e;
        src17 <= 16'h5596;
        src18 <= 16'hc1f6;
        src19 <= 16'h59bb;
        src20 <= 16'h3c17;
        src21 <= 16'h429c;
        src22 <= 16'h860a;
        src23 <= 16'hde86;
        src24 <= 16'h8883;
        src25 <= 16'hc763;
        src26 <= 16'h3388;
        src27 <= 16'h110;
        src28 <= 16'h41d8;
        src29 <= 16'h54b;
        src30 <= 16'h4cde;
        src31 <= 16'h5115;
        src32 <= 16'hb92b;
        src33 <= 16'h3590;
        src34 <= 16'h8bec;
        src35 <= 16'ha1ff;
        src36 <= 16'h2e03;
        src37 <= 16'h24ac;
        src38 <= 16'h53ae;
        src39 <= 16'h4224;
        src40 <= 16'h7214;
        src41 <= 16'h9d42;
        src42 <= 16'h39db;
        src43 <= 16'h685f;
        src44 <= 16'hb89b;
        src45 <= 16'heb5a;
        src46 <= 16'h149b;
        src47 <= 16'h91ff;
        src48 <= 16'hd7e9;
        src49 <= 16'hfd2c;
        src50 <= 16'hd773;
        src51 <= 16'h4f30;
        src52 <= 16'h6ab4;
        src53 <= 16'h2dbf;
        src54 <= 16'hb0b2;
        src55 <= 16'h164f;
        src56 <= 16'h2864;
        src57 <= 16'hbdb7;
        src58 <= 16'h339b;
        src59 <= 16'hc3d4;
        src60 <= 16'h1fc0;
        src61 <= 16'haaf3;
        src62 <= 16'h7e5f;
        src63 <= 16'h8e9f;
        src64 <= 16'h1e7;
        src65 <= 16'hb3b5;
        src66 <= 16'h8ece;
        src67 <= 16'hf641;
        src68 <= 16'h1736;
        src69 <= 16'h3df7;
        src70 <= 16'ha7f2;
        src71 <= 16'h4348;
        src72 <= 16'hc0b2;
        src73 <= 16'hdbbe;
        src74 <= 16'h6959;
        src75 <= 16'hb95b;
        src76 <= 16'hff01;
        src77 <= 16'hf3a;
        src78 <= 16'h437c;
        src79 <= 16'h775c;
        src80 <= 16'hcaa;
        src81 <= 16'hfae6;
        src82 <= 16'h5f72;
        src83 <= 16'h6f70;
        src84 <= 16'h159c;
        src85 <= 16'hbe14;
        src86 <= 16'hcb86;
        src87 <= 16'h6c69;
        src88 <= 16'h93a;
        src89 <= 16'h43a3;
        src90 <= 16'h96a4;
        src91 <= 16'h9584;
        src92 <= 16'hdbae;
        src93 <= 16'h78db;
        src94 <= 16'hf85;
        src95 <= 16'h97b4;
        src96 <= 16'h26b1;
        src97 <= 16'ha81f;
        src98 <= 16'hef23;
        src99 <= 16'hf653;
        src100 <= 16'hc242;
        src101 <= 16'h6038;
        src102 <= 16'h74;
        src103 <= 16'hfccc;
        src104 <= 16'h6c9e;
        src105 <= 16'h4992;
        src106 <= 16'h1b9c;
        src107 <= 16'haedb;
        src108 <= 16'hc516;
        src109 <= 16'hca3a;
        src110 <= 16'hba92;
        src111 <= 16'hd4b2;
        src112 <= 16'h465d;
        src113 <= 16'hccc0;
        src114 <= 16'hcd0;
        src115 <= 16'ha426;
        src116 <= 16'he42e;
        src117 <= 16'he78f;
        src118 <= 16'h9ee3;
        src119 <= 16'hae0;
        src120 <= 16'hb8b;
        src121 <= 16'h8d16;
        src122 <= 16'h447a;
        src123 <= 16'h508d;
        src124 <= 16'h1352;
        src125 <= 16'h99f5;
        src126 <= 16'haf60;
        src127 <= 16'h61c4;
        src128 <= 16'h6836;
        src129 <= 16'h29dd;
        src130 <= 16'h48f2;
        src131 <= 16'hdc1e;
        src132 <= 16'h5007;
        src133 <= 16'h2d86;
        src134 <= 16'h7dd9;
        src135 <= 16'h3d66;
        src136 <= 16'hf54f;
        src137 <= 16'h9ebc;
        src138 <= 16'h5b84;
        src139 <= 16'h569f;
        src140 <= 16'h1fa8;
        src141 <= 16'h8d25;
        src142 <= 16'hc575;
        src143 <= 16'hd0a9;
        src144 <= 16'hcdce;
        src145 <= 16'hb358;
        src146 <= 16'h42ab;
        src147 <= 16'hd78b;
        src148 <= 16'hd75b;
        src149 <= 16'h9fa4;
        src150 <= 16'h1a41;
        src151 <= 16'h45ac;
        src152 <= 16'hc7db;
        src153 <= 16'h72d7;
        src154 <= 16'he9f5;
        src155 <= 16'h24ca;
        src156 <= 16'hb221;
        src157 <= 16'h58b8;
        src158 <= 16'h2bf2;
        src159 <= 16'hfa7a;
        src160 <= 16'h73a9;
        src161 <= 16'h6a5c;
        exp <= 24'h5069f2;
        #1
        src0 <= 16'hb371;
        src1 <= 16'h8c59;
        src2 <= 16'hff68;
        src3 <= 16'h3a5e;
        src4 <= 16'h61;
        src5 <= 16'ha63d;
        src6 <= 16'h2649;
        src7 <= 16'h92f2;
        src8 <= 16'h11ea;
        src9 <= 16'h925;
        src10 <= 16'ha3ed;
        src11 <= 16'h46a3;
        src12 <= 16'haba2;
        src13 <= 16'h7404;
        src14 <= 16'h7513;
        src15 <= 16'h3f6c;
        src16 <= 16'hd942;
        src17 <= 16'h6e0;
        src18 <= 16'ha4cf;
        src19 <= 16'hc1a1;
        src20 <= 16'h1647;
        src21 <= 16'h9301;
        src22 <= 16'hd527;
        src23 <= 16'hfe48;
        src24 <= 16'h1a42;
        src25 <= 16'h10c6;
        src26 <= 16'haedc;
        src27 <= 16'hc69b;
        src28 <= 16'hbaf5;
        src29 <= 16'hd1c0;
        src30 <= 16'h1f9b;
        src31 <= 16'hd664;
        src32 <= 16'haf7b;
        src33 <= 16'heefe;
        src34 <= 16'h65d4;
        src35 <= 16'h5dd8;
        src36 <= 16'hdf3a;
        src37 <= 16'h99cc;
        src38 <= 16'h67fc;
        src39 <= 16'h64b9;
        src40 <= 16'hfcd;
        src41 <= 16'h4887;
        src42 <= 16'h9e2c;
        src43 <= 16'h72b7;
        src44 <= 16'hb407;
        src45 <= 16'h584c;
        src46 <= 16'h2a69;
        src47 <= 16'h46b2;
        src48 <= 16'h8c8e;
        src49 <= 16'h11a4;
        src50 <= 16'hcdb4;
        src51 <= 16'h4254;
        src52 <= 16'ha452;
        src53 <= 16'hb170;
        src54 <= 16'h7e26;
        src55 <= 16'hdb94;
        src56 <= 16'h3fb2;
        src57 <= 16'h38ce;
        src58 <= 16'heb9d;
        src59 <= 16'h2631;
        src60 <= 16'hbfa2;
        src61 <= 16'ha743;
        src62 <= 16'hf94a;
        src63 <= 16'hc747;
        src64 <= 16'h2531;
        src65 <= 16'h4737;
        src66 <= 16'h18db;
        src67 <= 16'hc713;
        src68 <= 16'h709;
        src69 <= 16'hdd08;
        src70 <= 16'h199d;
        src71 <= 16'hd846;
        src72 <= 16'h298;
        src73 <= 16'hf114;
        src74 <= 16'h57d7;
        src75 <= 16'hec27;
        src76 <= 16'hb4b;
        src77 <= 16'hb052;
        src78 <= 16'hf482;
        src79 <= 16'hf66a;
        src80 <= 16'h862;
        src81 <= 16'h6e60;
        src82 <= 16'h1e2c;
        src83 <= 16'h209b;
        src84 <= 16'hac7;
        src85 <= 16'h25f7;
        src86 <= 16'he2c;
        src87 <= 16'h5a7c;
        src88 <= 16'h6e52;
        src89 <= 16'hb992;
        src90 <= 16'h7cc6;
        src91 <= 16'h8779;
        src92 <= 16'hd25a;
        src93 <= 16'hcad5;
        src94 <= 16'h6490;
        src95 <= 16'heb04;
        src96 <= 16'he2cd;
        src97 <= 16'h9e1e;
        src98 <= 16'hcc06;
        src99 <= 16'he378;
        src100 <= 16'h74f2;
        src101 <= 16'hd21a;
        src102 <= 16'h9bac;
        src103 <= 16'hf9ee;
        src104 <= 16'h6074;
        src105 <= 16'h768a;
        src106 <= 16'hecd5;
        src107 <= 16'hf05a;
        src108 <= 16'h1317;
        src109 <= 16'ha43b;
        src110 <= 16'h6afd;
        src111 <= 16'hea47;
        src112 <= 16'hb480;
        src113 <= 16'h2b78;
        src114 <= 16'h3dda;
        src115 <= 16'h433d;
        src116 <= 16'h6734;
        src117 <= 16'h70f8;
        src118 <= 16'hd629;
        src119 <= 16'hd067;
        src120 <= 16'h54b2;
        src121 <= 16'hdbf4;
        src122 <= 16'hea4e;
        src123 <= 16'hdb18;
        src124 <= 16'hb7c;
        src125 <= 16'hc58a;
        src126 <= 16'h19f3;
        src127 <= 16'hfd9e;
        src128 <= 16'hde6e;
        src129 <= 16'h81e5;
        src130 <= 16'hd71d;
        src131 <= 16'h8867;
        src132 <= 16'hf959;
        src133 <= 16'h4ba9;
        src134 <= 16'h2ab1;
        src135 <= 16'h2045;
        src136 <= 16'h17fa;
        src137 <= 16'h1c6f;
        src138 <= 16'hd651;
        src139 <= 16'h2e8a;
        src140 <= 16'hf1af;
        src141 <= 16'h1f1f;
        src142 <= 16'h5d96;
        src143 <= 16'had7a;
        src144 <= 16'hecb6;
        src145 <= 16'h31c0;
        src146 <= 16'h3941;
        src147 <= 16'hb659;
        src148 <= 16'hcaba;
        src149 <= 16'hc97d;
        src150 <= 16'h6c48;
        src151 <= 16'h32ef;
        src152 <= 16'hc769;
        src153 <= 16'h156b;
        src154 <= 16'h54a5;
        src155 <= 16'h2c0b;
        src156 <= 16'haa2d;
        src157 <= 16'h40d2;
        src158 <= 16'hffdc;
        src159 <= 16'h97a6;
        src160 <= 16'h224c;
        src161 <= 16'hc540;
        exp <= 24'h52da3a;
        #1
        src0 <= 16'hbc62;
        src1 <= 16'h3a26;
        src2 <= 16'h3f21;
        src3 <= 16'hac93;
        src4 <= 16'h5e0e;
        src5 <= 16'hd2ac;
        src6 <= 16'h9048;
        src7 <= 16'ha419;
        src8 <= 16'h940b;
        src9 <= 16'hffa0;
        src10 <= 16'h2ffb;
        src11 <= 16'hff68;
        src12 <= 16'h9d9;
        src13 <= 16'h4e90;
        src14 <= 16'h7740;
        src15 <= 16'h30da;
        src16 <= 16'hd158;
        src17 <= 16'hf561;
        src18 <= 16'h6bf2;
        src19 <= 16'h2540;
        src20 <= 16'he4b7;
        src21 <= 16'h2933;
        src22 <= 16'h1bb1;
        src23 <= 16'hadba;
        src24 <= 16'h4518;
        src25 <= 16'h9cc2;
        src26 <= 16'h9c87;
        src27 <= 16'hceae;
        src28 <= 16'hab24;
        src29 <= 16'hfea;
        src30 <= 16'hb81c;
        src31 <= 16'h6f9d;
        src32 <= 16'hab95;
        src33 <= 16'h4b9;
        src34 <= 16'ha267;
        src35 <= 16'haf76;
        src36 <= 16'heab7;
        src37 <= 16'hca39;
        src38 <= 16'h6971;
        src39 <= 16'hda93;
        src40 <= 16'h6fe4;
        src41 <= 16'hc158;
        src42 <= 16'h7469;
        src43 <= 16'h79d0;
        src44 <= 16'hd72e;
        src45 <= 16'h59e3;
        src46 <= 16'h172e;
        src47 <= 16'h6b2b;
        src48 <= 16'h1dd;
        src49 <= 16'h2c60;
        src50 <= 16'hd76;
        src51 <= 16'h1681;
        src52 <= 16'h2202;
        src53 <= 16'h3b35;
        src54 <= 16'hc7b6;
        src55 <= 16'h9d50;
        src56 <= 16'hf5cc;
        src57 <= 16'h6732;
        src58 <= 16'he3fa;
        src59 <= 16'h190e;
        src60 <= 16'h1faa;
        src61 <= 16'hb76c;
        src62 <= 16'h6f52;
        src63 <= 16'he115;
        src64 <= 16'h97df;
        src65 <= 16'ha2b3;
        src66 <= 16'h64f5;
        src67 <= 16'ha2ea;
        src68 <= 16'h8648;
        src69 <= 16'h2548;
        src70 <= 16'hfab8;
        src71 <= 16'hd18d;
        src72 <= 16'h465c;
        src73 <= 16'hab7d;
        src74 <= 16'h4782;
        src75 <= 16'hc4b9;
        src76 <= 16'h870d;
        src77 <= 16'h1748;
        src78 <= 16'hde0a;
        src79 <= 16'h32fb;
        src80 <= 16'h3630;
        src81 <= 16'he9d5;
        src82 <= 16'hf7ec;
        src83 <= 16'h5cad;
        src84 <= 16'h9b4f;
        src85 <= 16'hd3c2;
        src86 <= 16'hd54;
        src87 <= 16'hc82f;
        src88 <= 16'h2546;
        src89 <= 16'h9d09;
        src90 <= 16'hb898;
        src91 <= 16'hc399;
        src92 <= 16'he34c;
        src93 <= 16'h9e81;
        src94 <= 16'he0bb;
        src95 <= 16'hc536;
        src96 <= 16'h6c45;
        src97 <= 16'h85f7;
        src98 <= 16'h8ce7;
        src99 <= 16'h232b;
        src100 <= 16'hf970;
        src101 <= 16'h4917;
        src102 <= 16'ha42c;
        src103 <= 16'hb60c;
        src104 <= 16'h913c;
        src105 <= 16'he538;
        src106 <= 16'hf3e8;
        src107 <= 16'hcce5;
        src108 <= 16'he1c3;
        src109 <= 16'h4151;
        src110 <= 16'hce93;
        src111 <= 16'h5c6e;
        src112 <= 16'h5cd9;
        src113 <= 16'h3f4d;
        src114 <= 16'he253;
        src115 <= 16'h75de;
        src116 <= 16'hab7a;
        src117 <= 16'h45d1;
        src118 <= 16'h6745;
        src119 <= 16'h9b5b;
        src120 <= 16'ha014;
        src121 <= 16'h713c;
        src122 <= 16'h7981;
        src123 <= 16'hd9a7;
        src124 <= 16'h827c;
        src125 <= 16'h3a93;
        src126 <= 16'h16c1;
        src127 <= 16'hf144;
        src128 <= 16'h9e72;
        src129 <= 16'h3e53;
        src130 <= 16'h22f1;
        src131 <= 16'h38d5;
        src132 <= 16'h6e58;
        src133 <= 16'h867b;
        src134 <= 16'h43b2;
        src135 <= 16'h516b;
        src136 <= 16'h413d;
        src137 <= 16'h7d88;
        src138 <= 16'hda56;
        src139 <= 16'hfe2d;
        src140 <= 16'h7854;
        src141 <= 16'hb13f;
        src142 <= 16'h4e04;
        src143 <= 16'h9e23;
        src144 <= 16'h84d8;
        src145 <= 16'hb18;
        src146 <= 16'hdc93;
        src147 <= 16'h5ab7;
        src148 <= 16'hdd5c;
        src149 <= 16'h81df;
        src150 <= 16'hb4c7;
        src151 <= 16'h36e3;
        src152 <= 16'hcf36;
        src153 <= 16'h16aa;
        src154 <= 16'h50b5;
        src155 <= 16'h7596;
        src156 <= 16'hb0d8;
        src157 <= 16'h4d45;
        src158 <= 16'h547d;
        src159 <= 16'h9749;
        src160 <= 16'h9999;
        src161 <= 16'h334d;
        exp <= 24'h540fd5;
        #1
        src0 <= 16'hb3da;
        src1 <= 16'hd95f;
        src2 <= 16'hb550;
        src3 <= 16'h33f7;
        src4 <= 16'h335f;
        src5 <= 16'ha041;
        src6 <= 16'h3ed7;
        src7 <= 16'h8b91;
        src8 <= 16'ha86d;
        src9 <= 16'h8a50;
        src10 <= 16'h7cd;
        src11 <= 16'h5aec;
        src12 <= 16'h7e30;
        src13 <= 16'h9599;
        src14 <= 16'h5b14;
        src15 <= 16'hb919;
        src16 <= 16'h784;
        src17 <= 16'h7d6c;
        src18 <= 16'ha15;
        src19 <= 16'h4867;
        src20 <= 16'h88c0;
        src21 <= 16'hcc2c;
        src22 <= 16'h466a;
        src23 <= 16'hc3a;
        src24 <= 16'h2664;
        src25 <= 16'hd794;
        src26 <= 16'h4462;
        src27 <= 16'hc150;
        src28 <= 16'h5899;
        src29 <= 16'h7927;
        src30 <= 16'h3d78;
        src31 <= 16'hba36;
        src32 <= 16'hef8;
        src33 <= 16'h64ae;
        src34 <= 16'h9d45;
        src35 <= 16'h75ab;
        src36 <= 16'hdd10;
        src37 <= 16'h60bf;
        src38 <= 16'h166a;
        src39 <= 16'hdec5;
        src40 <= 16'h7d99;
        src41 <= 16'h9681;
        src42 <= 16'h514;
        src43 <= 16'h9260;
        src44 <= 16'hf2a5;
        src45 <= 16'h63f2;
        src46 <= 16'h88ef;
        src47 <= 16'h55b4;
        src48 <= 16'hf2fe;
        src49 <= 16'h79ff;
        src50 <= 16'hfc9e;
        src51 <= 16'hdcba;
        src52 <= 16'ha651;
        src53 <= 16'h39d1;
        src54 <= 16'hd1f9;
        src55 <= 16'h1c3c;
        src56 <= 16'h4964;
        src57 <= 16'h6ca2;
        src58 <= 16'h8003;
        src59 <= 16'h3948;
        src60 <= 16'ha9f8;
        src61 <= 16'h1d46;
        src62 <= 16'he383;
        src63 <= 16'h6226;
        src64 <= 16'hba7a;
        src65 <= 16'hc6ef;
        src66 <= 16'h25a2;
        src67 <= 16'h6f99;
        src68 <= 16'h6807;
        src69 <= 16'h9de5;
        src70 <= 16'hb804;
        src71 <= 16'h4590;
        src72 <= 16'h8601;
        src73 <= 16'h3d80;
        src74 <= 16'h382c;
        src75 <= 16'h876f;
        src76 <= 16'h5185;
        src77 <= 16'hb639;
        src78 <= 16'hce81;
        src79 <= 16'ha18a;
        src80 <= 16'h80f9;
        src81 <= 16'hbb3f;
        src82 <= 16'h9b83;
        src83 <= 16'hd5f7;
        src84 <= 16'h8350;
        src85 <= 16'h9f85;
        src86 <= 16'hdf71;
        src87 <= 16'hd322;
        src88 <= 16'h49dd;
        src89 <= 16'h2bab;
        src90 <= 16'h2dee;
        src91 <= 16'h59b1;
        src92 <= 16'h8bf6;
        src93 <= 16'hb0b7;
        src94 <= 16'hf646;
        src95 <= 16'h2c52;
        src96 <= 16'hf888;
        src97 <= 16'h40ea;
        src98 <= 16'h9ada;
        src99 <= 16'hbadc;
        src100 <= 16'hd6c7;
        src101 <= 16'hf716;
        src102 <= 16'h31b;
        src103 <= 16'h895c;
        src104 <= 16'h4791;
        src105 <= 16'h8a41;
        src106 <= 16'ha49c;
        src107 <= 16'h313d;
        src108 <= 16'hec2d;
        src109 <= 16'hb8e0;
        src110 <= 16'h5dd5;
        src111 <= 16'hcdae;
        src112 <= 16'h4374;
        src113 <= 16'h77f1;
        src114 <= 16'h2035;
        src115 <= 16'h89da;
        src116 <= 16'h39d4;
        src117 <= 16'h84f9;
        src118 <= 16'h3c60;
        src119 <= 16'h8424;
        src120 <= 16'h37b5;
        src121 <= 16'h1765;
        src122 <= 16'h5f7a;
        src123 <= 16'h5c5;
        src124 <= 16'h66e4;
        src125 <= 16'h6401;
        src126 <= 16'h4e18;
        src127 <= 16'hd909;
        src128 <= 16'h6227;
        src129 <= 16'h62d4;
        src130 <= 16'hadc1;
        src131 <= 16'h447f;
        src132 <= 16'h66f5;
        src133 <= 16'hf589;
        src134 <= 16'he736;
        src135 <= 16'h4000;
        src136 <= 16'h34f;
        src137 <= 16'h7e53;
        src138 <= 16'h8ec1;
        src139 <= 16'hd187;
        src140 <= 16'h42cf;
        src141 <= 16'h1671;
        src142 <= 16'hdaac;
        src143 <= 16'hf2c5;
        src144 <= 16'h9efe;
        src145 <= 16'h1f8a;
        src146 <= 16'hf68;
        src147 <= 16'hbe84;
        src148 <= 16'h61af;
        src149 <= 16'h51af;
        src150 <= 16'hddf8;
        src151 <= 16'h1aee;
        src152 <= 16'hdb34;
        src153 <= 16'h79d0;
        src154 <= 16'h6560;
        src155 <= 16'h2f69;
        src156 <= 16'hce9;
        src157 <= 16'hd35e;
        src158 <= 16'hbee;
        src159 <= 16'h981d;
        src160 <= 16'h8e4;
        src161 <= 16'h8e10;
        exp <= 24'h4dac07;
        #1
        src0 <= 16'h3a8;
        src1 <= 16'h2f78;
        src2 <= 16'hf572;
        src3 <= 16'h9914;
        src4 <= 16'h3724;
        src5 <= 16'h3786;
        src6 <= 16'haf52;
        src7 <= 16'hac2d;
        src8 <= 16'he88d;
        src9 <= 16'h834;
        src10 <= 16'h2551;
        src11 <= 16'h9ee9;
        src12 <= 16'h540f;
        src13 <= 16'hc936;
        src14 <= 16'hafd1;
        src15 <= 16'h2b5e;
        src16 <= 16'h4596;
        src17 <= 16'h111;
        src18 <= 16'hd42;
        src19 <= 16'h12b4;
        src20 <= 16'h4dbc;
        src21 <= 16'h5724;
        src22 <= 16'h3908;
        src23 <= 16'h8639;
        src24 <= 16'ha6ba;
        src25 <= 16'ha43d;
        src26 <= 16'hb0aa;
        src27 <= 16'h1f7f;
        src28 <= 16'haba0;
        src29 <= 16'h7ed1;
        src30 <= 16'h6efa;
        src31 <= 16'h310a;
        src32 <= 16'h2eb3;
        src33 <= 16'h34d9;
        src34 <= 16'haa6d;
        src35 <= 16'hed9b;
        src36 <= 16'h3c97;
        src37 <= 16'h6485;
        src38 <= 16'h9e7;
        src39 <= 16'h645f;
        src40 <= 16'h2cc7;
        src41 <= 16'h8c8a;
        src42 <= 16'h2b36;
        src43 <= 16'h164c;
        src44 <= 16'h9693;
        src45 <= 16'h3695;
        src46 <= 16'haac0;
        src47 <= 16'haa4a;
        src48 <= 16'hbdf3;
        src49 <= 16'hc678;
        src50 <= 16'hf8cc;
        src51 <= 16'ha95f;
        src52 <= 16'h31c7;
        src53 <= 16'hf53e;
        src54 <= 16'h6cc5;
        src55 <= 16'h28ec;
        src56 <= 16'hb03a;
        src57 <= 16'h5fce;
        src58 <= 16'h9df2;
        src59 <= 16'h3c3e;
        src60 <= 16'h8fda;
        src61 <= 16'h4c88;
        src62 <= 16'h5558;
        src63 <= 16'ha693;
        src64 <= 16'h16a2;
        src65 <= 16'h75bb;
        src66 <= 16'hc9d0;
        src67 <= 16'h2e07;
        src68 <= 16'h30a2;
        src69 <= 16'ha4ec;
        src70 <= 16'hb8ae;
        src71 <= 16'h9fa;
        src72 <= 16'hd737;
        src73 <= 16'ha098;
        src74 <= 16'hc242;
        src75 <= 16'h5ef0;
        src76 <= 16'h2ba2;
        src77 <= 16'hac82;
        src78 <= 16'h2625;
        src79 <= 16'h9468;
        src80 <= 16'hd9cb;
        src81 <= 16'h8577;
        src82 <= 16'hb69e;
        src83 <= 16'h984b;
        src84 <= 16'h4539;
        src85 <= 16'hd1de;
        src86 <= 16'h175;
        src87 <= 16'hb17;
        src88 <= 16'h8796;
        src89 <= 16'h78f4;
        src90 <= 16'h38a;
        src91 <= 16'h1e8c;
        src92 <= 16'h4c67;
        src93 <= 16'h4610;
        src94 <= 16'h1fe;
        src95 <= 16'hcd1a;
        src96 <= 16'h3eab;
        src97 <= 16'h6655;
        src98 <= 16'h2265;
        src99 <= 16'hcefb;
        src100 <= 16'h8b9b;
        src101 <= 16'h2ec4;
        src102 <= 16'hb893;
        src103 <= 16'h6218;
        src104 <= 16'h5700;
        src105 <= 16'h3596;
        src106 <= 16'haa8f;
        src107 <= 16'h80f3;
        src108 <= 16'hcb3b;
        src109 <= 16'hbdb0;
        src110 <= 16'hd0b;
        src111 <= 16'h52a0;
        src112 <= 16'hb96b;
        src113 <= 16'hcb8a;
        src114 <= 16'h3b48;
        src115 <= 16'hc48b;
        src116 <= 16'h7b66;
        src117 <= 16'h6979;
        src118 <= 16'h9e3c;
        src119 <= 16'h6586;
        src120 <= 16'hcc4e;
        src121 <= 16'hcd19;
        src122 <= 16'h414d;
        src123 <= 16'h2464;
        src124 <= 16'h94ac;
        src125 <= 16'h52f;
        src126 <= 16'hb60f;
        src127 <= 16'he3ff;
        src128 <= 16'h6c2;
        src129 <= 16'hc05b;
        src130 <= 16'hcba5;
        src131 <= 16'h4093;
        src132 <= 16'hb01;
        src133 <= 16'hbd3e;
        src134 <= 16'h3d7f;
        src135 <= 16'hc75d;
        src136 <= 16'h1dd4;
        src137 <= 16'h96c9;
        src138 <= 16'hfef9;
        src139 <= 16'h5eba;
        src140 <= 16'h5df7;
        src141 <= 16'h5474;
        src142 <= 16'h1a9a;
        src143 <= 16'h7065;
        src144 <= 16'h9575;
        src145 <= 16'hc3f0;
        src146 <= 16'h4538;
        src147 <= 16'h7f43;
        src148 <= 16'h5181;
        src149 <= 16'haad;
        src150 <= 16'h95e;
        src151 <= 16'h3207;
        src152 <= 16'hfd1c;
        src153 <= 16'ha24;
        src154 <= 16'hdae0;
        src155 <= 16'h16ef;
        src156 <= 16'hde42;
        src157 <= 16'h42ab;
        src158 <= 16'h8090;
        src159 <= 16'he472;
        src160 <= 16'hb6c3;
        src161 <= 16'h84ed;
        exp <= 24'h486243;
        #1
        $finish;
    end
endmodule

