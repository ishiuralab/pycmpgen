module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfef404bca0a49509;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32bb159b0334c280;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h403fb06fa8dc4877;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b087a4997d51a70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcd4272cfd78cb08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86713a3bd0d289ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd42c5876aca9714;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ec5d911d1db4cb9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7c57954b808c7dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1b725a3a90221a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40b76b2fb2a2d2bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h777ef56707e524a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64ab2022cef83a4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe6962f4e24f543;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1cf0e66c5b8dc8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h792df8ac68df3e4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf2e14f85cb4ec76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73cde79cb475d4e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacef1870d5e21f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50d937dd25a9d6f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f46bf891d86a87b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa3ff6aa2e5ffa6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9509e97461d1343;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79ce2745162d3d31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h957cd3dc4ad99cbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4db509ba3682320;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c6c7f18adce21c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a87c349f400ecd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66a34f17f1dc7e2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5728c8ab679dfd89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12167eccc10a3dff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbf25b2d3688810c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ebb9ec846cf2148;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h127b3a256c43e60e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48c088874691bef7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h865c8a2b7a208a81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98458eefe0cc9958;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48d9f5da776e0cd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h900ef98d8b91a34a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5f64d78267f1f73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7ad5992171903d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66db2f98b7838ab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b7bf6c861faa78f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd55243c93141dc45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e6f5009a295d938;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h610bccaf659a2f3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c3f6aa28156c53d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5142e01aa9975426;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8c156603e9b8710;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h729447f0d7b13c85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb810322bc742192;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26a11c69a20ba61c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a25e28a62df5da4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2643060f560e513e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87bb255f822cfa7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha95e5732454d46df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7dc74a092f07a29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1abb31f210444ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7776cdebacee9bce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habb387c6b850f54e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54bfe1b584f13edc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9acbf3e07b37429d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb00676d39661c827;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98da84afcb785128;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63f46ae13690c927;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ed021b1227ca43a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26a5200ab751ac60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cc02473c7dbebc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e641c89e346567d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b21c9b91d4f1931;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5bc8bb42b9982c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h622747e61728ccb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0031f5c515e34e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1153a5ea78fd8abd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0415ddefd18b41b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42ff9ee9c42a9678;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h875a571649b70bcb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h786783f304558a33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47421096b9e8aad5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda17ea41054f5579;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h383bb18488e949ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd39a8a5ad884f7b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe6b5028f7ec27fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he40164b6f2a37f46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2173362dd3de04f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e0498475d05c74e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30daa16e143884e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11b016a60cdd7292;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffd71ebd0d8fd471;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1dc81cc7a4fd0e37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27a7154f2f444ce2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cc6d15ef0065f99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c2996566de4c6c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he788a4fcfe4af4af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ca786ba41820b9e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42e856f2c0e28244;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58b962388ad2eab9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he577f5d1b19d01a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6e198fc1bf6dd4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d704c6a1760f3df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2cbd9bc5d000e4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8d01508cead79b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2eb0177e81b60bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb92cb710f5c12d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56a7544ea8de52bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he18e1cffa926e0db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbff51060775024;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d371541cbc2b867;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3928e997881b3f31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4ac1286e955ea3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha94684dc2c55e03d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3b9fb83e6961f31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab518f34ee6acdbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d348946fa09ca0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d690d5878514a1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7de4eb08e7f49404;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcffc4fd8e195fced;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h812c2a86c82849a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca16f6e9e27dfc67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haec5d116b1467a5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h693d2de76812f063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5ce57c470f2e07f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75f38c5da5dc1c3e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h528ce4abe41a0dc3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3398e080567c7024;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5e24f2a9a69a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81468c0f6b1f55d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37009ff04f7e763b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc74fa10a848eabd0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadf02f36b8e4e913;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3297c966214841b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea601c60b90fb4b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9daf2f584e866782;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddc31cab7909907d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8315a07f6d099412;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h336b033675c01d34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b9a74537817e717;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h432030586fe3701;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc636406753322a15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bdee3969fdd1f1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c6e1abd6e7ecd34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e6c102be6ced2c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25e0b7739b05053a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he638e92a9a248806;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h406cc918b47ec3be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f88b7cfeeb77d26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d60e7cfb2155c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haacdfab51d01bf41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6de97d89b769c34d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h507a92c912faabf4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3adc2b95d48bcfe1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44fedfb60f047613;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab84c4b31d344f82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a7ab8de9f152e21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21c9198234ab01b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75cc2efe92de67c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0f2989649f3e30f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c3ea054104d52c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e3998efdd925ef9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c921fe6355b3133;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78c87a12346c2516;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81037d658346b525;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3322f5f784b8de53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a24e15e9cd4273c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a5e38b0afffb15a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ebb695ed1da6b59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae27dfa65ddf1cc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff449be1d0e973f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4707369d0d169c6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61b8a754c427f8ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h842363c2ba572387;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c40bb6a1111179;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h526bfe7750c1a009;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e0ac6781764529a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc065cb27c42f1d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15d6791be108015a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96855c655baa22a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h863a27aea15ac1ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5086ef4fba2bea49;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8e8aa1f0513e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc29c17b444657c9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4326f821c661c15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3e680bf09335318;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h495af1cf49150fc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h115ca97f6805b9be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb00b9f1865fd1412;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8183a4d56fd956a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2604eb3b1f1bf841;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98d763201f6aad14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde11018ad6309ae3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5120cb2700591678;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4acaba3b47639bad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8db86b6f1ba0d0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a0717865f8c70f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b6a0d1c7f41306f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33e7cbb2c095e3d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49b4509461811fb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecdccdb3fc42d464;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb463d2724939e5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b52ad5dd3a1011c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h128161e5bf3dabe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8511396f05044a53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25826561fe1a769;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h350e8e2b11e4bff5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca2f8a9abd667b50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf48ebe6fcecbd8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6025c2d74dd3c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92296f828f55d87f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51d58cfa48e731c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha77d6075820f2161;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc93a41357fc4d451;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3871cb4141c3c08f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6db88e21f152204;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd368ee09b82c5770;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a9d078afa3e25ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h832ab6f3874ec9d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53fe4ea8367b185f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46683c697f4a7eb9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha62ac5fe7bdc442;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57bd4e9705907d92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h348147e2eeedda5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafb1dc406b39613d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64fb7db24b5d554c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc21be76c84a689b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c0dbeab00b06697;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1709585bbfbcff62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecaec5aecc748f82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd482d9df7db2d404;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h769a4411c94b70fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0a9e37de05bf638;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h483645aa423e3d4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b0c69c66382c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34803b494e6b86d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he77f9b0504713376;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc95cb106e01b8e1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6eb8ab66f9f8aaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfce691f98fe7f6bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc9bfe9b720cc30b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6e445d368c3d3a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca82e17dd00bb2d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c01cf1c1704f171;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3e111d3f9308d0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a97a6ada485004b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcac98c65a38ca5a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b84a0660fcae18d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h524a4f2fceed63cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6116dad97f1c20b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbab374343aa60dd1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86deaa08e70c79ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55303393afb805c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc75f3d1e723087d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56acb386caf653c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93c69142e181ff13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ed72a8effa4a364;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f021d6355f4651;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd9471bcc1041988;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8e08965724fb9ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79b07dffa5d89c89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h373ba9fec8081dfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h794cb1f203618322;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5bac0e2e8e4b1f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73b086cd5c59073c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8964c1d155bca77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb463fec14e31d63d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfbd971b876e4c03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae480601bb73962b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51fbb8a8a30bad0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb7a802f2a2b5bea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd03d3f4393fae21f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49c7bf271dc0f24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf77354f779482fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c3770798223daf7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4967d17da2b5752;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dba174dc64456ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1af951f648f63c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb075c44b7105549e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81e24b432522de64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h243c770d9bfaf2f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12f6783324ebbeb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9d3b85df536124c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h116f15fdf9d4c1a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1af0e9218cdea56d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17bff694d329d93d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h433b2f621b06c46c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f119add02752e0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f7cbd4345042f40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he92d8f7bd09ede5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1413a2d79d29e13c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48befd6217092faf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h928259e8ffa31724;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2ebac6c5c4c66b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3db19f8261eafc4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd300ae9e6139d6bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h835dc10548a93bf0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2512a74558d4e601;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84e816c87bb9530f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc560593bf66b24d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f3deb9a73e8d87d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59a454fca93ec9d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h496440d6a0b133ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78960cca03426cae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19fe4e2c04989264;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h402466c0feae750e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f3e0e388da5812e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32a7e10e539e83db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9db9a864dd03d846;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba0e1aea6cd52a81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h613fd41360a27cbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2e4a998444bd232;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9c2f28f93f992f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd47a85a6a0d181b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf96a073b3f8b020d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6287e93ca7426a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87132e69d841cff2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf77b24ba402bc345;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d4094108e4fecc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6774eabbe4a0f5dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42b6e63fd219eaf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf15e1a078dc58ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1110fe16540dd838;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8b5215171a7b05e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74281c60cfaf76a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd97ce96accc66e97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc58386c6884fa085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49818d1bdf046875;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fc8d4d1173afcf8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fdc044cf2d69e20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cb4a421801fc631;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39034f276b44590d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h825931bca3481946;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he80be648c1eb016c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3fc2622e35d4ac0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h818591ae5b9edc51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3870c46985529c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43f0050028c10172;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a065a4ccd48a53b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee4418379980dc1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haea88241e132563;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7e41d1132f55a6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9acef4e4c4bd7fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca3d9a511138a71b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560a7ae2e9e673a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8af5474e857a0df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb500fd437658c99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41d7efc5ee995ad2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he589788f1cb734f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3400f4b5787f3883;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h878e631b3d7bf15d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bde28634df246d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha914145c03c5594c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48302f59a4c6e3a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcda304a6cdd36f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5293ccffbacd609d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3f94ef042b79875;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3516adf6bff95f50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8aff53639d2f2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44d6749a5ea2b20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h498e8f5a94fb3106;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcad1234c8aad4513;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h416b47b3b9f3c0e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5275101083df1c92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf915573f3f2df3bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha875b625ec3f902;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c0b9a659a764ec9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he223f43ebaa37ef6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4f078aecf4d8e56;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab91b0ed8a8cf11d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd93e30307b34367c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17ce3351832a1357;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f62a4a5a41c8fba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadd50275c4f45b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h160e8d9d40a6a9bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d4c4233141e4eba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72ad8039aead9a69;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2c824a4d63c821a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h235e8437f06add6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61725786acba2cec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b6b5f721765247b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2de95169eda14849;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc76a63e3e6e283b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38fb46a0acea68b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3780411651d68492;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98d983557efd9216;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4821c654da223162;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbaaf9dd277dc8f91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4ac95a2fb02706d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h923645dd72583fe3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1aae5ac70ed49ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadf2a324d0a0179a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe304dd78df047b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3ca209dc3b244ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haec3c92043b03b41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h884dfddab987be3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h578e27168aee56e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33872f4f8f0a7d0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he55e6a57c8fe8b51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf46268941039cf9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28696131bc3efe95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cb8c998fc8c43fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2a9d61768cb95ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee5f07e877284553;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4a6396f6183f7eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96452726785a4373;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa6f37e979e0b9d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc13d6c6470dae19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fa0425bd4d83740;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8652e57bba7e5cf8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19b8a86da4214563;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9282d7ef8853c67f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha764fd6dcb1766f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda494a6728708099;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha36d56be603bc8ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef468f4f3e17d285;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16ef97bee3b142e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e6b1fc867be2048;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h952fccb4242a0d1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab25b0628c31d48c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d56d8794e9170f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93d55c3a0a6f868f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4645bb16ef01f47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e5da95715b1b1ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd18470398ae827d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74a2a161dd6bc072;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b11efb7de0c4b1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6c7fcfe7db6baed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9be1d5323611414b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he652fb2d4d9bc127;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a29a21046aa6eb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88ce829ff6b13be6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcb43363dcf4bb53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81969cbf634c23f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he00b1e9552eb4512;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f9544e5e6b8c1b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h212360805ba7c120;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48f110f47a4e6f8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce1bd50306e9dd11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7cbaa0ca626276c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a0b9f0227d50f25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee0fcf08de260d5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20d05a372c64825a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfde461aab60469ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda9427ffb9cb55bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h159111097a5ffdfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h571eb99da38f0020;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c3648268b9a760c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h471f546e12762683;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cb6614bb0479252;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34855f660478767b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb03deec56c5d22cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a6823d2a413a44c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1dce169188d59a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61e3ff9f898a26ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffad146019df0be7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc983b68130b34104;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc602066c290a0fc1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6e229d4be5d138e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0720229de2eac73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85039d806021a8f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dddefbc0c3e59ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88a22cd01bdd3149;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h142d56303b1b95d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d5af9e811128840;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefb35e391ca6a87a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h378d9e94a97b3e14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he721d90d3b7877b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99fd3baaa295e31a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7463219945561e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h776cd8345ca7e918;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee587a3892142063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf23e0424c04e43da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd21ccd66d6606024;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd04990789ddf0cd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdff6f3405799625e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2981c553543963b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcef0bd3c86d67383;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f4f2d14fd3beb16;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0e4ccd125a055c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef5040f47478f087;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h478ead295850e794;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae2252afb756680;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfd267ff24822abb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb611cd12a826d88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5fa4460f371c723;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0e66ec55be9d000;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17e4ff605dca8103;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6871b96ffe2563a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5bf6190d52b5489;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ce99d7e6e6b01cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb7397cc91d8b2df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43a2e2f032f874d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb68bec8a7f86cf86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74a273144a251aa9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9b8bf8b1c4b1d68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbb6cd8768a58495;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0fcce091dbd3f7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5660758abf84f789;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3670510867878f88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72334ccb0286bff2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb64d2f4ecd34ee7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca0ce198cf1d7792;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10b843da36345781;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he09d6b91747ff9b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h291463e1061feac5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2aa9edd5e94f5892;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73ce7936c73ea385;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21f333844e4fda49;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb62eafc58dc694a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4da9d90a53ce4bfe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7feb9b524486e521;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3371db5e179a4ae8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c24c3568d410c9e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0d5868b4a96dfde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb52581367c444b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95d6fac6d88eaf1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h542ad8522e084d5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93d0170391f20836;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha49ec6c5c2e88d59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc5c50a8b6fd57fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62ba446eb8bd6c48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he84d8a1536036b5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40db21081e9e1ee3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h976b8a4d1ad670ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59586baab5144ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5479b959db4055dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4e824378914c816;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf32ed086793065a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46b944db0f57639c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h200d1bb252adf55e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38a247091f88d476;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb8f428b51ecbbce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10ad69dfc522599b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda8a88eb65552038;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he925eab2cfe8dc52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbde32315b23450d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41a390c6c6760d87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfba104ebdedc7a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h538cb429b57c5af7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bab7c5545f7b32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h882e346dae2ba8ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce4f9984bec7a964;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h800ebfa443794711;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6449564e5be0de02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58b557b51d4443d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5968f7df539c48c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3201ae0d30bc5cb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a03e8e487aced00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbf9ee8365f5837c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c8d044539e11db9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbaa0b607db903f3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c964908cc55744b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf89560140f2cd484;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6174fc57e2beecfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5a41b9e07530bb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56a0dc1bb4c5b71f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had83fa78b01d9284;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95cfcc15a6c73793;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h649767622f67a813;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc544b60094a1dd01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb3e3e65bd262c6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce5a9c0c67e7f352;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1acf935f6311a12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f0df1113332a840;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8785aaf334c321;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b8e434eb3860b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h829d1fb65565ae97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f8dc4eb0c48d5ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa642125915cf3f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb44fb1c590d844f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81e148531d205807;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4243f7377c6f3e73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h251dffa5e3542b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff9ebc80e191f64b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f56f34c2a163977;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc88252ba9811295;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4adeda28a39b9508;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ff2bf7f5c9c2659;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha95c25b6f9e1edc2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16f6dc0ed64f6ec8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73eb6e09e2d0b36d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57b37a38ba97d882;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he29e1255ff549ca6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3d230bcdf8bd4ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b6723318df1763d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf6b0ba0d0f19eb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h370c8b4cd98829b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5441671a4a366683;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc98547c7363098a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b9f7c5fb617949b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20a9259e976a8bc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8827e1054fe796e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a9a9f05db97f00e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9293c7e4870c04d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2df3a6a20f5d920a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdeac7f0be597b98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c2d227940d7fc83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56c4cd093c619dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105d31211b49455f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aace31f049f8898;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8cc0dfd71320711;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc795d8aaa75c2562;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f211ad7571a91e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a07ea31c9b53e89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebec5cbe5e16a829;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8014735c48bbff2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a83255f10173c89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea2f7a24cd891ff3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67ced6b63e16510e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7ce560b38421f9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3ccd0d54fc052bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbeab102737c5c9ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c1b1f98d16918a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h173eb654cd81490f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd814bc0d98a29cfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e0821c54a71bf94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32225b7e15aae820;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6309c1fa8cd0627;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f337184c5271bdb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8619b16d9921043;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6391f50e9ca055c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98276277614208b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h418c21afb4a0780b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb413c9df755dc26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h380a9b6848d17a72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5521d141639b1d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he35ec11d9dcfe3a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h873a6d183fb5c4a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b90511c9250c8cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbbdf6b6d4257cc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had3944ad57f4d199;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3257ab32f4c9c5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ce7a14599ca2fda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf51a14e2d1a02a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54716a0721e188d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had23b66644d7ef63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7745bd6c04f72a91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf83a21ff6b48dfe0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2edd1979c66eb553;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2f492f62e3fe4c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fbbf38b254c5299;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f73b8c94e735524;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4594062e59b69a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47510d114492d4b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94e4b21a8af55b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec086e3e83978278;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9aead6bf466678fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4146c39ada848986;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a948c2412ad9d66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd71531bdab71be1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafa862ec82346c70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92be3222980df6d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fba1bec0de4048;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a8218113c26fca3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2158e8251568f7ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb523aef8e2c6995;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29812ca7d6bc80f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5fbd2cf13565248;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h585c5d422d68fec5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a97c8bebb7215e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha60f9f158bb5829;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed33abf2bf12f1ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81d727012e18aed3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h251c4175e55db43c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59fc304858d59377;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48d6ae9bfb25497c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fe1e0d26b62de0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd29e6af4312a214;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd26200e15d14313a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd04784844a6d6a95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcffc56191922f9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97e19e6e74b03792;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h607257bbf4c8d51b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf78a3e840e926933;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe623f823b03c95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14c43bad34282421;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e0aa820ccedecde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5842c1ca5f7dbce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24f50e4261916adc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6f36965a0f687c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c02bbaabf2a2b8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h344ac7bc615c870e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h677b983e1817cc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba89db1e155bd0ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h158b1083265c79c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb28a331dfe3b17a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he70bee5375b86577;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h955ae2b9dbeb517d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf88ddc893c937a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54478e1ad49e6d4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf079105f30c00bb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7168a1175d597056;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbac18d9a50eeb40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h177e5214d5ae9a30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a77d1d30d85d0e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef273a0d6490de29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc9d0415ef5b83c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha417fec868003983;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefee267e92c52066;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8ff19a1e1c7df39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72230a1866c78b5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h212be36c5bb1fa95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2037d24704361e63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7a37cf3b2141a76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbf7a5a74f55b085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9067b922beee32cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceb1c5f2eece8e0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ee20bcd2cce1881;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9fccc06128baa5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2625a983fa9a126;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b91d9eea3e80dc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda8d52be21b8c59f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2fa2f316ec6e3f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88797f7865a90068;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9fbef74d64cb490;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h902268621bc439d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb561b3b98a227f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff47ec0cdf06212;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81f1614d68fd0de9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68590af489a5173a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fc3675a55d9c1c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha64f66dbef59a979;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97fe9dca86f307b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd957a803eaf228a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4e2e9f8629c3c95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e5a574ad63b88be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8d6dd4385f4438f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he42386721f37e718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd3d0d832886181e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ee853682f3e6ed8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6baf9ff6797302a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8b90c186d0682e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h199e3b6f7e27382d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ca3f6ae5dc54dbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4118a28a208ea1a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb80c0a2f996d7e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f20aad39b566225;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe5dd07a996bf1ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had2de29195de18ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7498ea49ca983c91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58243f4e7a873983;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d0ef6b94ce091a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5b40499a7cf8347;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfe8502cfad9ae2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he14b6a7a932e680c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb611e2e0611f57e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a7893ee840c1dae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa5e9b64089f45f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17cfde538716a49b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h704d92d75595b1f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb45188c6fdbcf4be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc12def49827607f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff60dffcb2e18816;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2aeefbc321428b82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1db865988b681822;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde35b9f242f27a33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57312b4c90602b72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4766648a5a3269c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7433cc52e0d8e9a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66b29436e5e8631f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h138e56a07d22adf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39b1cc47660a72b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfde55f38a1c684b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h280626206ff9d587;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f381d5040c76f5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67f04e2a598e7207;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9640672f7bea1da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43da165a296d9482;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h289253d3ae16840a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf476479a2b2d1f48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b0c0ba5ce509abb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf330dc53b335cedf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f700321a570b052;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce533e84c6453c0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbb4435d49d81f4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e280f36465bcaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc463f7b9d636ca6f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9f8fac382420a48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1496ecc1e5b8bc37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb46cac49199683ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha16160a0b94c21ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13608c0ccd85112c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h613d787688731593;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70e7c914c5fdb33e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha02310847aa9ed9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7897a987303fd718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20fe319aedb2cc0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h609f50527d5af696;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560bf3c4043921a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd68f9c0034577ae9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90421a76f3ae4b5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfecd87d74c4d46d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43f75ca7683d9d62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h121da55908a9df90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d22ff70a8e8820;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h141912313bfae0d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9240bdab6126a347;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5030d0bd3f15400d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha38327b2b069c555;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf7a18d96731a002;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fdaaccff4de052b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he202d5df3280186;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37148cce7041a0fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88a2e47c86dfb622;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6263827aae2267af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d15ad7d56dda45c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc738d5dd629fa516;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80e805c44de014de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddc852d999331968;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4774eb16f35fc1eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f14eac054c5c82e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fce6f8d8a59409e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h614d2f6e37a51d04;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1f16420c78df5d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2109d6923c2c5874;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9c356f3ea6cbb5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c0a132edd69404b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69451d3b9e12cc15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8c0b011ed8b40ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84e09e676d367ff9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61d2128ae0f1652c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd17160d3386b2e5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd27cf2e4f39417ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d86af5882fa0439;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d679d0ea1f9d67a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h994e118c2ae12886;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3c439beb41c3bc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h183a6bdb3f586863;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he26a339f0c7fd06f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacacd6a1f63cb4cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58524cedc0422762;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1e51237adc5376a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51f4fa2cb4bedf91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfadfa79e98733d9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4ff767979abe2c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f6deedab56ff77c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36104de245e2fdfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec5e1ce9fc7b5e68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49a81d568ac52a0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79d59aa9811442;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h256c0251ba7efa97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed570c16575d14b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7f5dc938cde1df6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c1da8d162d39b02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c76a9c8702bd82e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7742f7db42ff4b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff5d2c6ebd13ae61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h970adf63a093e4de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8f566b41575bd5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0ebbf9d78a4748f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he15099b303974a80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79d3306299733719;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ffe3fb0538739fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha40de7d3d689cd4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e6536cea90cb353;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85687fef17eb4fa9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefcdac522cfaa4d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40ee1d54e22062ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h747233f11f151274;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h112fb9076a0943b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2784fc0f1f5d6d19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe48c85c80bb2e03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb46f86f90e09b26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b7e9ef090d3a655;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd5da5c892638338;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfae80f2d679f972a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b6e803296c091f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb1a8529ddd54fc1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3fd32046e0e75b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c3d8a6f574a346e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15227d8b0daf06f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba62124e17fccaaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa2fd640f14201b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf7db95ee260ff98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h143f416017f3df7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha557db73b7393245;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7b3832a9ad4cbbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9123ab8f4da7b1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff96fc9b47bc4284;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cee8de547c7375c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b5940eeda2920aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h747a33d03726d287;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3f152ba296bc08b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45471d365c4741ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7447b47624be088;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf76dece3ea5504b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dd3e43bf7d6d62d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h248a05d710259960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79dc487b7b2060c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3527d6d8a51a7028;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h466ef95c54f9e2d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he49feee112de0693;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7a7b0efd96051ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed3cdc8d8685d3c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfad8276f8da96429;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8c266db7d848889;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62931179c05f7a68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e41310b3982d9fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bb74997b75d4fcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8dfacddd5aebaa2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88064a0a4a7dea8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d7bdc1f6cee1d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb337c2e5cfb50cd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66c5b7368e5237f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf15defce9f44122;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cd67b3742daa173;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he104ed3035a6dd2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h336f09a6a724bb44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dd0060831e52d23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f4a24259e3117cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2067b5fcba969e3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a37f77f929d4885;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a3ddb145cda7d63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc20ca30997519811;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11f0959e72c04930;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8642020e4516c27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc39a9c4db14b383b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b83fecb08911ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52424df6382509f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45e5148de4cd2e72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h430f4c4ec69da485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h366f9fd2d163956d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74f3d9bf558e19e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a5c48a4c3d5ab55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82fd9923f3a25dcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haced1007add1bd96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6197d8d03ab906aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha824450a68eae2cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80b4907cf05c3f35;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h634c72c4c0e5b4cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9df612675c50619;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94f260722557711b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc89e225f348f3ac9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24e412046eee6172;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2149d85a3442facc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c7865c3501298a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd61ac9c17c8f9167;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8677120f95cd4b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9afa71b1a3d9f20f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb562a99ffffb2866;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91cfed0f5b86e2c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d86553272c5dad5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5811231f81194f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e6d61c81c778a7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h893fa7f423695c3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29a531c40d94d6f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4eb3aedd0d8d9e7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e3ba16f8d750664;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h179e3422260a8271;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e513c13542c8833;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2240beba2fd4f98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7077dc752d5f33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c5407550673b264;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5714322a2a705da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e290f3929e3f00a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cb2da51013423d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6986c1287daba5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce3f2f12a483600b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72921c39b2b8b26e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5b19dd7ee490ec8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3da528d9b70636c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2d1d0ddd9757a9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff913099e86b7f20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf69dae8d0a34b77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79bd8d1c1ad06abc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4af42e2962eb39ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9d68f5a81a21d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4aa54bd1daecd22d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45c246135d4f8c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52aefc502c0d882e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d4d5132fe261c51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbe3a07bf10e5b2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e0a5bf355a93d6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59d17525aed1ef8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3ff87c38791f671;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h335351ab09a27c8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34bed9631dcc6c43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a43c6da6223e2b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1289676a46a28e06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3642f6091ddfffe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbb139caecc7b7ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5106790023a9fcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c5bceefca2eded4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8b6fd20ecba930b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2e0d4f68d5dc409;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc94741fb9b2da2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8175fd8b09e2e22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h213ac6a33b55f9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfa99e53b33fc90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab8b28753fc0e5a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h585c6556b99b25cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34812952094d5139;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ca41ced37f174d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c309b47a6e3d59c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h864684a617e85f2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84dae467bdfef935;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbed83b529e9bcb69;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6f2b39b3aa20ebb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd8d1eb354aacfa7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h719088b7010bb96c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3573c2e39a0f01fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h534c18fb88e99856;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d0da849439ad488;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1c0d50c1695a5e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4701a1ed0c7c8ecf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb603d4303a982ed3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d8c0c56564cd521;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92225354a2791da3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f7a9f6846f2db0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5d0797056bfa787;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32e7271997174b13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dbb1aa5909b86b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda8e98f76d6b476f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20e97725c687554f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h464e64faf5641674;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5014a4fcfecc8cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2623d6278b875d72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f98c0bdf7fa469;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hede4dbd7317d48da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h802062394aa3a469;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7c2b65ed407454a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf08238c413faac5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bdb3366745c49b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c9969d7f614aec4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba3dab01612d9465;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd142e99187fa1eb3;
        #1
        $finish();
    end
endmodule
