module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [15:0] src17;
    reg [14:0] src18;
    reg [13:0] src19;
    reg [12:0] src20;
    reg [11:0] src21;
    reg [10:0] src22;
    reg [9:0] src23;
    reg [8:0] src24;
    reg [7:0] src25;
    reg [6:0] src26;
    reg [5:0] src27;
    reg [4:0] src28;
    reg [3:0] src29;
    reg [2:0] src30;
    reg [1:0] src31;
    reg [0:0] src32;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3])<<29) + ((src30[0] + src30[1] + src30[2])<<30) + ((src31[0] + src31[1])<<31) + ((src32[0])<<32);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h964f03ca4d62360f50291a7f37f4ac5a6d4191b6a2609aa98ceeaa997600b4139583ccdf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1aad48b424ff21a4f4f8993bd92afbc7c471fbe7e735434931dca4c5f4619d6a6c00c0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d15d97233b0c08a1a5d38dcccdd00c049dead8057704ffa7ecc7cf0caeeae97ccd69f758;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cb814bfede31e9804bda0fdf8f2aa8e2ae8f047c0f8dd2dae797a19da7a0b08e14787e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4165f9e806ba7e5d6f60411e88a1b87ab5ff7f5c8006f1a4a81bc72bacd7f57b00df2e99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19263291d68ed2c2eab5a2fe725996696d35dfd66591cf6404d675639c098e0b8c29b021;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50f58a278ad87dc0c4cbd36e484d240b65e6e05b0684f4c4041050be3873f868c6e284a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee1d26180c3488d3d5c6545cf6cdc9199197ac013b076370abe6a401d4ba4ec3da6b2aef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26f417a37a6f10bcb8fdab377647a4b8d68783d3c85426c80a1bb6df821698dbae4d379c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190876b99d5130426baac7dbd5c8bff6705b8dd3c40022d53ee4994d1316f772a73d39eac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1844dbfcdc752f3ad3735bb6584d894d0fbaee2811296b9bf68d8b6b38a5475e6405dde89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124c35ade6ab86712d0e274023a42f5f7bbefe827a92548d0fd06f534073e6c90da94fb60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e3f78f151ee7cb56a55d0b12c3130a92d8e55db18e4dbeb36df08f7c579adec859e8d4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2826b513f47c58d7c8fab238e362f9a049045cd05a320786f0cc9db72df0f1bf1fa51fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104ee4617f392241d6314b39d94ea827e92d4d62e967e490c55e581dbe9e8c9535bf11bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65c3461942b129264507a43410e15d1ef337deac64736c09bea5cf0158a7ca491e45bfdf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1d7abed58c3296103a54f390ddaa219328900ded4ceaebacc6812d398d6786d60c999b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1e9882c7fd66abc2d780a0542954935a41ef213ea4fc094eb3dea9db03531130900c72c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7f72baae4c8fdd24fbf9c877b3ea9fae5d5de152f5d68a9f9ced812a34c61f59b9ae2fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135aa9e37514e1546bcdad8c318b1e80a0b1f4f761e893a1a84b9efa14660ee843c2fa2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9317502bd1d1e50eabcc2b2f941fa8d5e05fc240951efd909775e36341fc7ebfc65669ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbfefa926ee4633ce29e21384f621d3377d222337297902cfb2e98f46f89315aa690fa75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c74a0623ab44ce7c6de36aa3cd0c60ca7683f58e00aba001713c1bea6f7afb71e4a27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8265eaf2cbe9fd4f08ac4f55e33a4ff6f084080aa2a0b9f4dfdfb7d941d1df590f58ee6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131b3ab8015cc9e947e48d2ac99be8f1096a0afb055b6f5d92a3b6bad46d4afed1d969c56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144866c80c7b749a6f98880d9f86e35942db586359518a5dd585862680d5e095aea2a87d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1684de4494a2059b483b1e9cda309db3fc89912fcd69a2c1e5438a41677e086c8300b1d64;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf521052607d3912c57f8e3738857d71b6d24d321abc73fd4214c500f4c04aff4352570;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e525fa91d767b22fd5fcf8aa21ddf2a23efa4954457a8ce9bae30a02ae20de7c57bfef36;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1250eacf5cef53920f653bc7ee2545d9181736051e0d9a9ab0335a1553d12ad2130456b8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155245928e3f38b13096323b04acd5a17698465190e6e64d28bf1128cb1d96bb02b9dd062;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1470e68acda58db31f470256ae26922f1c9a4ef4eef693428e61ca9a2b1b184a81079a37e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef99916445b96cec8939d0674e0db0fb7f56d943d964a462efa3a78fdc30e882b7c9eaee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4defa0fb779412b77046dbe0d9090d217899a5a4c0c3e1d0a1a172a4f664e58f3fde707d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b42fb058c5ae870d8e4cac4fe79ab8db34528cbf967cd6cc44d7de60dc4542959078f78d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d4556a854f33523abdfd59b5716d3b1200f81fa788c902ffefbfbc2db8fd895fd62c9fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d68ad931d4da7ea3d6409e828d3b24a8c3caa433d7a0911bcd811972912ee940b7930fa1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98962a8523e36720d6be19795d2e3b11042388819ff4ddb3197ed7ea643aa7a445dc2c33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72b79109d8080bee94d4414f61fae70cad3c6a0224ff66ebf6417d31de555ac6e296553e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c1c86bbd933cabcbe7af055bd0ec8e73d4674974296e488afc18d390a93437c8fdf5960;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc185890c4ea07eb6e25e47ccb62898dadea10fc6c1921b15fc6c6495d71d33127d6dcc7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ddcff99ec9542361d5580306ee086ce4dd82dc807dad083543496c593a14468c6f64832;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132f09aabbb3d83a55dc160398cacbf3d2ba1c9f948e0151c24cd4602fdb99ea3a07dd90e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd594e33649394409bdd998497a328294da382b4c9f1a55748d3b7589457e72cfea340a5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d2f0628d6dff044d9c6c215833a8df2104735bfb89d42f24cfe5ca3ac18238ff3baed30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77a4057d6cbff760ce27cb7fa1fda8c3aa4c5c5338e14b1b45e5730a025185436e6422f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64d971445fed943ed86cb95f472045234a5557fe68e90d60a2763f04fd3ada382ffe8f53;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ad115e24da81ff6dbeecdeba98cee6fb72f1f1379d8ab8f76448cddb7d6dbad12104f46;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d1e761a53fe89d747ab208199390643a443a3f2591ec338e39074301cdd1572cbecfc93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfd1dc47effaa01c4b874e3b951e653af793bdcad0d995a63eb2d6f7a4e56d69cde38ff7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c198b8f05097486b6a835ee62d4e48735781322c037d2de29bcd0d4a9484926f81eaa9d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ef44f2443b95d35159eb6142c58a4e8271002cc7d37a3a02602b6dd8dfdd4afbf4fdd6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8ca614de670feb91066943ecf662a1c2bac890002c68bfc198636d77f4e6ae40dfcd62a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8a399ca04f858aaaa102b7e4631e5338238494fc8893c302a1c41621d64d90cd7e73b36;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haba92133aab72082a83e6ff558735b8ac5bd8a52d28062e99861f3a44109c1ea21a5b017;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a8d2b7c402bb69fa606efe242ecffbe8ce55a703ef7384608a1eae8e559499ecdc43946;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1accbaef83b478d2e8c6bebaebd0c83cca57c2072cca495266e2858fd6713a601f6df6a0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb464855a7ce7ec0aef794a72600c48a8a847a2afd17e90f6622ab3a6da113698f89e166e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120f0ca31e7afd1fcfd7ddde529988f95e51d476e98c674cdbc8d6f25fdf11b09b79624f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf1311e271513a8d772b811bda99a022d08a02065e75e244a1d72d320aedf758cfff38e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a6da044289e06bac3e6c047f240629105116e6141a11ecd149e8024df406e08665d0ead;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0c537dcd824791c26c9e7a1df59d14011964a41069e6422aa82375fc8d4ebc731711b94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa942d3c667bd619561c7a7770a31758d2eec9ef099741ee24eed02deaa7c64c694c4ecd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h993819128fe3ea67fe963f34318ed5a76a55be8569fe1574f695600885fc96160b18f303;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71f2cdc64c7200b477a1d57a1689c9f46fea41f10b4c33be91d0b79d01484171980658d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he18de1eb459623d59c71d7892c51c936b5b20bbf579f78b46556fe568c5d5941ae804432;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8fee2d6e94f4c40c18dc9727455a51758ffb08fa30e492c4b24b75a460b7d9d76c493de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb309bc35094dedc41bdd451ce966f9ef5de97b256995e0529d3dde67b976dbf85b030bf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc58eda394f773b5482416c8e545257f24ddf0a34c0ee5a00d467ee4d925039a6ec28672b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b57ef64e4d8303d73094cbbe7f05ff6a36d4e6b23f9c9ce5eadc0835aca4281cbfaa848;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe99eba9a6c7297941793c248466ab3932646b2fccd7dbe897421f73c261a14611e8f1f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe33c5daf702ad80073022f2caea851bd89ca9e5b880c5fa6d9adbff6ef53477d0bcd0b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9868dc34cee709f94b99249ba322bf015f1cbcf19d374af4646984a9931299f489aafea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h992610eff84905c081372a6a3b2c6579dd37ba9043a32b6ce13542771f5cdfe432ff59a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b13efa859f1fc43aa0c34983cf2700ea656124ebc3db68dcedfbb902a39db633354846c5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3a69621521e6bbf118daf89e405f7acbea23550aa7a127279c82efa4a96e9f133f59357;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1046fa541b1911fb45d0a30c50205b91f2bf26328128fa799a4a0e437c3e02cc83f1a4813;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbcc57f35a2bfbeb7edd66a38375b45079cfd841a5d404dc14da1e9e445b5e7d70bc442f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4552630822cb04262a081a5050519a1870f9b6ea113515f28f7e97fa8e116136140cd16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f82cb9fd4aee30eb568f3601ece5f5c346519347deeba17fa411111b00fad58aaaa9ef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2d96d3d4b5359e338bc4b5ff0f0f6f5fdde3f87d4af327e9f01d664479774ea23db6527;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65890d79cc6f4f9e78e7240251c3e9641d486e0c0f563b86e8392be0b401206562d5f5fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e2e3aa7d5e541d285affd1b8ca7f2759a5d9d97457330163aab61eb1c95e1ed2cd8517a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d099872c28fc805c9b2faf51a6033ad58956d82c65ef98e7e58386afd2d3f149d8bc207b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b0c12bd39199c38cbb97c6a490ed7f33eebaa5e2aec992bc43618269776787116d7027b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h785f12c1b53edc99bccbb60774f8e0904efc2985531138d4c5fbb37fbe8a95a66ff2a574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7e355670626942abe2838076434d1cac9f1379e380816467d56483d3bff8b3ad97b944f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5de9a1d76fc0ed4ab3ac65bc3115742cb7d39557ed5fb2f57dafd6e763dd43fa5685ef59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7ae2189be067eb8750977e1329c73966315741bc2d3c7a0aada9b8f69a48ec7457ae78b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d2485238d61d3d639e9338a09f5c2cb9d93acf4e75171f2a6de8e527a0b2e9545aa8fcc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b47e9edb4314864f6a123e75bab368a570150f1042e835645c2f2a55a1604c20c9557402;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bbcc8b088f68f0137f791ba3b3ed0f6fec7243647f8711579ffb8a14c97c763ceb27633;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7f3e65523c38994c6ad7c7f4a7b09386261cc3d35748b21cf3f3d659fcf6452312d9ee6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177d5f7cc23187920dd5dd0595509285243305e325e24227db8c6075b9da212ec06d26cbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed8a38e308e0183fefbcbe422ec01043652b4e15e432ccdeb83ba890bd33d3c04195972c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2d2a28446a2660f78ee3415c1c02602b0c5c2d6abbe68cb426998f222a6a7de369cb3ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cc6aaab9974e6e41c615c964be6650e4c18d13493caa6816e56b2ce0a281041b64aba43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc790f32ba4b758f7c2d5631e86a380dc51e8683fd6099318779262772f2f22eb290c79c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22ab5ffcc2a19cf6a63541e54cd816745993651c0af90361290060953a21c42abe5a0faa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6c8b0625d0d689107f30d35f6d19dc11aeb0c816b24aab7b73dc52f212519cd5ae0ec2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1340ca58d7c79bb2993999da202063222fb04ba0c313ee5949409805e7c4a9693ff2c5e4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea9247a3e1f5f880f086701d77339b175aa8b8f755d2fba0245588462a1703f90f002c3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33cefe5585f20a312dadc28a1230c2e65f7c6877335601787525c4d5626da7a07e37eebe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7d80a68c380fede8022e31b77735aeb31416bbb44206ca23ae1df1a1e0e25879654fe54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e32e4b7a4d14e9ccd4e4391732b4d1bd472c0b962e2c9c4b67c320951cc3d39fecf16d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a099d71076173a2140e14f75923bf9e1c59e0d1156cf5e91017726124d9c205890b19e70;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1325ea5819c128977006f2d8063e1495c0fb4c64d8cd71808aec096ffe0b45b4aac09d5a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd84ef9aa18eff01bcd9a9552fecdc30c37efb450233082ee47c5fada0d20d57cc843a64e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h533bf439b1fa620242bb22fadaaf283b554b549b4d5c0e7bcfc7dbf1df2f2d2f8a2e9c7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h401f20c9e7edccd98ffedd29a1c113e5ff1cdc4f4f42245b719d74fd461f377a3b7ebd17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c04a255fc47a83c685c1b7d9cdf53ff2e78ad3d567bac9ecd7ad419574882fba75df8ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1939905889a11df99b86bdb0fe58e300cd74896b314c0a766d7e7006f7d44cd4786290052;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1385abe721bd2cc119bc8de053b133d748cd49bded758c91763682d662dff499b09a712d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c7b4d4bc5c37005ce0a059c2090ec08eb586dbcda500d51ce5bb42aa39f6df4fe021e6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10739884d45b9d105325be8db022aa2e9fedc73f03c4ade7791006c4679feb03c725c3902;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef8452324d1099468d76ed3e534faf92518fb1d918f07defdaf694684b591b39485fb1b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144aba90214f8a349ad730b3e54dc0b415a66b8764315e585c1569b62485d29dec32eaf56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a76c3fd6337a23dd2047de24bdce2b8f41022bc165dd9913385c6b4becc00a1e0748659;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13894b0bd0dcad3ce43a7eed05437054f15a89bc83c94cfc2c392de52e8a04fef458d8b11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198898fbe3e1d59963d4a16d18cceb6b12052bdd2f73be086afc6da2b5fa043efae00a769;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da5094c707442430c26a0a668a373d3c9b1ad0fa555f2db6425e6e49586dfc1f6a84fdfe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d88a7cf013fd3feacfb7b0fdc0064c2935daaf21beab9d9a182adcbd9e6d608a41e438b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181f8df0441933ed7838ccc52ef24621a51d18a47b8677eaa84f95b0ee70362bf572aba35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1416fa86825f98ef5f3f38ed9c01daa4406842116d2e73e0968d45d899af3665ba14d6d26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc4aea538070ae7edfaea7463dcc963882ce3d163721a19b2f768e43555bd8a155d22c129;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d3d0357d5c4cff7aa13e94db0d28164483b4dbd308f4bf247b4964a1f22c6296ae4f229;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e24164cc093649d1ddb4cdec015d5e3c86a5b2bc84e290fd2e4603df66990a2c10d8495;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126e68eada593819fe850b9731174a931807d82314a728ba2fc6ec4d5d617a90f03d895ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191baf628572ab8a5cab8fb5d3e6ca2c0fe150c8e9370a2da0cad6d633e5758d223ea91dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c81bb8fc23f5abdf246752ce515bee1407a12799acd95be281ba3fbeafff0199a8381b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11da77e3c2bb6f7c0effe971f6e2d961d23ce01bad087ba77b63b8bc5cfad9d705a7b1002;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36d43234ee6369917b22729eb4ad39c253b1e7bb7bfd747b948698239245ab8565ade387;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d814c4758918301596dfc74354efa40bb85c29bb878e84d27313e5a67eec9a40868d8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e249601db66a8bfe2df0aa7c9effac8fd7582ec6877859bf419909d550017547c7b40d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c7de8f2ddf5d7495f63e92f9992f6cd68bd12f6bb4f9eba5998ea5435e9443d213d8b60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b48b8eefe37e6bae5ad0018d7ae328478b1832ff9050ccf16f2b9bbef5d5d6bda9d31b07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d0eb2ed3f98c82deb61d2c85fcf0f397f33846f38a859b529dbd1605d351c662fbf2706;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae38bb1a98b42d37f39071a7db327dd84839aa3e6bb951320b0cb51952e502255a136ee6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee540fa776a8ee26c2b4b49ce1ec827d7d2d95f066faa333acac2482aed1ba142e8a56e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b2ab73af8c932e0de92f184daaad8024962fd69df77af3c908092f9e8bdefec9e809725;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb204d707ab0c1254f6ba3f0fe67cf53eac50a38fe6e3963bd75cdea529d7646dc396d1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f169df847181b9e978403620ac6f4887572fdefb824f8d960a1bcc43ac6597edde0af9b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99f533486fef4b2c349e4d15d50a49da49b6ac023cd67bfad507480bbbc075fc17d1309c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11185727fd13951f0e8ef4ab0deedd4a70a5873ea6bcc01e9b76de38f7fed5b6c76a4fb97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171c7ebcc8d21b2b04ddb04ca09ceea45667139861d87e6df139c4c1d7de540307fa9b47a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1504ab03c63f0ed881fbb76ac3c7959f36d90884730092fc05daf4db6d30c0f895271ec77;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23de1b3fa123feb5db15cc8aa196cf36a678947a99598d6a4499854f953c023702115967;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5d32ad13e823f5599580749b3b9bb89f0e7246dc99c44d10acb6e39ed049837a377c324;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a641b7998cdb30d4464d555875312dfdee6676c7ea44262f1defc49522924e0aa5ffe87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131b1d9fe22d4f873d041926857cb7c6d65b1b5cb5cbc9d28d56a6165e3e995bb2bb624c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf0acc402c7090fab14c7e2b6c1bdce529f01fba5e631970d006220f9262a566e6d32044;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e54793748e3a9ba5e846550d6777b1c398b50da672db7fba40df2af6789a427333fac958;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a96ff5237addd4541a7edb8d29f908aa2a9a802d753aa90935041fce81d9581f5a86426;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136d1b980a745b32119a5147ff209deefad994cb2a7ff54c3c626175daad278f5e87c6fd5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h762ac24d3c51089ebe235c181f3b2dd43285cdcf44f2c6436f822fb25d9a6f724ff8cd92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ea50137f07a9e608c418d1df6a0aefb51491902cd580e3edb22440845828c0e88aafe55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c38d82f3cbf540570280489e8c321712a1ebd76ae067dc6723b6ded2f4ebd603b2a7b44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a34ab2826195cc1d4b65c763d88cf2540d43c8007d7d961c6176177e53ffe6c8ae0bda0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4c0a7839b5e71480781800983cab1bbced63d4ae3d08d3927c99e8ad13c7eff78cce919;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150d8e97ad65b53fe8e6def188a279242eddc67838bb2907b6b7f484d10b897698290b283;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16db824b2889ffbe9eb1784ad50b0dea7865bffa61d47ed2a41f4d79684d460c3aa69fa30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78580860581f0df0e5cab68cdf92b6f94dd1176a1c2d153c22d8d54ce40720099e209bc4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h696ee43ede37168e5d3850a6eda4b20c7dfff623f7ad0d19fc769a7e598f93e6ad54b5b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e70e228fd005c0d37fcf0c5e978f370ac7fb63d99ccd245383959b02f6c16c39b3d44f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55066c76c7908342b595e99ce0636fb56d5f491693934c3f4874bdd433839f12c1541ad5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70b6675e022a878f11b41dc2a8161333d02aa41d7c6b8dcbe7529bda63161b1d41db591b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf4a750095b13504d498f64a320b8402e0ba05908b256e8d23b44f8f1a5217541cd6d25f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77474f0e3d68248df8dfe3f3a795e241450de3906e7451e9e4497bd1e3f142539400303b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dde677104181a38ec50e79eb1b146a45f7c9a83030bcf745032b6fab127ba800cd712767;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1943b27537937806a2eccb95f817d015ad1f0c118b26445e2cbc2c1caad4aa3f4de9252c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9aa99ca5da794a52f0b59dfb660ae1e918e199782f2a628f1270492ca43828ff876c4bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d201ec11f2def73f3d2824404574de3798c80db11241008c6d7852cd699fad74f8c0aaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b60d90bcb18fc2bfec6a8bd03e47d246cde1a8e296e29095bff083136ff013bfac5323f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e95ee633d96cff81db97f51229ae2fdaefc7630b94b93002dc9ce8f28bc8b19c1c5db27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19032239f07de7e5f7718ec3bdf961aff67ec6e8a21b5906e3353bf468020a079dde5b7ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3aced6e777f1dc42395ca92852d2a44b6701981be413b60678ef4422d605c8b0ac33854;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cb506f7f6cc0a24e00084bfb8d8cb7f96674c79f53e71bd1aee8da7920fdffdded1f0f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc528e102fd5c1d124bc56d2991b1f972bd88e6b5ed0885db3be9cabe3ea6e0a443b6ac64;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1c05ecff0f91d4cc3e08f83ab413cc434711275e8dec72d01aa8f15c7e51c42988061ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ebd8d6b57a6ea2f6ea6a870859d060b06f81287981c38f59c1caeefabe19998a67f9728;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17466aebcac909b62673effd8ee4978ce66cbfea762b6094f44de87efbb24f07d90fd53f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc771e6f9988245aba66813d94ba4a631aed0b9a84ee108e89ba2e4aba2c0c0505228d38c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194d464d51ef41e733908867296872d82b59154a9875fd881716eb21e851ae24e9ad0520f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h332fa6bc7c27cb9322791e778c80c83f2d2908fb762941cbb8efa5193c737b88b0ace5ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cc796e6caa882e4709a402b43e1aa42fdb47bfe4dc8ceba99ea0fa38da215269d621799;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3fcad30d4f1b73f2f3075729cfb0349f7d09c49609cfc8faf122bcf0e5da169612f65cad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc89363db044f25818358839f718922a70ea56abce2344f8e3128021b8309c5d3c4f287c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a85bd6806fcb8b0eee45b50548a76a5d40596a3490b23379cf9e5ada00e89b657de131c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64bcf24b88f77878161ee7d9505350410abd166f089b748da1d6be9877c60b188b0e0c6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae5fdb6c1759b562e634fa2e3c86cf0b5b1e0b2704a3e94d9beb5763e60851d4e85c2c38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebc4a212898d42d5310c5d63a74c108a278d37132014f2937474164ea28f95195ec3729d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1388ccd582ff7a6e48c1172839f672b77c4f6484e1f959ffc274be7c2f31055536e83ef9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189f4539ef920cea84e487359a36733cff6fc0b2187440304efc37d8846689ef97f3f3679;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55d5fb6aba0ddc295557beb3303afc9a694fad8dae047cf17f20f3b85de857e2f6768dee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28343f5893af08698fd7ec7df807563194d454eab3e5b5409774addfc8e8ae1b16d873df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aba36bfe02f27f31f39317f83d28ab38a9a0a425822a2e84bb0edff81dc79fc18a4ede1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h833df2c115c846ec890f210291501589a52c78ec480ace4f4c1db50fe28e4ea04a0dbaf3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b8740ea013cce38332a1104af946b089e7460ac3642cf8ab33d1b8406fd52c54a105f78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a73098397ba0617adf45a9c4c9ed5c84f31eb03a9d9029f3c3799ab2d2b283d75f02a27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1250662ed778a365bcbc7383997221b53902dc3b483e13935b62b0bda551307d31c557345;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d589e8d2a97e5589c342d81bbefe8dbb2f6901fcdaf81408f685c2d7f8b20b117f3c074;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db450178adda4993dfd3f95653b2f2b7715dac4acc16f4a755b846abbf150746e0091786;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8765dd53eedc55b7f05412578919d3aa2b177e20f58e4199c8d84ea17b72c74a0538660e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32b6e28c64a291fe73962f24efea9276dccc97314a84e30da48448efcc2e3341432752e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0bab521ff142d74b4612619c9b2c733d7e99a68866de08043506022b19be4c8adc7b65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3d556e7e74b093f2fc3706141660367b15f1613cb11760119cc795a2f94f590d28438ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h736068c481311562f4dc60e5d8fa05fdd3df907cea433a3bec66c4c2c331939f3f5ac3af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd040d1d59a173cdd71134dd7610f7daf9eb677a6146136ccffe2358c762916ef030fd278;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5b50e1d0395e27fd4d13a4972887cd10c2f62a82a644412136824f442d79d98f608aa4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ae2d946a85d6dd4fc63f6b67a53739ecc1ed00e27dea1a373db4b867d083d2617c0559e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cfbd1fc08290b356edf348467c77a7245ad5007d273db8bcb438699b6a6b9c344e580d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d0bd749ae175bb3cff72f8480963f6a6c48065962016d6179053e42b7ba08b6570ef388;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49ecaa8d62c76dec0a7c3b45ae5d8dbfa3afd5e9ee04dc4ed9619d858b51c5b17106b7e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d85612b63c20be848952270cb2ac083f9ef18535d67c355425709032f97965e466c7ae2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f6b262a244dbdfecb54c93ed3fe7b5e1be9497e18dfcba10fbb3b98e9b55fc9b583fbb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d3fbc03baabdce758692439e2b44baa63e3e13730cdf48c1ac3e9e33175d920147c0f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda0a28385f5fd6ef007a99fb67e71d56dc8ff8da7e72b135b4785869cec62d4648e49712;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1159ee71ff402ca8ae92e85e39940d03905f889b2c53da0a92cbc9b74805325cfdc116c91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc36147383568d5fcd48fcacf5c8bf9213e5d69e86d19b79f4bf9d9446f2929214d1a1bd9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1149ac7541360adfd1f83676f3d0b12c23d3a981909af1a2e8ba4da12d85fe15682f85c52;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h619d2c5edda39438fb5fb7a502c71e02f1a4d234c29b2ce7ec58a0b506585e1c56652c4d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa925d54d43a914565916018fbbe633619f5c7b1d2ab4bafac62b788ef2566b91a2c4f0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76ba8a9f7a41ff149fa7c25602f2eb806753b8d6dd3869d025f61284bb0d603c3bc01677;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad9db39a14fe400cfe5ff309c2005a62a4b0924e2a3ffe6aa5506836a32e1d8c04dd83fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146a193fbade3092947ec3fd8320908e5e75713dba8ef9bd77349700869a6b756e4294c40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca8daf5cdc20b5a61f1b7754c03b36da5f0d559759e9da57a2a64b300afa04a6622c323;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h499ea25741158b0b321b3a6c70531016d0e311641001c1f1f33c7209a493702ab0862d79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5b734e8e4b3fbdf5183ae355cf0e7f40f0457eca52eadc6e75de6ff9d247e305168f53f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d162175c5721ed0242a08593c5b90118683e1c3a211a08391cfc54d3cf07a34ef8fab81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd1e819590a5ec040641d7662467f8a49d181315c0e7aa69b8e097674cdd86f8dd8c27cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfaff3b09953c39d24ea88183d2ead2922dc60d941790b8e4068ac9db5186824a949a810;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe3c4e7710e725c626458b3d0da1afd20ca03eae6b2b9cd5552b6f869c4680ce61fbbb9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1304bb2b82b11965e86de74abbb7d2c349ca2938232bad3f8e2b19e6706d7b15b174bc637;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h399409e1e2e421859531e887e190d6d4d0fd3cb2c7e50a969ec35d2152504ab8dcd6d7eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81471c38ac0dd26b64ebf6603066b282c02a0ab76cc0b789ab695ec76bfcc4223d5b590e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d431e1850ab50da79086ed2ceff4162e4ef1137b2ed876bd267bb4ba96b2b0a565608cf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1228cdcf77933edd21948519ed0d038d85fa9ad39686d8f79d5e37e6601f2c8da037c695e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e2a643b1782d9343cdb30ce569008a7a3a11fcc7ac9d2feb0059185b0b1baba1cbde300;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ccbbb3e7fe8f26d7d2ec6d7d2bd58e777e01556e104f1527f854d8a4d1ee4713efb08e9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5e108fc906374059a22ff74da510de05a36dc4cedad65c0c843e4b116da94239437a104;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa93a01f9b59c8d1d22528da308438a5b11cd34d4ccc48f269ea60bef387e12022af479b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104814a1ffafbd7b45ce39f850e0630f5f7bf038ca061957ef3130ce412600d5507df7a9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112e43f4bfb1bd37e35d7325bc0e4d060c7c9836f1e451a06a245fe0e38ead2e6149fd119;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b9af9985303c4ae0b07120082b915a4f18b1306345070117229ff8d7daf500191d13aae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1467bf85b3ea288855406c51ecc98820a7239b315c5e9129819425f5f574543bb0f9b0a2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff69189fd441e73cea5bd8d844f1085dfb76920d33a7cd2b8a15c1ca2503add8f4518272;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b9690e76922973e6b2524c39ed9fe60a83081efc46489ebd146e1d86f08ed9015f27efc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db53e4959aac26601457849cde891e9aeb22d797b1ae557d8b129940cdcb29cd5752b480;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182c3d9d55f30ac734df3bd02500e369d9482cef49f91ccf69be5aac7e9ea66bba79d2ba6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bafe2505d00471bd3e4efefb27f29c313d5ff55b5543c7c9282985c0db98d75e87672b2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1add0720b4bed348c2cbe72caa82a4b774f3a8724bd4e34613c3f98ac1b69c5ed19b0ebfd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa397f7f2082a95526ff6616e7c522842d016fe2c4764c22d9ce96cb40dbbfa3e9b3418c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c61458ace9488e185d593833054cc05570e4896596b603b0c25d2d70179bbf9fc3fde304;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9b226fab9478371581e0dff28bc6617b80d11e884a1f557dac3bb90c4caf3da598fb59b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfc9e0c889f7935df46f11070e1bffbefb99e9186e4e349ec3e0dcb9e403657ade70ec47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hada1a6bfd82c3bb39ddb2faa97ac071b0360366f5f3fd229bbeac9cb4e757eca4e69ca3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bedadda57170ccfc0e754f67a18dcc7afe0e09bc9054f2413ed7f06fecb2be8799fcf611;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbeb38e8b762cd840916030817e72b0ffd7708480aa461a0b91f3afef2144693717d6bfc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he908bde8875788b0b50406dd8ae43641b6a059473ae9ef378895b3c0c21af5b8e71000d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49cee65a7c4741acba9bf8ca738c53870677df257f9aec3dce7c2e0f8e31ba4a640a0080;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1653c99e2a1f9555e7ac1cacc529c85cf5befea6756ee7a9b8a17dffcb390021b9f15276a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2734ba5e604219582a76c1b313ee3c9c13db3bebb3cd41d800efaddfe6dba938b89d99b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1261982d574a426a72ba1723cf781d8bc899f69ca5a48c03f01dc1654a18ac2807138e15c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19dc06a0351a2c1c2a4e1cc081e9e120c70edca85b503baed13dfc928ddddbb5607cbe779;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ca5b1e5432e0db9c2d906525efa34d7277e8dfd770507965d7d5a1e69d1e50745ac1007;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6eafaf89bf4a6bd32905cffcad7f7e05cf62c9a80033cb51eb8e7ac892fe93cc6e1813b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1613c39e4e77f47e5933ae80e9fd92b690e455346f9c47f96c4fbfea7fc3c7144bc47186a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1804054d1d7e3596a40ba7645f547e4c04841a6883130bc5bf57b6e41ff6934fb80af69a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78f9cda47de5b9103b12464a89661a8e2f8dcdfd4867d43dd1a435e94b43ff8e66209dd2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1861d568b83a1cb2aa9c753bde86bf8fd2cfbe1d4292e1b4889015cb6fb0198873f31e8b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a8ff27ab0c31b442bb33311f2e60b307d2b00213ada256a1bab78d8477ddc896a6ceaa8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc763d82580287bd79f914b092b22b994763d328739b072ba4f2b938b64f40ec56916bb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e037b541ff5726366e49e690d38215bd7fc6208c67a4826a9191b5afe0a3f5fef2a1a0cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb27fc7d67258357dd84ad8eb032d3fa41763437ad661ef7a9e29af12919ca7d1bd2d096d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b0d91e825ba00ff136ae69bb9f7b70d72e875fc4639fcf6df4ccdbb209ce44ef97a9fe6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9c3641e8258ee4f1b97dc7d5c79e22f169ac4080e08dfcff3bdcc1fcfb1cfd9b8bf34cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91aa22c15c758e47fb4b959b078f25f4c227dc5e9bf7a1fcedf1b602d0cb1df900198ef2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e03fb9c59f85e78a6a54c2b08a4d0bdbed55880592fa45d2f5a7ca202cab1354c2a898;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf47d5ab736501b57c8f03aacfe2a7f22927ae70d4d95d3718ba8920ac5e086d949bca23f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c4ceb1c2a7e505a8f17b6f336bf1bfd5dbfef9077ca61c6af0c02ea30a06393db4e203d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdc20382d061b46abd104fed98550a421c15cec570dedc30487b13fae6281d761de9f401;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39a45b08b47b16c1f0ba0d5a91a1a5e677db001060a8f525f39fdabb625a9e4b8408c327;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b58aea6c9510d8975ccc33be57b75e538f7306a6a48f29c8a021b8c3df6b436950f103b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197f6ec279b0dc8e3332166b5140c9216ffb2848d0d31284560e64a66150576d30e6d6694;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc51cdbc474f6df7a9af2561a9841524eede64ce5104af0db309da620a1c0bd8ec85a27dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b0275038dd73bcc5507684f7a7dc18f0f2883536581be3937e75f49871e17a892a87342;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe6e2cfbed4433ce57e3cb6f1d39c545673806587ab66b0dbce11d2fffdb806f84c6f104;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1e722e76e07d643df5801e03386d1a61410ac29c8f1d189a7b85ed2d4210c246c0159dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cb49826abb96888ad76862322f311cf6797969d55abee3981632857bbb569279c33e5d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1259a48bdd87695f0a8ba4217e7a394481cca1d3a36883de2af09ab8766a9397a75d013c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75dbeb3625d99998607a9a7c1dc3baad5a5d4fd5b7337dcc083fb8cd8e6c1d21692aa13b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1caaeb376d795a602422223fe2d630ea4c96631c63d360c91d8f26b46db743fcfd93dec15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe4354a15f89f1d9ba420480f84fae80adb3d4ff80d43eaefda6bb8bad3916c1421aa829;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90c2527a9efdffc70665db9d52f38b83f3fdb5d9b988ea85f1f616d62d5736097ea6207f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1912a7dd98e0850b03265f1fd86d85589f0239b1ccdcf761aacf29bc948798eea3068e76f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc3e38808f53321f19b71f5316dbf86c7b7090e199931fe0c440a08dde2d6329ec6dc33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h245f3186c7f2b04e2ae522f7df8e02e37427106290389f876dec16d9c3ad9bf65fa543ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h743ed94a78fbb4047745afdbe30c95d1cb5be8f1b7a7fca22e367101f2134f3a10c011c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6312842892699d87c676b411093fc06b23598b8ec26112a7992ce6029b6830da9823de57;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae5b26d6f2d9626728b6c8295cde7d919a9b343597fa226e2eca9727460cc2fa71d4d14c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b4a0ea77a32be9f61c56557c9413176d0f3907156407dd0569f9ab41bf69f48e5156c76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f091a80337605782dd751dc299081e33b4f2a91b9f9357817623881897bb93adadfbfc6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e2424e6a2c9dc7cdab4c1e3b700cf807505a99b6f92b988554fda8c4adebb0f43946a23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df2681c4c3b11632a7063ee16da804862c5a1a5e7c7bff574e0300ff9e8a14d40ec5ac04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98f700bdd117ad383894af0a437ca46084d4fcbbff57a5bb7e63c70f60bc809564accef1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h558859f36f7aaa9d78d0d35e55c102ac7617710737059b9d94b88a995ffd573451f080fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5249ff5ca6c7ca1ba652a8122a47778442210d2c3cb3d91dd8e79af45e3d255be89dd14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97a63b886c2025ca3597e40b52c3f6e30c6c97deb31655a7830ca8216a65fc791c947998;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab4b20a26cb4a3a3f68386c55d6d662748947ec654bfeb0d25c716b68c26a28942d6f7be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hffe3fe2635c675d7bd6fef2e404697b8bb225b1fd006c18ef01b3ba9c1e85e54eb18734c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6ee8c6013d45d2c630dbc802f966efb8cdf601dedee3b8a6f928f3e844208b22ceb9931;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b56f868fd1385123115aae61498547f6396f40590a5b7008d800e0e707fa7686665d0b72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf4efeb05b95b19e8e75122978b35e43e28bf4a2bf8c4c87ea94a924178cd06a40ff7458;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha38524db4aea3e16bcc3013dd60253ec304064b458e4d30bc2718e0e327d9bcb99781c2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1477f63670d20fce7c14d960b279310c0d04e844b0082aab25b7d5c6e6ee69ab3068b2b02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1845817d1a7f1cffe836e7febcce66831e6a2b38a5ec11b3938ceab14a9a84e7cbcfd3bf1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93d6545691179f2fea3b7fb2198a0f2dd691c8487c65d2d4b150cf52b6dd7f5ceeb05c07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f511b0976445f560a9a4cc208273f2961fe7dc4d9ff5ea5c977d96ea26ed5b1582b89f42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55424a42f39699be655b61c7404426611f1a8374d8012477a31d7e9ff55aba0d0a083206;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18541790a00b274841128cbf67f2ecb8969ba0b3ddca1432f71fc23a99e1b18d6e8adaeb7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f2f8eb1c4974b1e1bad08f3feaf46dec5300d1ca2542b7618c7aaa38bb67501e5a9006d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdd353d3b0e9a855a720c18f56560f33194da9ebc60af2876dfe27f1b838ab474dfe1dd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d438f6fd39936e21dba21ed9d451f08958879029b85c44aabc71061426d06c9b2c4f5864;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13651c32754d67eb9e614f0004805384c23007c68f9c2fc631a51bfb821d92ac71ad03c70;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e33cd1d11cac89543d05de0508ee4cec3c11f359b5747e87072eb4d008253f15a04db74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eca1e0a2534ac007143ae604fa674ffcce550bbcade394f0f7e46a49aee2b481fb9cee2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1222cd69dc80384d6af7b8b1e8d6a0855501907728a2943c4bff94b200d136e7da5aa332a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd384b59bbf4a38a48216dd4b893f3135563628ffe61c0a4dd7c7cfc5f73bfb79eb2590e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77dbba000a9e467d2911e68ea039ac351c58925fe5e4e9c98047aff61de480c33ea09593;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b7f68094e30c7b3d15fab586c67f9a71895eb7a4b14796b21e58b550c6f2d9b16ed4334;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aeaf8c11e410cb0ad4d62f966612664d02335ecca05d82b2ce464cc9941cb7e481be60a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa0b92f27448316ee3a80b18eb92852780815a118ad1f293a0d06db00db2cf9be00c7128;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11238351624fa419a65a764e020508afb65e52a8afdf8d3dea16c8f597afa59cee22cb795;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144d2ad2462e2852f9220964ed738aab91fb92aebc5ca99557f00ad5da61dc5e91336dfb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc80c18cd28779a1956673d5b12fdba5dc74d347ffd92a8328f7d12ff063d26de1070585;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h383dd89f32e8df56564b5d25b6b67a3e179dd488b102db090481865223690e726a88cb25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7ad447bfcefddf532b2987af104b2cbf78f8554f58c48d414cbe201e920c52a383ed978;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c43e442fcc4df9d0cebc6e62b785c8524bd98edac89b627071519f57855343041162fab2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f676d1c55570a0a88d6b45de2fa84aab9cf65a3a5907593caf6b695cb81bb439f668ff8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0ec9b60f2246f02a65680d718cfedeae2e314ad760acdbb1e646bc8cbfe5ed86ea91d15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aec0d705572a57d11aca5cd2763d90c65a3c5f0fa1daac276d4f3a0c4226577e8f5ed699;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78439a7901390c7ddf138b8f20695a28251e7219e3c6b4f3a83359a9b2c619a56dd6e8ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1562183116a0d734192524a91c64e5617e4e542d3a59f1125b0e157291714d6dd2d02b375;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9675be8f2a4cb0a1a4796d9b055c32a3cfc74707d4c35f1db18d58dc1f3d2a04463d719c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1847e6975e11d1c935801d3173efdf3d36f5861b749a695f708a25c5c405a5f57049d2bbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122a3a0f3175b32620994439b0a54c94d869513ee12ec9f7c4279122e9600e02aea61b2f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9bae00fed34e0a404fec32926dacc8f2a638597c001c0ba1b20085993ee78a591ae8d5c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbecfb9359b01f96ad80a0021319ed3d9a3c7eac287d1a831bbec81b94e2ed74e6875342f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a076b80e8d93a07c84a87bd663eb1cd1f248bbf65bd8f9da5a9b1776bbce142bc1922e03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59ab0eeca121a021e43fbe3b4602231cd80356c98f306e60256a110e485afe9044df23b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1effcf7e5244e18e945f0ee8e53e8f0ee977ee4b10780e7122a8f39fbf22b6f2bf50a2638;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163dded08b59ad2fceb2f4ff0694e61f75235bbf07c941a6612f9907336db97510077f6ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88ed46e1efe36f3f7c3a19625b3edda6fa2112b4160fa453feec86acbae8fe673f68282c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he244cb5c80e50bb65c1102014297e478909a857efae96d1dc1b72f5fb21d17d63bebea3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fad1ae66cd5f4e52be11b1a46e2fa2122c291f64cd01e9f46a9c7677386d095d0b14558;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha339c3164867795e0548b22f332c6ab0bd58e96e94a36c50fe238b1d73721a955a414efe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec4e230381bfd578c586646b29936465c80c82fb4d62524fa55c5490282ecbf57c21711a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb28703d228105969b2753d140a5a0dbc99170e09d1bd479039355a506f961b9e3c9ed3c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d1cf19bd1e9f7ba884142d710572aaaf0f69a57474abd01e3bebb79b7226076d003f0cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0da77e9ce7a65331b3990be08061021ed49d638b54ab38afe9089ba2ffba8bc0b25c3c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8a1b52a8780c6f7af7d05a98056a92f8314ae217c13a1be31254d32fb1a64f7a3a91cae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed6e29cacaac7bf388bf0b54c951d3404f5c5ac646b0e5d057fbe66f74e3f67fb6833f87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea51d15c00d31f0d7b5b5297ce9c26ec4dde2e6f1be02bf3d02c8fb17b9efe098428111a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b37251ca7fa39eaa7e99b2664ce8d2201d45340b0ffd2efee699e931e1d64a0587a3c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f774fdb69ae3b4c3e5c78a902b2c086d226bc253c468b9fc7ea800d5469e2e8f7e80580;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed689975cee07ac2dbc5f905269eb978596dd18e35be097bdaaf701ecb8d43736e088f39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18744eadb2395cf866e198b73d6d5812983e706bf32b9f29b06419c4088dab753a1c89f1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182d99198e7eeea8f38082741491f8d1838716c8390de22efae21ba81866deedbf6d43502;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba8f1bfca7a3fa1a0ef3f434afa033975d8f9ee1fbe87b053fb9de3abf98494d72b28413;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bf2d5a2ad4462713ed64478887c8270484bdfd06cfac86617c0813963545145937aac86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f67b1519e32337e8fc707ff9458b07a08c63efde2f472c00d28236e37def99e2c5ea9fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fbd5ba9e6b2d08713b8d9511c48d5a537ab729ca17b5f5936c76322c3337e4a1085ae6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db03e309b0f295af42a5c5a5b1a16757e4d24d69cf86bfc30827c1cb24750be5615259c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2679f8625d721b47790fd86425b2e1c0068eee4146443d690927f80ecc4322a08c74c658;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb5fdce51f7d44c100ed863d847492f7578fa88dd52e545437c9ed35fc51b01211f442ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h700dff4728ee42b1893a359f320e4a7ad414e3e4292f21cca15f9254c53c8a6ebeffe249;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3b65412b5a9388c7837119175c609f875156900a16dbf3b8ccebc74faad7f34b1c6c768;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140dd63d3791e5a72095391aff3c2e36d5c7668ff8c00bd2588a79412e8513dd680d7ee4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1867cbbdf67c3d2355c19f793ca9ffab1c081092ef76e7db5deb798edd52c76e1b258978a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79892df2115e80e7d103bce03b19a16651911c8d7ea56701effe574047276491821af8a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1210977a75aa202e8fd877c85bd5844151fab6600c29ebfe2bd7f7f1b6ed87b86fa3655;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47d5338c714ea1aad6abd09d1f19e1927ae946b352ec9060625e43d14a2b836a5cb05075;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168804c0a758753f24be0a161a543dddf6f809f1ec7cb7128803d9b74a01551df09f0c283;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd61b141a18eff646f562ba027215c895357d170e4eb0cd7b0309a54e58de04ebcba6ea3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e30104cb7cd06a1528a27a158505bc80ab4b39050deb5bf9f5d59345e45447aed8ef588a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b50d0047479d8c596b97b8484d895fa16e7cd388f83bec7bf0edaffc3599fbb6d0ad6bbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95673ac1dcd6b8202e63a2eea116e24047fc9987f82312f4ecef11f72e799e36cd87c6b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc91ba91caf01d6bb975bea1ffce954781cbd87b539c01c40c11f069c9ddb57fee1bdcb3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1230c456d80fe14eea72350567e520b830248fdd662da37dc59aa852d2f05f2fb87e7b457;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a17e3a7f9b4380c42a3f03f73058222a8fc105b7a5df94e5a56d1bc4700826e19deaf38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7815a0827c6403a0e4b99937150315dd55cfd6552386ce9583489f3b3db53d0198571e9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec86909fcca0998589f61a4076e631a99ca77c9d6f446cc0acbeb54e9813408839339655;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d67d7cb2a2cb6178c72f1e906c3189c55c2561e9f61eb69e2b7b44522ecc09fa1a84bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e39fc6d776e588759c59f2e0f149923863568c6d71e0b4574f3cecd1d0fe7745c5835f76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95300788829d6d48d0e3e03ccca2ce5e99e53cbe80258219efcf0ca6ce901f0da8bc509a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h205eec82f562d73445b00d9c8bb79967d37f6e252eeffed2bcf750a4271b0983e2d57e78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117bc00260521f6b53245ef2765220d1df3c5aa441f9ab0dc061df3aa9cee9c1bab222bc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dabf56e87ed2691a089a845ef4a4382c7bae0fe88ef26149d8807f711b99cb75efc9302b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177feb9a8519245f6d44559a36aa278d01c900e1680af669c2ea55eb4877cbb8a4a68f89d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15641a3e7dcfa3e443eb17c03b500a9f88ee3af8c98295ef599a7e648770673bfd46857e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd433f93bf3d6c1b83283e7e6e86fd15111e3594f04b9a1b79b33cd8dff9bc97872d3ce67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67ee3b878d4bbd6fc31b7f40e699c781e0848a33aa13b6ff96c597dd4012859dda5ea497;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6b16ab78b1bc892dc153b2f6478a49be327d6582efd71f62b7e29924da846f70bfc0824;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c83812276d90a7358c92678166fb8bf9565f26fee565725da68fc62f14b99d39d05038e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3484a3f2cad7a5c2e60539febd09b50ac665b5a4a1e53e623336157317f119dbf0a44925;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43ddcc49ba2cf7eeee87020ffafe59e2083d4c7aeaed01647c2771685ab6f7bddef358a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f43864bf8f26488210afdfcbbd38772499364d987923f42af452329c3117c4d43e71c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125d21d0c8d5c7cde9247e970baf4655efde95eb059d6d59a805d3541622abf329ee4b046;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1474d6d95269114826d86f7326717e0da892a23a713f99c1b43524c60f027ab532c06a115;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5c616dbfce0c1e1fd70002a9b775570f73e57bb1e30ca08e52923b7e8690e000cea7a99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bdd95ae12f74b2fc054509ce8e63c07fefeb6f2806cee513b677598906331d57be78c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf6652b7cb9f3ac52653d17a7dace40ebf5a9d1c58a5bfaede59c6f62ccb3500c76527c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15de4e27fb0443bfee802c0599c4c1ae6838e2a67a2681c1ad3c73de5f848ce6534ae7d38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd03cc5e652d8131588415a127c2a712456036a82c2e5c6f970996ba6b0af1093fdd130e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0f12cef13b52221a0dd10cee5a8b520d1c4f722e4bb00c81c397dbc2bfba55f1e8b099d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bea587692c1b360199fcb948fd741d28924935cf44629f8b3f95a448c31a5a995c4919e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a3503c1c1dfdb5a4e4bf8c299253cfdca5ec1ee954e3f63e012a07890dfe31c79a4751c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f354d2bdd8da1b9ba284d67e0075881e264fd05aead48d876eee9d5a8b08ecd4622fa7bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1819f3ee92959584762cfecac2201cd1974d4fa9ee8a3c2901dac89ac530b897d497f52cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c5e07c826704217b403993520cb3f6b613f7784895937fd899fa4b4bd30c2887077c122;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db90ab8260bea41e08bcbe6d0e06f96fe221baad938734f388319075e2ab0a591c782aeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5662c0f903b6599333599bf769866a8a2f0765d0ebb4bf625f115d7a62f656ce0e204a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb05dc524b9a036a333c86f2134e660e691da42f457371a6c3bb6e6f0c0d5bce93b0b3f6d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec19ccfc0c7049d7657c7d7596f875cf9552a9cb8624a7f7368958b23d566656e5cf0ec9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f6f1af34d75db1f72dfef7b7712d45f84dc5884ead11187c3ada1001ebbca5cb3faf042;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dcc8fdef9384a7b83b746bd013d53c11747d6584fb5dd95dc5a9cc146c96a46d9a0a7e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7c5bfc3aec157de3435b4659d4ef4313b0df4ae03722325b0892988c6b0b8e6b682b016;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18de27547dc16ae16e6883e8099cb9cd9a80a8dee85374ec9460dfa8175b6a3f1aa0cef85;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e928cdbff6aa64c15ebfd7af9efc7afe59df112e9b2f01354f6b385eab77ad171524249;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h679a7d8cb096afe773fbfbed1223566a4eeace2e105a15c497addd8256fa8d09a1d73a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e55d3403ed379d10ae8b7026e87fef60deb98cf9493c9d37dcf874365f56829a87d5677;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6df0683abefd767ad5e0e51828c3579adee19d8fe5552155737d9dd77c5d03bc55df21d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ce137540686c3af937f39d1bf419a44ac227181880a9cd26fe5322357b85a89f578434b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d72cc239f63cca0a54554b2efe74bfe2b0756fdacb2376ffa9e5b2e25ded09c8cd758a54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1819adb25dd6229e28bfb91fb4de3156a80ffb423ea7b6265e4df8a3a5ba5aef3da0826e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cf25133462d7dad2c0e75ec2ed710b27a0e174292014eb1a57389c62b800715fecc2f99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ec5d5a306da2bf7a65a584784dbfa15c523f10d0b2ba896019608c5ca378d787bb2265a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166616f19e45d28eca04a04da66b5466812099232dbc9e8198565b320c9027b23ba504e1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b2750a924a2a6c67d772aa6a1bc53a0a0ca25307f9ff86ab5e8c1a4add1bfefac81983d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aaf059252aaf7478949ebd69610340376941a0887094946f01be8950207db82d870b051a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f4ae876e8933de800135a8645550a88ebd77a480258954a4729543e21dc4d1e552b6d49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1815e3f875e1a35f58f290ccea5c492c40d76021eea1d44c2aafb4a36353be1b520473e1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef0b0306e721355b293cf27ef20369eceb953c5eb7d050b732bd1916526f1f9b1e2ea270;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f50c576ac353acf3cc622a1255e7a49eee34438eb0f5cc8a6a0b26431b3abce999b121;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54635eb4e41ba5dedd86825787c10e1e82612f72f4e718193ef20a4a89cba8261c24a1c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda9a36edc7e668b255ca3a978efcf581a1fce38831ba4ddb86735a4809352d9ba40c304a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfacd1b70b69c6ebbc00b241ce1995bb9177ea15557189bd9798371b82c74dee1cd0f1c97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7aabccca9fcd2d641c5bf9ea9d39b282421332d244b2a4893e5b92c7b4dadc42c454690;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50920b8b7e3922c4a3f107bae8c3e4486eaafcd9a0db1e23428fed6eddc7e5bfb375f904;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1120a2e495eee8e0b998221eea73bd4e28c52dda7775d19a6a40f7e8e2c3808edfcf0dcff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he89d39dd12e30f3d837d154fe1c4bb1ce141b878849667807f354f6e3d5edba837e894f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160e259a014a50f9e70a27ac1c11fe617c9cbe8a0815b2aa8888d97de4f4cee634638b139;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1182329e3ee06bedeb34614446abbbdb5a35d2e0b2af579d1573fee86e44fa128347b0736;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d75bb37b6e2d2426286276615fedcbc15504baa92872c6e0d89d76e0bdabfc998187d2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e047c58a1f3cba31bfbadb8d72eaccdd7399c9a64cd67a19b2231df47b6ad42d993ed9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7dcf2347902e6a302baf4218aea53923c58028696e40b341f6644e3d5d11ce6e4ed5933f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ef8e324d63d24ed0a240b7f632128b6e657e5673cd96b6907575d2f1b13f4b2bcb1a82d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d50077e17424c039c461e5740b72f5edcced78a9d3fa7765e1d354259bf27062344260f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c25906579f916589a6c73b310eaba29954ceb011c4a25fe0c86e47c7db52973ae62a2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7072d5fc5c06239dd11ac0437380dd5828bf216ae598b4a28516b344708d0cecf182a235;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10551dab3f70cbad50174773a08f0436f92773db872683045ee81ebfc5b33c7d6b2e2b138;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16525b750efe90ab6b21f8c54b12709a15e40413f1fda1a6e57e12d266f436bce39d074ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1635025d7c2197644f8180c434ed58acb72009469b33fe4592e23e88096efa37f9a01250;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d10a1f637b3d65314ad7e8432ae77ca080dc6ac2d557ef5272adc75bc61a7e899f574544;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a10f5a72c2c6f0a88625a204f4a416c54b8e4d689b04b16d9212516d47823b3c038496;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e76cd8453019e729ab2960cd1e7342a1edf713ddf7bc42772002cf4c3b9cf4c934d76be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd958c884734bfa8a2de65ff2bcbd7a34f662e143647688d94ae0c8e2e114ba1a8cc910ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1465207f9fa5b6ec532794612fb2b19dcead1f741308b62f2a52058004d7df1bbabfbd444;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d76c0e5a45a3c6d9e7a2b041970a7f440e443b01b47d92876063bc00ce7004f42bf034c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h46633270d79c6769be5943ad1b4c2ec47cad8dd0e9335a37f7f88da88357096858ef7387;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f9d4b303525973738252ffdcab341caba9cfdd66b80ce695dadb22577712cb75416d9f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178c5e4c01165abc86a3a3e4868fc26a38745493c5112f00546ebf4ef3a3e150a0bf87f13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2ead7b8d95e9765f7ae565dbeaf343744662bc5df4c123cf3b443b409f3ebd9d2c0c045;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1828a9c1bfef9d2b2ab2adfba3b4fcf9f67945409f252a18d76c8c4215260dff098f6ad88;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1045c19bb55b6f3442b8973d2801fa7b1a6e10eb291606acd59200a6f26e2ee2f0b368f0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155eac412537a152c378149a72902f5b3466a417d1bee8ae6b7fa72ec8658bd9304195db5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2c9ad285a513ba44ab430f6544776016d699d3c04e2d0465f5b247bcf01b4420823c7ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d566ae1a9226f590b4f22be75d9d5a247f5aeabc2db94125ceeda61342a6721781a2737;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b76dbd72847e6711bc9f327181fef3fcc84c17db88e7fd474afbda4544a855b5e044bd3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1838009cbf5ae800863ff35705c69bfe6c8173940e270dd9b3f3a6fc7815f9e1ebd1e58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e98f433916070bf57aa28b309d2b8d1b1b51c59bc892e7b89880148b98a166078a41ed75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h92e693a9600a1fbcb70590704c526180d5551ef41e989b22cc666be12635b18ce46428c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ecb24f2eb1732ec4d8de5c1ce9405b27b4570437358044c65cfe4e78cd75ce7ac3dab3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1349eabeef7778c3843c4d9240ee328c3093fbc3f3dc1ffddf9178d7aa3f87f6e153b7a71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1707dbc3be849a91723849e3e13a9f740963b25b1ab08e32f1a8bc6ed40b1ccdd7e25d218;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e016f0c74d79f4c17eaeb97613a968565367e2f72cf7d72fefb10f7023bfa9d00747041f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d8c4798464f7d00dcb007f85d2cadee09d9bd9966b0eaca689bdaeb9135ff1ba24c048f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h592577d2a2ab7ca9977759de9ea8a44a5d34f38d26b4e83663744606821e6b3d70bdbd78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f5fb724c133c8b758cfd0f1e2fac9030d0ddff5fa3964892e75ddc0ac43f65d8453b238;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a940a53a7739c6a75cff682839a410bf059030b523a88006cf1d36caf5a1ea936d3c30e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10dddbd61280ca10e1f21e2574acc3c913baa7db4b8ea76c5cecb47fd37b79c16560cccf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faf7f65a69184f6acba6f83ec449b2693f9c71a35fc71666fc8e965b61d6da9127aaef5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1106ea2077979e670174a51ddee77a8c34bb1b639b8f315acb69e827253970aea1c4232f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1128e4d4366cb594be53826547b6370535cc4c8a198ddb93f5d039855bec1ffb103c90f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b985f1aae3fcf46e8f5ef4ff94a5b95fb0cfc19e529860ba7e29aeffe5a2cd42ba9d20f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fa07e318b57b543ea6e72c0d11e9b0124b2e33c46fe2bd6c48755ec6c83767fc47690f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42ccc6685ad5ae2c4a9f85090431929b432c3fae773fd21e6559502fd7ba7631a4190cae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h128ed01a2c892137a33072d826e6e9a5a1ce37b22dd5a2791b66593c5c5cb56ecda8eef89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194b4fc982556f1c4e3b24e54f029f1cbcd664a29164dc41d3a93619dba40fc64ebef1de7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1052299dbe3c2836faf4179836fe8257808df09cc229ee2ffb9fb0ae7875451cb418d617d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha95d925e42989a61031179cea13eb8448c7b20f514ad68239c91e583a887af5cac3d9311;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179cb230c9ea674345d1196331192e6d86c4baf6431fb2b0760b509c8a09f0c5beda50186;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b10b63a6f230a881487e8b24cf1afbd0cb61f21aa0e45cb1249b187cfd93a914a25f63c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h552a64bc309e1a2d9be03481957d5e735c8af3e80dc6f8eb0df06bcb78576f3b36fdd06e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f4bfae81cfbbcbb7a2c7d3b1cb2eadc021b453a12a8e2d6bbcebd813332b6c558668da8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1526d79748cd5e838f88f19cc3993a42e1f18cd2c98244585a454c47aac19a40c5d3784d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cc017311afb7607d6f49355deb7269530e17f06c0b416eec568ccf737a5f072c25ae07e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189e1a586a40f065447a20be66a04e59fe5eb9fa74bd4723cedb30593a82344156f180369;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66901d328eb8848ff1d44c62618e68d0a24b329c5a7292f3b8c791f7665d96008730464;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc68a3029959ba947259b9c0d8b7eeea09cbd67f56203484da9c5907c353bb38afff97d35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc52c66c6806456a04d3fc1945b70fb6d74c324ab0ecc5ca02a5cf44c870838ef3e6d5248;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc2c8a4d99e5889a065404a7432ee7bc08538dfa3ad2501e9e89fe20f5662883cc162799;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c9daf52f19af3f0029634cc2ceb27d1bf2820c9e32a070fc10f4f40cbe2072c66cdd1e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4a1fb47b406ff976bdd4b4f698e042efb6aa1169f567e9e546527edaf9e77b3521bfa81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed1346b67b04131e85c177b44d63cf8969d727c91a41837b0eb6b9987649d51ae40f62b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18464f10228c4ac2e76585ee3739309700968a8bdf0e114d6d07f0cdcf940dea484107080;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116b172bd82fb3b71a896a1d35dd51528e710237cdeb1b2ff107e159f9d3f75d6550d1f23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9ec0ba53245ca7ee3e9a5cb0b4b71e864d20fd0afb12c014b9990d882805d525ca4cf7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd458b629cfb874047bbb2cf0bfbfb013f08c2e7eefccf79db15688512f16423032bd685;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1177596e1ed15d21fc13d22e1a3552202737f444af49a573cdfc1de977702dec55c60b29e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd0aab345ccaccd65dc80743f956cef89fe9c6b9adb2ad0993c8bf9906b2b37a26e05b66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc842385b26167136adf1219b603ec8152e1550eb8e056cebdb1b33ac504368b2d03efad1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd30935cebd85202bac1f0e163e19803fc7ebcc1fc72ad1fda53a6ac854d24051c1e75a15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf0d4f9e209b0d3084184f9ac598236064de898f4ec7de663f7ff113e2a5b512dfdf7760;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78d07c75d9a86e12e424812b061f403ec27eb12861916edbd16a95185291a99ea69b04c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189bb11f0f360c91d61d22d0f8686f77d09d2155b5017aa00ea71db00e9dc9ebd1b1cdd10;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182fd9b459ccfad465545fed96251c53aaee4f98967fb7516682fae575c190004949fa382;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bdd955642c41c6c33f04a3564d54e9dc9550515f5c8a8e9146628f42424056c95b7f79c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha19e5136593b87928147a7301b426dd6be180210aadc535f1654ee63d1e44dc831f32627;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197dc30e72e20db1b2b99474528bf3d4299b42dedd206966a91c94176dd2228264c995fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e898d08a457c8f325752c68051371a11ea3b6fb3e2e137c61f5c8a903ff453487903bb7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4399fd9188846f3a49f0a2d4542bc4b5e5ed78dd6e18c8cef1d28c0b64d0934bf62a0b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfaf2b800cddae3b315021fba2037b4cf823b52b24c57f249d2d8ab1c111a7bd2db94cc3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57edbe73a36c024abffae88ebaa684621f2e8be8324e5bf3ac47bb89cd3e6c77b3f08fc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85410e8c23242c03993ab0872752e2b648987f77803084c291928c1ef3b745cca2517e1e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dfbc3879805d5a6a6334d4e9a5aaafa10d4e1046be8a106e97db218b4036e31194dd9b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a30ebe3478142739621125232174d40a8852bc87a880bc37b9d7cbcd90b0e0655b9ee229;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59e38d1a26cab7d5eddb4265a6e2c35e808a9a8b2265c58dc009577597bdb6065c0c8c80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c2435667ac51e392d8db0a49a447198a4f4e465764be26fc91fc54d3ac405798d2aa3c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af691a6fef165cb94ca4abb48d0fd0c452056f479775b7ab28cc295b6360119998272f7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65bb4e0258d53eaaa37afd15bb0ca75dec33f3839f2b1d7d8e7539f2ccc6518e00864c27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bc9814f95750d3cb6d6da6b2df387211a7689bc5ea28da8c7871e3f71e21f9bbd45008f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94cb4070ade871f3be86da43dda1df0c61d2db84e0ac86204abd3fb753e027d73edb8d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118117da47e119d29d639377eb71f4b51ae50ea73e907db2b9f8966cbf308e3e9b076895;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1669f2b71f6aba9fbefe642222a01f61e908e7dd9c0fa02375852be186f27165d60d666dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83c204d6c0f886aa4c4c99d73a3840db4b7ac7dd2fec837fabf6cc072b5ce9d521df0a4d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9cd936d35bb8479968918b66e92536c5a16486b3a1ea2278d69cec0cc1b22db8bc1afc7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109d9cb70cd6c53c665c0f0f2730e9c0419f4765b99680c8af87f27adc3f8cfca38045dcc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193094bac698b14c25754232b44c0a221530ec1cc8e077774afc88336662884916e1f2017;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1530b107c95927c0e900580ef185513900806c642b73f76f71a07d313265f1ec607adf4e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b6212084869ebfee5e8ae9c66895992398ae42010ea6de1d012276d0145c21f60af1b82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf35c034c81b632c78342b1648ce2b9d85bae4e73448299da7db5dcce8f2ff8fd4c143953;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1445f609196f30dbe8c70683978b0f2185da4eb0134e007590b1723d7d6df84554106e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36d98c520c228cd34fb6b16be99e0dd974eb7741eebf5dc73acf8dc060544cc2a39d9ba0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe9099e6fe11bbc6d4827198724ffd61faec498479c33246dbdd19288d59ffe848eb0f6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fa1d4dcb34a0c7855d3f5a6e082b4f74ee7fefeccf8bc66a756f85fd0f77aca86af9afb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115af7a858b5f23600238a290ef4f702c338648bb4f1a1824d28aed9fe616bcc1bcc50e13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe4f10104ca56ec38e20ca29c403951c584e1dc6f3ab5f4ed948432c5457d7954aa9400d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5fd654da8c54ad53c015517043da1569617cf2dbd98f9eeb5f1b41af2b0b607f6e35836;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1078c2d4cfc2f88bcdad5ecf9a2a2de0a36b00e0c4207098974051b292db45f97da7f9555;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba8063f1d6a438b530b92527395c3a5b94f72945a82d1c95f9d09646a055659c26a7b24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b8e6faa30c7784e4eb67e5077ac8f4c82223e966d6738efee7161b172acf16bcf341630;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1759479b610ae5c1744ad1dd728bedf116dc2f2af66e93510a9010f41c736df5c9222f746;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e71daf1c7cd02e98cb5e986799a6e6520404ecc1e5f8014fc0bc1fb541fe14068ae7eb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fd597904b26b5e140e7926d07006082316a957e226ce45bf93b9a62d60804e4018b790b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcad838add1fe5d8d554b407294d6305e6d618e55a590808301d5e7acd466e7cc8e43e96a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c91b3c09bfefa78866e9054054629a6394ef6d1b83dfc4e9c989aa8ae6ded5fe9254892;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4c7fe226509917f8d5cada24a8f45f4069bfee14e31e45c8f5afcb5672f6084c5551ea2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfda236d215b0304af0d37cf5d3f0d12c5ddfb5db265f3500c20b8a5db13902b311cb714e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138ff92fc0d9713f39437f319c0f46c479c9410bf34b6b6eb1fe8e2a8b69d881cc9fba21d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1783352ddf22d286facae1d5c2348671d1f31c5e3d1ed7698977935ca1656b45a8c762d50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b90506ea93b26018860b67b4643749fd831b5014b8dad4ef173f4d5f188b5a8933b6f52;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e41eff1b49567d780f5696d4b3bc3f9af5b84804930ce826b9436cc8bc3119745d90194;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c5e72920c84ea2bca02ca11be2cdd9dccd509363b0fd2b16402f549148f3f0c0405aa13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e6ceda02c5fb46fa2558be3e408e0155e0cd13f2c4e46bd70b6cff7a6d21e55129b8e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12268afb4766fbb25638b3f91e50437712b0522a29f441663e5c9c07feb24ab57d1f7b189;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170467cd43ab7931e6d8a3b6325b048f49de275d6efd67b5c6f5f2359f94ab702323bddf0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94dd5b01bdf573620a1d6aaf24b8b31e8494629a1cf2abd42ebd7e67c6e6de4fbd203ac7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f881cf4f00a62997e519d32c85f2dd0e3fe408b07d0a56c2966913222fb6b8832fd106a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2bb4b2a6621b1d70825dda5dd602512e9d64c4cc66301fc4b1cd466b48956072b2cb96e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c53a59cfd9efaa53dab05ad0cbc1455e1745a80209ab450b71a316aac274b54c46bd4703;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b967b1e0b454947f51d6608ae915498d002eb5e135a1b539c7adb8586611a037da6d644;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1672a083ce60f3f829ae4de56657d2c8d006065dccee5304f934750657be11a08f866061a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e2f855966ea1585694f75c75f942139ac67e03ae9b95112f7802f8d92387abbcadfab34f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb6b3b6906081c4132b250eb9350f83fcf4c25677ae4d5180869493b3023ce65d43f53d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ef93705f22fc203e4dc28d9f13f80949800df3ee631c67ebd59ea96de4660bb340724fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172ad451e70c8e7a38f847af26d35628dfc006cb1556cb12bbe11a16200bb5b5fa987590d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c912a44eb981a63f7f19bab25b47125e3704b33b3b3f2b403fc75edc66b795d392b15cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83c68c9b0ed4393693da19cac2ca7a0215c1e1cffce3835598e12acd8639cf9a87910804;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h403f3949e541c4434f877284e74807def408ba888f031ad0d1ffcb9ada5d4aba147d9cc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb2db9b24d45c7edc8c201b023ec72e6620fd84e4d15b87adc7da98a4976ce362765d33c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d99b6bc4357dd387f1e6c23a8e683594ba18d33197c246a0d86e95953fbf571f5c7ad8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e17a3b17114aee679788ddf20ab1ee3c04006aeb03ca7e3bae381498f57ee3ff4528a85c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8176e433f3c6e2941481d056f46d839b16622368c2f14e626c2ca5433776bd0ce79e2e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9078472bad5e0d62b058823f849d05097db48666823b64812d71c80bcf3176e4429bafa0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haefe50b7c6ef2750b74f2999d0df1ed6c0a61706469fcadeef3126fcc17977b501606b8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a29d46487729b5204c25a4a886eb9f1a8b0104863ef02b02b7f1952004791abc9fcaa05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdae4cc43b2ddb3159573c291e5ac675dfb0b83a4979bc5f7a966a4ef946be9812db03a29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc725b58be9c4836f508ce0f621186634224ca1aafcc697e27e28108fb0ae8f9d2d20d31a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97873e02daa0704fb6092e413c95dd6fb1147986030f53741399bb5eb90e7a83778d3dbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f363078882995658d69e76f8bbc5d15cbb6a91615293c1be0fcc5d384553f22e72bc5e47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h930272ceac8dff34e75bcc5cef6b11c91b222f7be7542f832d8c0d6becd5bc5e933567a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc07e466d7b15d419be25fdabf05b297eabb97cd7ef999cb9acc0d29df90ae97e4e9fced;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cf8eb9da455f9a14961377ed640d10525a0f71c0a9b38314af0d1ab0ed63123374cb877;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6eee428967d8fa10e870d716ffe373a86475ba6899a54aa11e04416ce34d3d213d6946c5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca38407129ac48544baf42f868eb0edc092556bb5d9b14c9a58f6e2e01c6f7f05379fe0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109f0fb1c32f115a79ae1213bc62bb9ceeb2f2eaf42cd546f225f8ca86c6750c9479993ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d301076750a32350322f93e39312b5391894b13fd1cd056e83db8ece25cf00e934439cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cc872b211b9661b971a634a0ea9bffbf1521e56b19ae7e7e6c538e148cbee4b0d2a5a8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a3ef48599d89892e178213df68a3433d9ea0e36a850dda1df65b0860045106c0c9c7dc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce4b0865a202f437cca453224c619911549bbd6163ccb25f447e482678c69ed1ee39082f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2509d2fcd5faee9d75cc8b01f2809a37e961a97046982682f88c990c5392f8c6f87815e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ddad74947fc6a9b0ea593bf62991adeae681ecaed62efd5512f6a3d838bb7449ed772f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4100da88231c723ebd282a983671128c97067462550d922a88c83db8b7ace3edd2e0db0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7c86424305a7850999690665054c05831160c655551296545a69d71df2c2d8cd4932b0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c4447ac4f48d124b100fc3665c92a18e53fa3e8d540c6e172681e70176c01d5639c133b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha46d622f59cb1040041fbcbb26264ad6a971f89d5980cfdb234da9d0a445572fc4649779;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc28224d36ca45b913db48af7fe8ae827133b2fcd6485b98eb33d40ddadc683947cde7a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d51e45dabf96ca7bc6a9baeec6543993cbc32cea8d8225021bd56d7b9eadfe8d01bf880;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e51fc1a43465c29ba23b76da0854b8ef38f99e85a0e5c0dac390c425a63be12763a04e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8e8f8313c6b35ab30eebd4d7cc89aee619584729e461e82335de9caaf19f0773fb6230;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1880d6a31121333f2893acd239a13cfdc062e4166caba8ac23f9b633e05447595241380a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c9fc469f2fd06f07a9002a0c3c7587f44a3941cccc02f7fe36db56fbe262eca69486220;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94eae5c92499ec22a5320e1a8a52280f9c8f9182a61aa7be6cf1d86bf51338b85a0537e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124720d029a05bd6d282636f18c6cdd3fbb44a6c96f04b67b16c525915c9d91044ee8a96e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ab3f60ac0ca6a9f702cc0690e94f611c2895078c73b3dcbf61350d4314ac104dbbf10db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he486bf380914657280f3812dbba0b5fdf36d46a3254a1b3608f416f2292c60d91ed4202;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9007f06c21e183cec089609dff780232d0fbda48bff36fbcab237832da523527d37893fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc877a9d0dcff51c648dec0e6f88f7446a1db2173a4eaf044408ed90c6faed61f6e5eaba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84aaaf30824885642f24fd186e51851306c676e2a46ecda5899b559d0f4f548a4b9c1e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113f43058fa35f4d019c258f9a80a6cc9a98d5ec643f4e4f0ec6211aa924da5280db774e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0b5c9603d9aca70134e283ea4e1b1936372ffaa160407b786cc5f04e5c515adf0b63dc7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9226b700630cc65e5f097ec6a33610bddd4ab7aa17661360e35cab45408e11674f361374;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfe274fb4b6a0a4ef9986da1766847017abef0c66c861082fb04ccb2f931ba8baab2ec0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha295e95cf0fc5a1fd3d9b924a228b9b558a7963d09d0a21d0454e43cc6777c2089e9cd6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126a3e1b000d38f0cf0e6222b888ce252067816c6e1d44e733b46a4701f1c1a17f39b2a7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ac290edf519c4440141061696c96c5ac8e75b5a62d5c50c398c9b3cd1b69cb1f2d006ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0afbfe5241d3d4d1e14741eace9d9c2418e2f437b93a887f19e3beaa8e500b780ef52aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ec3c937408eaa82760ca21c4cab57446fff705ff385a3a7e48f8e3e36b453fb24716f74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98d275a14e4aee0a6cc67dba6c64804d0d412ee76e48e819496fc9bd7901de9355557bda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1510131002bd2523d89a56ac88f1fbee5da492c6851bf867cc42f6251983e907733b9c57a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haffd9703c1418e1ef0d9fdbf62221733eef5ed735e9bdab3137d870eab5d28be51b2ee3b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d7e9e98d374528d919df5b2b806bf152b4c56424e033c03d73f6165ade51f674c250ba8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c547868a35eaa89cfd8a0bce7ab6adb568775eef349ce86f288fe85090d9cb13a15a673;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83b24068440380e56400ac47525dfd24b16840933d775509227fd707a6170b0e66994033;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c955371435dcea55520f673d696708d6cbfff17fbdc1b2ddade7721edd3f0c1e13b695c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd9f21a8759ea11249d60ff66cd32ad6926952928af4ebdcc799015b2dcab334ecf13b08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1f1515597d7e4b53e91fc5f6c37c17c46414526106dd4e25039f8fcc565a140cc33829b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc1bef0edf8237e5277b42b1d4bddad4bc66a123489a0be8979f003ab9a8306ac5e53d4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b5832dbbea4600e84deec7ee42bfdb8d65efd895377af6166c76742a9fe4eff2a4db4d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1873a190a3cf506be27769190b27a97405e2ebd6bb09bd3d16ef308048e395683e7134b47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4309de4ec7f363191835aca4b92290f9ba7ed532af7375c2e5f0e3e8ebd57162cda3788;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36fe8842271abc1c1c9cb90ae32017a9eb7921435e2404861c698bd3476849f6be9f3a6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145be49fa0c159699746f99d2e9e231e8b3339f6b17350a990b4a2403a286e482fe693aa8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f721b6ec41643fabf135a3154fb0d7969f289786deab5f4370362058c2c587ed5b54761d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1909eb0a8ae72dee1247755cbc049cb04daf59e5401da5b8c2c30cf1745ac124a21f38386;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1943411085cf1144b4b45d46664bb038256b942bc9c33c40c9cda46a6edf3ea9998731b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11db72110b73c0153aea4ed011b095dac3055de01cbf528c520b7be6112fdfe185fa3d07d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc38d4d8b38730693cec549e22df415f21624f656ec642d8c147c341e78170694fc9ddb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98efe7a1bc3c1c9e32e2641453d20cedff85b6e09e9c187cab4f91df0fce6a36e48cf9d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27c9bb495b6f1f2de56cf27467057acd0d0ab83b7c4643e16b49557751b7fdde9be7e2f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f49eadb8de60e1ebcb628d9e67212f4ecd4266f9b42869277bdfb2b8a7cc090f995a2bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197bd77659684c592c5ce0a95955e90166c10b6ddf80471b8cd5896b9a1212de2ac3c218d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8defe9c328ae7b0193b70e58a1dd4dab771ca6986ee0e7a4adc8766193d82a8e06d8d39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19540624c77259265b8b1ee77c66ae5ce2d005b97f1daaa374428f356db89d0327bf691e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4b4359b15bafb2e5cad67cdadef9c1da850e9e920a81b3b18f25f01cd29ae4956559181;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1020db8efb85340e591e2fababc718202218571a6a0f910940ff0d03a50173b30e8a3c2e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1431e085ab24b7d6a1619252e5bdfd0cc36ab1a6c3c3eaeb94b1b2d603a62e42b01e7f455;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4acb72b6e73cb8ff664828a84dc6a5bcd3e5cbc607a358daff5735d04bc6c961c7f39483;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8130b99fcb7a372f31c2610b603ae50ce50bce54d126dc645383c855e25b3cea325ba9fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4425d92594058bc8fcbf843cbc6ae7bc9847b18dcc3d011ef60537d02db350b9165f5db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96454f9a7bf5498efe1f9c3092849808bd35de7b6f5a0e1651b2326e45e5d235b43162f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f1f848aaef0dea25503bc47260471d7bb258485b190c241ab4d1c7cdc184cbc80c59062;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2c6af7e0d742ca97c29bc4c37561e65e0502c8ef217b1e48749fa566e3156e9a40e7a0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf25339239c429bbe32f4d970b87661d4d14605f99ea6ad99daf2d0e78d8dce8d35787d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3ea12797bc9c15b3c0e6b24a2fbb8f4fb346cab200d364320f39c4f3443264d61fa74c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc716c33960f325313a3f795acc148a7523527e7256d1dfb2b1e0e8ee6f6d7352bec6f599;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he07ead38e2d5ca624c6c5060ea7e9c1b3f9418fa5fce4d2de8c9644844b0ae8d6617a96e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc6f9e37249f38edc818e25ff6695e86adceaec3f7df133c04946c8c4d20ba6f19f6f4df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0240babf8c57e5e4ee49d147f7f82408f9d421b3fc9a3029a08df8034328b13183717e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7ee820cd12927bae2706380a5ada23cc7e6d199b3cd4cdb5dfe5b1382846aeb6a6b1d54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112cf4bf7f9c46ec6e9495f0b5b10bcbf2fcea953951763ff06aa2f3bfdbb1f4703274158;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ede46fa79b95a88b342b20437d452101db5aaae2b049a6bd1a3eb42480bb49408fc89d55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6da42bccbe8658bb619a70758a820e54a5afce35544773b7c83e22a8171070195847dbb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88e218a62b9e9c6cb0a3c1a91f1bd5b9586b14c64480be59d5a421ae9a8be8851e1e8433;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1099051a5f3912013071b6dafe0647e6443904e27dc7fc290fa089f6a21c3a655a8856ee6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbddee51b8ffb8a3edd63cf985e5d0f5553d8b81a968ead6dc41a00b1c56b8680f601c714;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c582c1ec0c52f20103f6cc8363fe0b9f23b58c6a9c8a4be51a4ade066ec810610306686;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c292202851e87890f49f640852bafa4d2bbc469be62984845eb9ef898dd0bb5fc5417e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ad721fec08521d93fef09466d85a759f1fb8326adfd63108f8c63f70b0b79fb1a3cb906;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h893e6b7d6da9d3969aedb3fbc6af8b810e106c3e554f4df2b3e1fd5d502ccf6e987daf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d64a6a61b70548488c753f2bb5b788803de8129d8d47f8a19f347b5f3ad7d888b960baa9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd65da76190c6947854272145134a6a4228531adb9c5a89f5da3da165eefe997bdaee041;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed074908d6fae0ca00d3dc30a693525c983f29a31be968f2ae4e03b71ea50c7646efd493;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173692a55d2958312ef208f3dc17de3fef1df002dc089c2524b9c881af7202346e657576;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136c90658f7cc0bcffa2e14fd1883a829e87002d6f233c34e3c115135f4113a697afd5045;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155d3e27ab7edd632e3387b3bb81775ff7d8618e36f9fd0c9af6a626c169474e9af0f49eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1e65b5b1df904a275266979edfc337cfa6b156e86825388086ed46544735f0b88b5347a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h871f35389f353eb8332e6c5ad18c7c27b1ac0c6e7b3b13986a6862c95e47ee776e76431b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9fb9c27a136a9d68133d1a6a1567b6a775a0656f494f383562c2633b831f7f3933b8fc8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ae0ba0a6fcd017c2a4a02af7bad6b2e540de92da89d69ad429729deabe8fd97da172bcb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h781919d4683a3f9276b3a33836c8d6535ec02931d41d937006129406322f3ded90741111;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85a8e331f7393c9d82c33508305eb353952b966967d61c0196654bd9928712268f515816;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a160296ae86cacd023c444c91b6349a3ebb3e257ebef0be938de2a1a913e12be1a66bae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a00827a661bfb144491b054b82c312f16fe0218dd82bb976524c8e5970c0fb11bb645fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7023584eae4df777c046a7a38aac5240d3f0e7d0172714486717f010758c8aec204fa3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d6911d57df7cc8d18cebf0e198bd6c1f5adc61474237b53b83f443e3b0ada8693f6284e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c06b991f8d0b8c4c99cac1f946bf224f9f87c1642d77bb4f664add04b89c210e428a4b12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb118d61fdcb8a5721334e46648663724089a6f771757bcf2ae0d9e7d4aa6d10adbcdcff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f989d72614cc22df34af06f5ce829bbdd19c3dcabf8536d1377cd5ffc56cb8c612c2950;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb5bb71a55389416a83257e7ccc1cacc52ab62bd77d983221a3a1299e70fc8bdb04e825f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e99170aa045edb6b85af58c5af202703403fd543613459bc473f8c088eb877e759259bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b244e5d276218424363ca2abbb4acc0008b65d11fea1b259e200a044311cf381f772607;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bde5cf6c038cf50b9ba0e542b25eef5f1984689ce6f4769e04004a20fbbc92235fe019f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf035970fac21861b5db1a1c575bdaaa245a1052104eaed9295681844d14814cbdd29a756;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140cb9ba7e990320d8d3bd2c2a374e5d97d0e22d00f709d89158e1bb5a0efc21a188dc151;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h335caf747dbf7ad71917d1f2bfbd3473f637a9f6af3f248fb91e31292857e9c6607a94c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h229a0ec47e641a956dc97ecb68082910daae4ace340a2f8ffd897f02db55b40a28132aad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcad5342267dc5eeb00f22784d163c000aff053a4414dd2ca424e15ec503eb7f36a6eded7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f30857d32d513ef3459c2b14657fae3286bb59d24e07d47dfdfafbb18555a98643158baf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc3a7b3901442828224338b9a42c68d2ebbdd8e000272f574a0e3e28534ed2608ad4daf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16526619cf6599fda5962949fc8c3fea96402d2250c553b2197411820aca23ed74f114be2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b53579ba0df086fd05d9978fcb49160ab099a5d9eb3cb83d7a0ead6ccc08fdd5300e5b54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8707f767c583963d50ac6a3a94cc15ab4fe46e928d0912c350dec4ad3b475dafb05ef8cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb479c96eb544614791e65a05d6759d8f1b5a0ac098b5676923045c690cc549348030989c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h904816780a93f77d11a70d2f408861a4a9c83e8e3e3baaa1903837c9d1f4fb5d3be4168a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1919c7f34b15fa38dad38289ae1c4b3a8aa9aef718a88bc10e6ccec6dfebf42e6762689d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3168fe4be8cd2545fc9b42b706200f0a82413d8aff872ed65a6d3c9f294ba819a6653aed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1777b310e6f2e12d6ce4444f0de82d2adb8871f5ff0c99384d407926e258f05754988e52c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4143460d4500bca70ab212e76f5b52191b0fcaef4d2482006a42b615cba5eb8d7690e0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9223bcb44d31a556fd18157f5ac079afd97073bcddb0d744c0aef2004ec1b32801f6557;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce0d61f70e73fa6350d0ef9150c7b1a5610d4acdde51398f5db2d889ad60128cc7c0e8e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2aafb86719c051f0ac2ced9754c0f988930e5f98dc59dd4211c3641b1a46d453fff773ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ee549b675e82dee98379682fc46ab08d787c175cd3087f0a9091675b7972b403882455b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8c1d9a7f2ef62865a5392af4e60df6152ff544e8a162fa83509a5e591ac27b81a3a3c99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0cf37063e5cd99007de891fe5a22f4852af31ea459d6082c2c375eab4765a8c2be2534;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141900214e42521a4c5c930ece0505e426d41b21b9b21227088cbabdc18cb18ca4ca9286e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c794ddbd6eb3967eddeb201e7839eb6239211125efbf9644e69b2f715be0c348663824a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94d316107a8563725bf36716c2b4dd601da73c9e6706f80220e19126b2397b2c28fb1209;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18294eb4cc2aab4dc0f18ff1d244c348484e6156baec7106213a9807ece9655a4fb6d9b74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174aa80f2f99f2a4679ea779910475cd1f9de2ab4e088864c085aa93d94e162167c48977b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a8e6f5617fe58a79c5a0c10894c0d221030d1a8ebd47e4d14e6081b8117018dba471657;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a58b18e937495390c54998b05502f9c67621a2c34abf383d353349cd88e6b5fa0f33f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1011eb075125265e960a6ed37b00ea6c21c049a67bf8f1367696e791dfef28ddceb4e9bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd18f284e0a87ff84fd4e1266fbcb3db529c20fc4386cc556cab2b5e073e2b001005d1c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c987467ec802cab1118fd561eea59aea07af0a1c40e91b4f6663656b2e37d884f14e89c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdb79c8a6e18cefb03d0d65ba927a97ce8627d862d3a07ad9c3cb30caa5d55957dbd9e2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h508f90dfbb0c7c2319e224e24cff40e363ac49443d85e2b8fe169672e6f483bca96442ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17611053b750141e5737cd3f4af09536ec0396427ab7b910b136142c319c41b5a0c836fd4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107a4eeb667334f123b38c79396a4288296e3b1186f27700f8c0da196b748566dde606412;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88053c58302b00322c272a46567e307764ef0cfcb24bdd652f6dc530d7ad1dfc02897921;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f84b16e5ece1918b8c22d14f55565f8af757c77aac0f7d0158775788db44460cb715d37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1411993789312687571e1159805218eab97f14b651a1e607e62d461049a8c11e09dffbfed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94aba8d22f29058e07703eb8086cafaaf3429d974b384b02e6816b46d0bab0426b8a5800;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5cd42f95b9cc97804515c296c227bccd7983ed2b1ca2e4646f390caafbe832751b656dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h327e12f313423945a83744f96f68efa07c6781beab149f16cb5f01e2619a5cc0cbe4d259;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf14b0b0061dcd9d482ed8f13c7c3b49027a18ed90810847591c5c4b48b99a53e2837e09e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123a9296318ab528ab5a4a297f8e3c2e1069b13b162ae2a9f8d56d69f207a44a7c9b027b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd04e0218f0b563a6c458d2560dcaf8b6a0d0d2d97aeb2da50a5fb4e99ad7988dce4b04c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1474eb232d55de532f9f84d41efdca0a950573dd7a6cd603cb8317918257a5c6d9507521;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9a1e778fe3231c04a7c0c37bb3a291ebfdcbdb6048291a4bf0e3b0cbfda7f13c0b4e448;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1227436eb0ea344b1b856768bdb6bf0bcf9b9c12c7063c9595c78de7b7c8a2e8b8900be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1167049e9960facce9cd4c5a4b3d0d9567d3bafd5eab933e88946516aa09e7de1d127ed07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf645c9c820622bd4cc0a187a60be1b11669081283167d83b66938fb8f2ccf2e5257de0d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9709d1837a19c647a31a54e4df5f84a9f722f8299af4ccddf7fa7e1818ef2482f2b2fb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170be31bec6f009d57ac93b0d8f227f7073e85ba966f32f2ddb98a2a816a38e37b6bac822;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae922015ef60ca6d7f45f54887b6896bd94074e84a99e9caf64049ddb009597e017ca145;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc31071d56841e73b854f2168be98fa638e8c59e621a23151a62fb6072067147e86cab6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be16f1dd3478958b171c6573b71829ceb4e9b4b8af3886d0410c0cb1959ded377f218703;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7c42c3d4b2c0946de5625cb523412afbee3c5e0f31e1ac95f62487c81c29e1115dc9254;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81b2033bf0b38d493db968fb73374406c794d2ea0b836d842f86b4c39b2b92854b96d70b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h237b2ab56de8d3d961326a9b75e4df1a5e0f224c4fd11f1f339ea67355c44a52666e3f53;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135a77f9c14de5ae5f74dc203f016c2c3ebe35a2e7f0e3eb6d5a3dfe6a69c12e64ae207ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f19c26a2777835261b21e54af8c8c9ff6cec846e99019e908f974893ec9542c860789d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1594491526f30fcd9c13f45aa1bb22abc6d7eb1355251a8eb2a49b0ef660634cca034b071;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a7945efa11dacdc0b85a37ed82b5d3c247e309ababcbc575b98bbb79268a4f7ad118355;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f2982806b8b8a5dab194eb7a4ab4cec1d7bb00bd2f818e3311a3e63bad638f4ac2e018;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab2b311ee4fce0eeb625718f7991d1dfc8bbb384e3159b19c4e7e973418c7d594f1797a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7490df7da043c1e7616610d59928c0336cadb16d88ff192930e1f6d554793556a6da6ebd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf54021c4cb61faa803a7139202836936bf22c712cb13cfb36a510130f839621b641b948;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbb24ce9bf7ddd998740984afca7b2d1d9b103b90a0d72bd7c705cc54350eda141cc777d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49058c166d30cd0f7cfd7bb90bab6984adac644732f0915e2ba812540b1072f91bd7d5b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179c188b3264086ebd7f7f8e3ae4e43aee9811d41421c61d598ea4049e57adee11f94bd2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8a15c9e6a00365e10df8d76a875ffdae130d06645e83382a589421cb072cfdf899e5a60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ee1c4d9db33d7321503db8699052f98eb052db6741e1c41f7ba5360ce8f5255f4f7bebf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha93451da0f229c6c16615770e9482567973432c5d55332950a196a4829ad14c326bdc15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3baa0d7a6b1ae3b237020a8372231d5c232c56231a30fc28485f3a22e4d0eea59490bfe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b464b8ee4988799e1d186d53e601ee98db134800777a897b915c0dd9c7e26bc54442467;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7056c7c00157c19e143a906a90e883e9edaad4d9b059d1721f3b5c84d2c2b5aacb01456;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c4bd8a655d33b75d2b46d1480bea2544a323236038d0eae2084977580506809765efe94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd80f0fbf1916fe1e734ca752cea617d848459cdf62d6e510ce10cfbf225c0d1f968cd2b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ca3aff25dc8223f7af13c9dce348f6538a23ea3876dc820adbddd7c23c8fafee8241c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122186eb06bc3b320983b991e59119d0022f52cc358eed52967e09bc2d72f37e0503a6b2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19085c89b950b62da9fa648f74cb1748c3bee0ac3945625e3b1ea69bf32b84c4dcb2c865d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8af76d6b75664e660a083bf4a7baff4a7642a9f31a302099293a2eb3f04e386faf5f1517;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16528cba7f7c41714216560032990310ef464d6c6b626830a720490395f56783e0815d1c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1588a190f9fb7c1d7e02cc9f6f2c0f0b7f62a3bca93463b53cd3450acdffbb4096f28211b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9729a67daa4b5c18e81270ac89ae489810bbf666add069813f28bcc5a11446f2aa2a974;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c0d13475ab2c710a47fb6e1e36953e5850dc8056cb4c96ee81d0f2f2f3c0aa6cba7530d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8c8d0492bac3b48f5662ba562494df711361fdbf3ac2b3c495f369d67e0856f161bb1e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb627f76c993a70bd12c65b3f8b639056dc653ebc82c1e65917f305f0c735c412b37f916c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0b3bcc86dd8be21a60d409da592b85a5de63f2e429b27c55f293f99b8f7c2d50d860910;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h867028beae391ba0b652c67d6035efdc9a795b1457dfa64816e4b8a900b352ed60df6a13;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122cc0426a45fa4c17d515e9aca960f77031eecb5828f9a2ea11a8917fcd6826541704767;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1009c379711c051e93da7737c2b01d34d8793019aba04c5e81ecd653469e8729ce54b5fd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cac8e5e4f8ff0ee6a62d889790fa04a791d5da29391cf1d94a2b69e4ebf15d7857e8e60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16bc2202c2b038569efc9c9ce397137a11616bf3ff5f7d0522173e4b60d113718855fbd31;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6e15d7ef6b4e2e8dfc6975a444cee5c78dee918a574668ae39d3479e6b6489f7fdd8572;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1437dac58689c31aad8e8c38400986648076a9db3fd114fd35f3b8976e93a89bb1d009586;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c1823b945b8cfaeb307c966f10bcfcabeb866c0f288e2665e300aa471eb7bf67fb4bee0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164f86c709bf1504f16eeeabc66e658e6df75932213bc9e08040f197f2b216d0622b52c2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f91eb62e3214a1adfef61929ae806a8cb568013470096c6042295356db68e54e7005e5e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30e752bc461f583018333d7dcb5a54f91b967e110f208b0feb2436fc0a055a8fd43cd588;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1864da6f4fd8b416643cc31f8ec47429cebb000aa2d83932e53b216c70767c54d81eb3e7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h455487e242fca934841ee273c36b3b001d1549f505e07e463cb3c05e3b39277a589dbc6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb496968bd12c5a1da3d3fdfc248a1c601f46d25411751a9bee85b280c8adf70b0d9e5ffe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha68f9d024fc26ef9aec823f44d53e396640d1a34eb2b7c5bb112a55fdf706815cd412740;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120ab374e135cf44603c924066f1aebf4b68b9fad1b85d6c7f915817817158687238e0947;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1671b1f4d1ae3a8f13775ad8778c02fd3f6214436255d555a93a3f61c97347043e9062769;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heea4dfdde4347daf3e999df82a54cea3d6ea64d447d2149be41c7542aacb913cccc7806e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173caa030e2f63f5618afb07f50a278836c466fbcdef7df66def5b0812574fff3450f7db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22e5547b81fb574d20ae7514426f459d41aec51a2ce8cc1bae5bf07ce39f4b12409c1ccd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6a8c89395979c5f2a26bd9bbce7c1c31a9493c5b0779cfd3eadb2f0e00e4b02a495de91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3ed81f429a5cb901db7c00dc1bdc4e0b66a0d8da33f78e057e72f7c5d6da9891675b515;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1593424d798d0d7fbfa84a14e961de0594820aed59a88f7d425f0d00aba08e51ab0e6fc9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45a3d25af00b263cf3eddef19fde032cfb3730ef0ee42a6fccf6e43af7db3de0ef29545e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9976b35fcadf06ed72bd215ee65975fc61917ae21604f12acf356993a488093dd819216;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113eec49aa80923ba9c46511db11716459e78fec5cb2803d554009a58f464d2a2d65ae23c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8570311795abe298e4125fca5712deffaac3268f338f8fbf1e9a05a965cf407b5aba5dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169ff914dc88df35b9b39185533d3f777cde8fc2b94fb5442f5b05a939c51d8ea27511748;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h661a4095ef0b6c291d4dd79db90397f9a0109c92517c8271382cf971c8ff7440d1e8f2da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h582ab37b0cbbafe613ebebbe81063a265efc7cec4ec99692deaccd9b10029699953019ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h571217070bceaec98ca742b46ec18f261b243d5bd626e68c9a2f4963c0bac34303a791c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed22609d3ddf4a373b16cf520e3e01b3b025eb074970f19edf3b4eee95b534ad3422e8f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c0daa26fc91e68f91a107c14717255fe7ad2e1445e9906d0754a12157d84eca3916a58c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38c095d64b7f0bbac3b1bd8813729362f9f35e381df3332a124b7823ff8e511a0f59e00a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4a36d68f2155165683b1014f3575f7ba48e5482e3ab82e4f240a1a1d5b1111092b44f6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7db157b7223788770cffdfee899b9c8b106f258c833d6197783222d4bab8156f8d1c1fde;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1546e5b737a90cb22d531fa20a635b40a0efab92a4f16bde67dbc8bcb0ce2237e936a4801;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1449350bc6920527a502f51d38d1ac6856811a3ccb4078bbc5456c96ae92b18ea72f8bb1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b064a97a9c9dd4aeced53ae901b5647bfdcca4f284cf7e17489be60180f862781b06635;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd8501a5ab6dc52cdf8ee901b28c892cbf3dbf6e88737c51973f3b4bca07a74e60cf3aa4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8282fc24229109e6a314fdc014acddf05c8251d3342c9f5c758ed2d74a1de7c737774c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb854e2d88a626cce7200a54bd636ae0dc1440bdfa35aef948154b2e5540efe5d4ea1d92e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afc3ac046f8ca7479d69722e4933f409f2efc09ce1bfbd0858e00e2f68ae634b6bcf0892;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1016f3cd000a712b37905164dcae6db39b5ab181ca98cecf8cccbd8491440419b6e24ca66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd146e07a356a4af83bfab3904008a645bfb89f4b873fae09b0ec0ada66950d5203dc6f78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102589206a602aa6f889632530b1b50f204c07513f039db5be70a1a571f94089b161eee49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165c9f0a07a0caf8849141dba51729315cd26da8fccdb77838251c27778d9789db4496d92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb489d41dd353231be66f3763bbcd5e3471edaa7d51e6b01cfaea80078fe0a43c16620af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a854b5051c15775cd00e13b8073d616053eb331c5d2d5897fa571ca1b04a7b6140da101;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61b492a5948fa07ed63a65bd25da233d2acee88be5b39572be933140c1bc420e72f686b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2464addd465b1a6816687f26e97136f4941a037318cba324e7c03674e5725f2dc3024352;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a70eb49868836f1223ac544b9811fdf49a46737de57cf9be2c5b886fac74621745bfe6a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13eb9e43a01c841423cf742c810b0262d88065ecf9753ac7e383aac67c050763db5816437;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cca5e1f3317217fcf5878926b75b97df44ebddff89c9ac8583384b00991475a9def4876;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49fbbedc689c9db8599d87b35f4fa35d6b562bd92b851f07fd2633e4711a9bad67e69c7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf65c456dcf01c78723556c48cfaf5be516d24ac441e8e6a6cc194656dbbef1a03d708af1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b368b9087d575ebd2ec42b891aab1e1fae67ad5a714103455700c187bf80ca80399edc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149745bc870ce96e4472392fa9d2066e136381fa7dd415ae8be2d6f51191a38c3fe543184;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b773ad6fbdce9d2029c80888814bc7e8178e0d08ae10a419c3130a16cdd447f9f6fc640;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f1d215639507e5f75dbb7e2d0564ab849b87e029d1bf0e84b0a2ae99e87924c49c233e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf83b9a61ab8708a1e8a05ec48818d41fbed854736c65d2c5a21251dac872ef093c2d134;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c31feae31cc9068d395fb4eb89383dc42532667385354f0374da9469b9a746f17b53f58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce10cbb83affc619f2bb85de2fb9027b0f26b3582d33fdf1f5ea139b8a5869f3d414de7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1122f78cacdacc92c6c655b59d8e7878242823d3febe8c20591c2a6cc1dff7a96bb267e47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114106dfae8a1fc2b86d8a283501409987a98a3a5c4b696104532b15af26eddd6996bcec8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a22ea353a61fedaa5a9fa2092f7aa2714b458e92a52fd37fdef2af7bf177cbb7f67aabda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb8d09fa798e383bc697167e165e875a752f86e392da1764e39a89e917e4d5d71488d281;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14de61a6b1f0b314d61554e4c2a327857c0bb200aa308cf11b533ea49620bb70b45b57c0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1b0e67f80c35716858b7f846d9bc1398561cd7dee0c1fb3878e4d426cf19eada5cf1aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fc7622a221b24b97c9a99e27b4869b8710e33aee3fd1bc439ccc872970906002e1585d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h720cb95c77f99b6177df17cb7a965f7e6d301ba0b3edccb409bf49aca619db337b8a1d60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a18017e89ece352ae73f0b9d27f038a18f9010e8e88c099cb20599d3ea8c84888825964;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14dc0213f8a49c921b18b3660065aa1bc10072cade8c1c42fd99167407b6b7a37bcb708b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3715c69add4c2dc95afbb42093d1fdd3bf8f577398871aa4b956d1cdadb15b9e29c50094;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11f48126a494ec1c604f404849d007f801a5d6a8768708cb0cbfb30ec71f865ce4f1badfb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a375e83c9278d29501ef1cd4a489245aa79b5842cd83b345ee8097ce781a6b40df4fcd2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36d1e2bcbe262272e9a48a191565ce7e26636bc27845ded694cea3402b17452ecee63e02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b3d621902c20b19f419d560284cbf26e307ae26b6c9665b9cf45c554891a724b0fe1a6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b619772b24a8f6d533ef2b68cd3206cffdc3b5baa6033158ec5113c24fed9f8f3268aed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de4c31e89f5283c3f943a60c2e66a352df3d2830f1d3a764b79402425d73641ed7a0a444;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17798f63f38f9ee2ec55ae460ef2b1896b4b11edd0ae0889593ea5945dc724fbf5ac5a9c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbdde636c11fda14b24dc01f0b0496ed7a31e940b9774cb18e19396a7f72c603c0cca1d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebb2d30cdf09352db31d04210ae4ff7143e6e81edb4d45e0bb284f24e35bcc15f85ded3b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58a8bd6b94191198957678e81fd3ba01de482eb3ebc7e46fa1669a3c4578f39cdf280191;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha17f0c7f5057add8f39d02510a9862cf0dfc0599d100a972f595a5c55b3a11505611da00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca33333cb009081f8ed15b616dc024dbaf2704754cc56f7e7386349a6957b0af78b9e910;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2a4fd591e467dded9ffdaef53f4a6cc06a20254b13dfa7a743515745eabccb323058156;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79ab74be6efd7c3fcf353bc2d9b007f0f682cdf04b9bde9e2ae89cfb3a616d9b2b7b59ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc997adc3d1f97ee16c630376f616b3fabd1aefa87112bb52fe97f0cad180a5495c0ba633;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5e8cb197099812110005c2684e7d1d4c961adf9095012b5b769732f5fa5e49434356e0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa3e8d24fd6a5091dfba12121ed84b2a254811ed21d63b1a8dba7109593caddaa62c47bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113370a726fd79008f7630a337c6ca3de8250ae0bc285081fc9e37e2b23dbfde61714742a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e20d56d656e7afbda905f4b5ffdbf3fffa311e06ca3d5b9dbc11a8fd31bb013df0c73334;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ff79c9c14d5223ae8ebfe342cdb0262ce3793babda23de358d5bf3ff3b412fe0ce28637;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4435da049c12641400a76e3113b03998de577b76d46ed763d43f7b0defa33316680e5ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1603303a6458700a14c6479e2cba26df5ca7be5d4656df5064c4fb3fed49cc0236a5b0346;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d004d650aa71318d36f79430229d5764fbe63d08a7bc8c631dddc7a5c9f4a352ada47e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9b552f2613839062d637f597c65c2f0bbfbd235fd23d8011ee812fa920dac01b1d9311f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88136d6844907815ee6abdfd162ebfff3b1c3c57190bc6846c777f29c4b8e062e41ac939;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbac043d550be06473761bac6493aa9cdd0cd9cb5c94d95420279b7913535d660f501bac8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199f235c39f6fe9cba837676b28bd89111f6e22c25181ae8cec31d9ad7bc1e98f0bbddd51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdaacf720d709674adfd19ee41d311cbda20acbfab5f6a3d15725feeaee53dfc96d8e0356;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha55fdc7730a95ebe2764dd89b1882144f5a273376ffd681fdd4e58cfcef4135315c59331;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d90b02d24c180e4b52d9761240c5eb81593506a0e713a9e76538e6a60b99a191f3358f98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1c7897b427df93800a342813584644f57412bab4173a992b5c184931498ff50f28ae3da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39c8ddc13d509ab19bc34d5719859f55660b4e4ccddb7e49a999c648d4a9737c23989837;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186a0e71f1b86726ffa14a5b19c6f03da85c06f1038a1b594d5acfe7be6b0dd5ddde55f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebda0bf1281bb8d36600ed2d705207cd7e639942f16439da7df47ff91f5d9d5ef0a1741d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9cf54da1c670d200353295637468579e738c88110c6f8aa74c352b228c85b8d76d707208;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf7884a6f5666fbac2609748835a702a0d9ed5b60413a698cb44b2a9072a7d01fb72b1cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc340e35745c4dbf7183af4d46667719afab2ddfe863517323a3e111f461ca8dd8623dcbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d60f08a9f5b93f5cbe375a2fe6941e046577f69c33a10014c1dff7b1d42e95a6b8ab074;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h631e4521314497c46751293eacf03a40c11be0ce71539a0672ff9055760cd71defaca364;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b6cc07bb3dbf4830a91ff8cf4c101b3cc0408b7e1cc7ae0858a6683d2b5acaff4b6c88f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc4eebe2f39134655a267fa0ae4144f48452d6f82a0d341edcb9c40760078a458fd469e3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141c4cc64fac8b0f09429c337e083ad1155e609a5f8ad902f11bb976421d793f762ac25ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hccf05281a151019728ad6ecdf9f3e44b428120607514bdc9c39f3190c81d5f5638daf142;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170272e079f5403c850b9a9561126774240c89a3bb01e6867f5e7dbe1a09dc57075fddf6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba79cf9780abc5c0cccb7f5faf7a84aedb7c71971e2692b52e9276a807110774bd32f90f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f21738c8d5f2d07f8dbffd3dc51e89ad2d0f841419726adb723b5481e79c0b46b4e4040a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15de874648ec859f7ae0ff03adbeb692f3e499bd3a0730da3a1ab8e5dd29f72ce19240e96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbee096b2cdc7c8ff39316cf66c1ddb8b1e27c31119a434efc3ff7ffd3e25d287da1b1d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8803d9b35d5a5efbdfc578a45a982245cf90a9c660708cf971a77a2ddbf8617b8fed75f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9afaa1717dd345ff3def262a8ab5159b1969b918808bac9ae19097078cd8819358a2a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a5fe53a23ee7f588070d42486061cfa8d7addf386b6a07223d9e29a75ec54176eae177;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h827c3c2ab33f2fa7324c05f1f334132c08fdce31d67f14b7aede41633a0d57e67fae0cb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfbe2a7fec8adf499b350194ca1bda83beb4b6bea3874a95ef52ec7de6a0b9d1b8baf12e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154f01bcd1a89d3c26b3091ec892814ea8bbb8c28eb63de3027e12d5555b41ac3de52d1b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c677599347d1588cacb3000630bdd7d54ee8beaf1daa15010b700967ce5920b42f6def48;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f122b6e70a19a209e7e618cc0c2fc81545d9b314f428022d9e396e6a1e751acacfd91d9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115e0288c96674cec09d96c00c1f324f63a4d6695f2e8f68d9d4818ed4ef7c5a3d52f437f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db645f57f9d3a848f77e8607ea7ca4c4e44dc7855d9614054aeb028d2b5cbf92bbfbd79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b0ae1dda846ef3f5d15b467af94a2b757e41586265f40cb7c1e488b07049974a5c3a890;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15eea83c5ca136cf492c37a1f4cdfddecce748e58d285e338e804680769ed48bb37a13ab3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54ab8f900c2d84b0e1ad26648e8d25dd34f8c20b855d90dac34dcfe2b3b167f045638706;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9f2127207c4b3ef6f707e023467a4534d5ff2762ea53b0d9f0459af9caa07327b9cb538;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h463ccf2a4457548535e9de1814d48e9ebeafac17cf42c3219b000ceeac024809e11c1edc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165903ca263e9234af48e9873dcf488fc3d6257dfe248e409503ff5e77814918c8a387d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h335ce32ab2af02370eb9f5fe25bdeaca46161241e940c4de949a02ff6b72bc75447ee78c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61f3b09d3fc64a59e2a64affd2cd9330af8835bfe06ba1f54f05d696f58f526a240aadb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d3ba2820129abb13af73a5bad90ad01c8e77c3e6fcbce2d7e3cae09d03aa4e4c2fcc2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1293b1162efe03a531c34635f67cd605ed52a9c73510d6074bb092d86d94f806d432b0b58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e3dc2c03e4003f9778df8cfe2ef0d2ac3b7dcebbeae1a42c47fe98e88abeafbab072624;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb846f7ac75ac3b334496184e801777b14ac9a749160c19590511767b0888552e9af2676a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6d969328b5f42ec13c0afb316a52feafc08d7bc61c9fb1a0ebf72252ab2e7976b292b86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c8aa47185bae88a0f06947cdd9182aca84f9d49cf9f992d3a019d3991ac5f50bbfa2277;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98f52b72eaa17bf84254c186d5fe7b458c7540fba0c9a0bba5e4f861386a5be5d9fe6bed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h818f01326e7ac2e25f0fc35ec4b4df46857ab6af7b4fc6f4af272eda09fa5f4fc1014d37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1723042024c84f85666063e136a6fa6d65a1b8a1e6b1166d197ab7544102627cff483bd18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h472f406033583cd6a79c14d38d879ce73f1f49df41651366494fe2dc152262aaf0974989;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3399584f71c8c28c189f9e98dcd2163ed298ed0a395bcf3bf947da4dfd314f25c84e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11248b7d0d264104e8c14cc9ede2601aa8b17eace95a442412bae8800cb310545040bbdd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf011d86695e074cb4817506b5841e941fe3083541bab8a6332ff3e29920f1060bbc4b30a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7938424d07620d2b0b1f24c236e620772d66dedf8222263b9b74a4b9be4d6608822394c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7d7f7d0c6d02aa19c7dce0e5be4ee07e8034f15637fe92fc4fba4547f28bd4815b022c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f5262b8f0e0fdd5ddd28824a672cd24699a3054e47538d27cbf6f92a3661e29c709e328;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha92d599436a4ced9bee30a6b176a09b6194ddfc8dc197a0e3afa5c51cd2b0c91ead8e12b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd173b67a705c6c14678ccdfbde71829d7ad005d51a682dc471a1eda75e1121c40ad163cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd740a3ea14ab9f4bceaa0e65aa2151f3a7f74340bff0a8c35531d7680d398cc0f8105aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1543e935dbde06156c13211bab770d0f2becf87506a42f4b3943a5cc7c360b480909c363b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168d8e0d4e2e8c552dc614c64a7ce0819f39f42f3592a8ca5f1b791e0679b9f955d3cb9af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c68724fc30aa72fa60d7c9af050a4c45c1e6d349ddf305bef67d3aeae544d83440b731;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19dd010fc2bbecfe8e661483985626258385324393f77152eca197451622494400c33699b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12432ff93d04ba73d177f40e897e6326a6777e6f2927320ce9a9e3e83f4e6c6a5be2ee8e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha48727dab82d6da97ce3a65267d4fdeac90521d2df2e3a3435b575191bce44268e786858;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fbaa25343350a834bfdef7c6ad2201a85349afd2022f64d3b3acbcfa10d0f6e547e29f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126350b71fec9b4fca639d7ad1367091b70dc714f568448398dc7871b79e9f449f8715cdd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac8fd10ada13bd7ac1f47b070b2101a2f61a13d698820f4c71a612d9387429db7b13f0c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60878e6c77a73bae7214748e6e1f7297afaf102f9a0d7c9704052ed74e8e631b656dbe3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd84dbfc51541a2f2b8fb0b6ea0268d7537551f86369721b443f359b362ae5bfcf25679fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dac6854f7cb5410e9269446709bb98d6fa7ca7e852da6bed695b98fb8c50b09776f20de4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bc5cd84344608f56631c42c3a271b698c9c2be178f1abc48c1dbedb1dea97e6be030c4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c84a3044923312bcfb2675d0307079b07e3145ae372cf95b8c7237fa4444582fde1856b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he13774720218f340611ef17b3f8fe3397ff5aa74de943d834eb2c6c7430a7d6b83a3d27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a70f10472428b037fb40e2d4b19260afed2e2ab81282fa7ce063bb7c8b928b507b6c2558;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1accb3ce9d7809258a0298bd4baffb3f0d02d0a3fa775c3f01da6b844ec92a7780cddbab5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e305081eebe6587db3f45925fd3a6c790e5394bd00bdbf5b909ce714fc1afb84a3dc289;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fc66acd08633923a9046a37a57a902eae3cf28f480b9ef8dfc183b49a682afa1f79645a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15edc6fcc329ee7d4972a3f62b86ee48f76ea7b4338ad84672b648d401fb1109df4e5a20;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf41e26e0753ff2e3160748fee3d5adae06fa4d7f85881c028fd44d195f1a30a34d2a9e68;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bc424f5628b910f4be8c9e0ebf7d9534e53034c791d1a0d1c704a6fc4fcc3bb7cd76529;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0615caefbcc4cc9b59221ea39f32fd881ca86308243af78649272e02d9931e8029579cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5961cc022b8e83c99f4c1263496685b2b33b9c009ddc36cb08705f3493501db3e37bbc98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77b1f4812432ef875972151d08369157c9fd5efeb763f77a3c26d78a7c83638297f90699;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfd63d93af4ff09650ea57edb8a88633d72d786c3fddfbb465f5baae0bb56e6e73a75aa4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h723748c756bfa6a0400a954bc9323e3df1edc6dbebc6133ea784f05439331dff1a54f3db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137e03b1e91d5fe53876d710179e83e6ea60933b3c9ce78597852288ef1ce72dcaf7c23fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1620af922e3ef6a46ec409e908ce64f87233f5dcb3dbbaab738738a0341b6da4c0d55c5a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1feaac199c0e73f90409b874663076e585526ec865b21a3de45a609187ed0554349cd0774;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d48b9cd7e12d00dedc9549784e06f070d5fd9ce5c8fc9f97be686d286357096f0e61998;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d0545cb7048d98860e365a74a7a63f063cc94a7d8e6b7c9851c18c872e66864756c0978;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfe6be575f5efa8eb052cf7f45a378aab82a4c59baac5433395590ceed9f67413eb204e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce61681bcaf3d53d4574775d2832000dd6e57114bcaa20ad34b9916456ebdeb0417dd7e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b8683ddeb7d28603406d1e8588ef2ae40c24795af9f31420055ebf259d0af2278a642c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1659def77b38dc0193b405522411cdc57be111d35b8211db1ce58afb8d7620bd78a1026;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h887bc5e2e49761274b50a1268286c882336c959fc7867b7a54e941975ac88e41ae0367bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc05ad122ef27f9e7d0b9530a6fd42b43640e179d92e8887239af79635262ffbd2efd38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94797f758fd2d64f94dd35918d0fdd5ef6e2b333adfe126195a62ae404bca470bcaac498;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he71cf23e5cdbb2e512643a3727aa19414ca2031a9a03abb5422c0d61c930cfe8cf7f4715;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc894eb979905d9cecc37b88ec92b8bf99dc81bd4170977da08da4da785473a224d4328b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77842be9e03474125b05a815df635fdf6930699b11c98cbb55e4035bd42a8eebbda9613f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ca795cd586ccb7da3879b975be349f68ab5326e38007655da922c1d7f3477fa56ef85b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42d2f6c9ae42cb0bd5b3ffb7d8474a5b5a441961b2ad9ed39cf7db56a60f666165b22ec8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fc45b778a39fe83be8196d45a8fca0788b679a33f9c58b147960515cd9263c43e954949;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5f4c24581d5fdd110888c3a17b7673206f2650080450e1f1cdbb25b7054f01bd9da4b3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ef82cc2877c0105ff4b90b534170f7f1259d19b86796472acafb13c2b9c26a374a8310d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d263d9df05a6cf0da9538e97089be656b8a54803933770e645f42f3c9d1bdf22ed52fc3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16accdef521e9ec29c36a33f99ee613661fba9247fbbc60ebf9e5ed34aab42ef4c114211e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd938b9e25ae38a05edf62a8a1221d3999d90506490241ca055c177aafd17a0f10a86539b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76fc413250306956d3313936822fdf05e8986b49c8b0d2331c9a1f485442e859420147dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127a2c440134e9a46934eedfa3c59c81957ccecbbbb428d7a810b6f945683b6e1dd7b3f72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca8557aaae22ea33ee50aefc1eb00617dfc2249918476d5ab30544427e321a487461bfc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170a02e9d72f4414297a046f529ee16903619d50f4403b7932cfe7972411f883161e83d8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100362ba6c1662c662b107d79b7befc95d1802f18dac9f0acb8d1e99a59ef7ee003a64811;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd63605a6e059ea61c7dfcec29ded8e8d2c7e188d83591bb607c1f44d0a4ec8a688ec4f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5468963e9c2fbe4c2b9d571ab17258e6bf9232f99d59f70ba5b2d8924a048da490c39ef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61aac0944114a8abb7a23be3eda3157eb9079b9bd5feddbeaa870018502f6a7dd036deab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101bf404d9bb79edb2574ba38bc5a5acc2c20f65f2a26867368d6c3d3b7af6a990dbd8f66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6666bed3bd55a50e240b09a3ee8a78c7a1b18a054e359a6713cd40787c1a22e8dbd17ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ac845dfa89144b3a021499f66d85c50801f44f53aa0e5505355d7bad5d719dcc2da1c30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a34d29faa779035f72bc5db04d167b21628d741464e67c205480725e225eb6a7a34c7600;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9db04cab111ddfcd5b402b99c84f3a9c028d0edbfdd3317be77ee2e5d0bc3dda823a15c1;
        #1
        $finish();
    end
endmodule
