module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [10:0] src12;
    reg [9:0] src13;
    reg [8:0] src14;
    reg [7:0] src15;
    reg [6:0] src16;
    reg [5:0] src17;
    reg [4:0] src18;
    reg [3:0] src19;
    reg [2:0] src20;
    reg [1:0] src21;
    reg [0:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3])<<19) + ((src20[0] + src20[1] + src20[2])<<20) + ((src21[0] + src21[1])<<21) + ((src22[0])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he849d6b323827431a28d4c9e3d710f689c11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d0610a04f5f8af5c2c3e03a205444549517;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5675693cd7361018274fd4989f837cdbe5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h676fe8accb58849b5706d7d7890202d20340;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6635f80f2b420b76ae609eda19e08c2fa26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ad277b1db6dd04c239a3b0b2795b1b830bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b82d9e9f486132a1694d9d343259ce43d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h814456e932b662ebc7192cb209696986090a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7193435dbfc578d71920dd079504d95d01a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3962c800c9de90604349019045b94a1eda74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc834eba2e186a72b6284e25835e011fa56f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f05ef5a151243040efb407c1c49b972ebf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27ea0fb358ebe2246d30553d1fddc6a1986;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heeafac8654ef70dfe44f9b810cfa50c137fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h696489b20abed4796c88f447929c2dcbc646;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd163971a1d0788d699bff153bb2e012393bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa4f1e67f0f73ddf10844774e02d0db904f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f9673caaaef80b294a50c55e06f43c55d6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9546ebb65e24a329e1f06943775204c2ab15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3e4b177647846c00f6e20cc89370f946eda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ee582bb5be7dacb0612f2e55517e2d378ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h403cd55d581550771038090e4e51a27ea85c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8756ec9e15181345a75cc04e3845bebc5701;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55994e2f8935a83abbc26a19464a2f3d694d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9589148cab12c6b26fdd71fcfe1fd44a12a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h210fd11f712690ba0d89feb1b0bb3728a83e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c9db69eeb4e211b081b420b747cbff8f476;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ef0529953bae1fc4c4529ffdf7686b021a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had64bd8ac9561aba4e1a20d360fbca1202c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5959df73d4888f07752b2d6a91fc8942676;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef1f63fa4c9c6c8e7376d105f54fd2759e0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd22750cfb07e39e376cc9bb86b20b7791dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2780e054f9b4b3b3d0a01880ec0c45d28f7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1635f504743ef62ab5c34b36227d20a9301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96cbb5febeb1be9f8c58882bbcb78797cf20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf8194de986898c95c38985f6402f9eb1b32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd96fcf958ccb0df268b7c37db186f15015ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1a05bf93dc7a71906c1adff6b1c68e4c0fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0edbdefd1cb9cc7cc2d606e6a1c0bdcc5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he50d9c3808e28ef4e1bb4b9f3263fb9f1297;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h478e3ff0090da5007e10528d69aa908f3af7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7103a79cee5283e8c6716734814fef99766f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdb95bcec91414734d2de250a8905a2cb20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5aff2b038f4b8de3203badf27da53e18905;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7f2adde105ce2338ee4cd028716c4d27779;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcded4b45ae4a36ddded2a41209e3571932c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5c8cde61b65060300e639878ae6df30e89e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64d1df27a7a1473a09bf185928a443f8c7dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h191e7cdfbfdaa2265b2cd039cb1676553502;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8020127527f2b46adc99c81fc8fa3687329;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5496492bc9c30a336b9891d8834c894bdd7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf56642987fec71e6a4b99f5ac566f76cd8f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d05b08c987a939bca095431dfa6bd6be68d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb24ade24bd01d643402ec3342004e0726ce1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha47d3a7cc59326bc5999f7e9885f40cd3a46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h580619b4deb2bb06e82e795094d09bd9ad9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12d2fb01b1209d69cc51ba7aa1cb0e66a8a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he422f7dbbb12bba8eb7a1d43b726bcd448d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf009490935bfe2fd927aa6eaf88e882ece3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h517bca8736352166a9a3ab73b7dd48939c6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c52440957eb982d9044b9e037b16cc4002a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff645e514077a2b671fbdfe028c65d572132;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37af73ab069ded8bb80747415f22d10d6d3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b24db168973374228c19bfcc2adbc4cebfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h654b783ec37c84be234d4c7e45cdeb9a0b6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c90271bfe9fd1917e1a6f9198f40c7a7f1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb55dfaccbd4c4029f8a65cfd96ada5bc21c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51b5ce0c7177eaab45b2e0fd0a8982bfb2f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca59cdfc174b02129311430cab088b823379;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef2131a77be1ef0de44058ff1a01917c444;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1743bd8d03634d149e08cc830a2d6e3d2bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h403d0e8b9f287c96f29650fff32b5a3bf4e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4a0911d25db5054b1264e46ed42318740f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e20516cff7810976f999f8b8a868e712575;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fea9c09430741711568509003ec060ec29e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76e395122a9919c554c97be6bd90beed4596;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee445cc9506f8b6115ec01f1d54752775191;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bd454786c92799acfa11b67df3749aab1fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf57d459c34ba6f4bc8f02fda188d1884ae81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd2707afebbfee4635abc763ec830c7d1b2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6eb7d535fc7ea6cf311e0fb04fd3d88b4203;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44ecd9e273264cfa9bf9c55260e10d31dbf1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5d1968d6caaf0eb5476ba976db84890656;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46fc8264f48c1a45b22047cef62dd40603b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dc3eaee537aa455b75666c089fea69354fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b1dbb46a607a11fa01ba8681a17c2f6035e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9f117a75e0ce325799d912deb5a11b34537;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3273909fc66ed7e0f0748308c13b2015cf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dcee3f5a0a39d60d8b44498f9b4f572b3ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86c547cbbd245412dcf881ea74b563c1b43e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdad95d818d8ec6693cb4df9ea2689363a948;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a09271f13fcb5cf72065cb277ef42a82e12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65a8f194d65ec41052263b2f925cc5fd4b54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7dd9fdc1abfaac9d2b3bb0da9c42d8b29b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h917ba29c880de2689002a8971f0f1b0c7e5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a818103117d6f0185916328e9bf3bd89ce8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd4e07d6f030df21149617b186060d5a8915;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h688794cfca8cf58352e626ec3076c8e85053;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32cd13b6dbd342677180dcca310af52aead0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a90530fe56e2bff794613ea8640b7d52d03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd32b9a148bc165bdda5232a7093969de6318;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6790c621a18ae1c9f77262169931dca5af93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51f9b6fd2694f43e11767025cfff58f7ece5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd05de4dbaa4f470cfd54873fa5ee21f7c68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cbcf23a1a043abc91bbc8b4ea5f97cee801;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b93d143421d90e2c42d467955b631f4b464;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cbeb534112d4dab3d3c7ef777b4a36101b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdff4156c1d878e4e720a8b553ecbbc8e66c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e3a17170446e4c94a48814c3641dd98061;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaa6bc74248ad7f97dc66b1619cfacba20bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4589e2eaf2f6123822a237cb1cff39ac65f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66d732e1e742abee518e603aba1d006f8468;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h778c27dda0d893fbb8ff23e0b454a9604527;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdf1e70a9dcb715883d55b98dae6d7b2195;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc2cb7b09e04ed333b50b57f9f78354e6b86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8e4ad58652872ca692b63d89692c11225ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11e90231210a05817db63a534288ecbe5b55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85299fec6df7b2ef4bec461f6911b60567c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd46bbfa098fbc2fe2f2f4bffe906ee58a97c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5883d3f64a91f83d8bbfba5cd19ce872a1c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h893a5b04e9484678a80672af7ddbfdb6c7e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0190f9658fa27592bebd886808e08efcdf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61625259e7cab22a6efc8c74b394db7db7a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11e990148f96a376ebc6d5d9863276016b4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e83ca365f5bd914cd11a3648a135251107a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb15c5f3b3a8101345bf1f65565343df74d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6869c3aa8cbe24a6fe3eb717ab31219d47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40ec903b77de81a9b63a0258c4f99c73782d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d9e3b0fe6bd6b0cab1243772328014d9c30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3745c4f213222bc0b70ac275d3c69712488c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h137ca5c7abad6fba6717f958ff72774dc602;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd95ec3a2f927d1a9074db40f57508765c6a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b4c2f0c50a5ad36218e569e341126075cd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h480dbdcc1014f84ab0a0105d6c1af0600a65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7d9e73eef729a9cab043dea2491b28bbbd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bd2d4743ae2ad30ead967645951ade247ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d4f064a857a5d6c72f9caff65d49bb28041;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h159b540acbfc0d35745b61779ab6b6929d9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41e93dbb08cf6146baf8138f7ea72dee47aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7bd622d3bfc0f0447b5bf69e459316a4d28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa7803f82979f893557dd2bf9177b7712c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39391ccf68d566357264cceba36428a5a2eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d9148e666d9e6a968ee84b7dcefce25b0c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a01c3aaba47d4bd64fe48ebf7e15417956a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85e35c95b50002564c6655dac3b917359141;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92a221f41708ee236f2b95854123ac01fbab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha69d2d04aacc1260a775334c0bb419771515;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2387bc532034b52e5a91fa05d3ae0047e35a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae733ff0d6946d39d709c95cbac6292fd192;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc91b158d7e49cc2fe1d331672aae090f9b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h495b4cbf6db5983273e5f51d9de920bb8784;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21a3aaf8e2c9a22451ce663e0e72a0839e0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d185197b7b3f8d3f1eea4f267a934e2fb50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3b6fccc480e5e5295f4c377c96ea5feae16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9ea2215964bde89d6efe4f0bedfd0133d45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb993c9ba72b627a27912a1fb40504ec0103;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b6ff5c0b07ebc755eb27bf40d18a47f4f60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1315d9253e324044409ed166cb4846a9c45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a36ee0b38733d0760cc3e848c2dfb433224;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d037d10cb04c2c02046239b9ccdb7873b69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h390e28d10d35bceb574d6b301d0f0b9c0972;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h549b2d8662dc99821b6e1d5642583767490c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ccc86fb9e1bb13e1e76467150242586fa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1750ab1deaee4d03073f610aefa91e30cd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha19743cdc20841fdc2650b56aa968e56071e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc929f97b9a6d5ae15989d621dcae0e84b9e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he238fd24a7189106446dd95890aafd229922;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f590df7bca96c6266c34fd1c192295a7ec3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2db88e110de06fc5cf4990db05db6deb7c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff744f27dd32184b525d914fa8ebc8a0c2d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0a31dd2dcfb0fce7c3b86c4effd5d7e347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc9386c1d57a932bc896c7455475ef814ade;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c2f5e11a00380b248e0e773034ac80e7730;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1ef7ac01162df62b2725f749fa4901c81ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b252405e0c6bd09c07e38b9992e956d8ebd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ae0dd091e4cf5ec092268ba109d1cc07ca5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc89bbe05dd8f42142f7c771d91ab70d19c54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h182a1bc05c087f1a0f62329bbe9b9e4e70e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7218fd9e4f554d5446723190723abedf0aed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3526989565cab173186b71035756827c7071;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8f920bd2b480c7658169b39b5c730f2defd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h532e9dad8f7980326cf91479b69462e57ad9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85a84ef43ed14921aaaa364bdf87d3ea4417;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61d1e45970b3d83fa14f86177d9ac95b0b9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a0f5dc32433781610aed63be97f1d1eeed7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf635cbb43c179c898f8659306dc9519436a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he63cde0f3630e64c4627d6b56167b175370;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe28e4f442b743669ebbcb3fe0c31ab604e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8928a29f388947c503330e0dc42a29f75db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bbc363f8380721e6e14059b3aa4242db4d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24e955b5da16d86e3b2754e3f887bfc6fe56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d62213f7ce0522f1989f1d169732bd22f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bacf36057bce03763e9752051684fe5994e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6190e7cd9efe4aa9ef098d001d9187b8eb01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58336e09f20d079649c02e2e6cb3764cce87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2a662209bf320043989abee1fe93c4f19fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1432b9abebc846419ef28b6e4b595a5ce9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c61b6ec66eccbc06ee9e33e8a073c4829d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41573912500790aad89b1e30fb5b7c6c0877;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbadf9e684b916771fc0781107805fae46a75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd234dcc87a1eff3ac9aa44f64f34e1acc35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2a330e9c633b445f3b6c240237fe91e3528;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb84e0e10a7438861a17ccd0d15e2e683b360;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd69ae4109612c515df4a6651b169c00146d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97ce8721bfbeed855924c1fbd8fd3eebdb10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc595398bf687f2c82776660cf2a77520236e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h324650b8d95b660dae8efa045b3c59d5b4ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e831f7fcf46f63a9c0064dd647cf0e507bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha184b08f2ed21350f5f5788f3fb8c77cf62a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e7a54794275ab69a249374dffb16f7815f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd36047fea747b06bea6f2d8c0013b71abd29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38457b584a62cb52184780238361ff1d5e8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3220199dfb2ee2c3085da08071441ac07302;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90efb99cb1e529222591a5051fea6b1b0a13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6125da1a90de471af8e930ddb6a2a59eae45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7069104ad2fb278ed7dcbd6123b027a68c2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1221847e7431f26559fada4d54385de0de9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5db7f4162dc1003355ed215641a7260c2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ee87e0b4b38999c03d1cd0376f7ae21eff8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1364bdcb187d21e4383e3758041d574cad1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5888837cc5cf3b33e853394cccfc71dbd41c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf40648cf83534f90efb10918222f0a33c462;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24f06b2ea5f834da6ba50c30af9d952ce8aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h172f14bc5ef617ee5396c439d187c54bef33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17c5bbc143dc43e2f3c3e2dc09d650f14c5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf9046d153dc9ffebf173a493775b0b4b9f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb3028a5c093da324b5f978af98074f3265f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5b310d6885fb0965846d0984f5d349f715b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2ccec30f7a570852a2afb657cd8f435fe10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34536d748bb972832781c25a84cdd75fc78c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9ee65cd5f0bd8d8c78839a2051ccf93870f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70ab96a1938c98c95030b620baa512d6e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h951bde8e1ce0a6faf679229572fcb4cf500d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2e03eb2cea6e875b27a5981db00e241663e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h926efc908004ba65b3f2ddc16b6d67cdc709;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h728e9cd978845bacd46c878ab6cfa31a550e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6ace1b4c5fd44d5730e4c2cd4288381da6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h692e94dd90a84d4aa872cfcd1d18e02afdcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd864ae0f0a8942873fa5c72742ec2757b929;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5d57594c7e9d96faf7c17ae4dbfbfe7e0a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4cbd20dd16e13524aa1fcd1d9b735662d48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h247a14bd812378b4543bd71974313046a4ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7d51f2bc54e60ebb477cc563bcec5081f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf063f1b30310c8439f74d6d9d3008c3469b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9585376e95d8b19068265abe3497f10aeca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf85239c64d984afb9b215a173f848f69c5fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d8f4929ebddc97fd3fa376f475d9970fffe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h479c446d5da800cccf8baff55bc93240c2c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7f6ccddfea2c9ccc4451455852653c235c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f715b15fa4740cbc2c0dcfdf20c5293fc35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd22dd44bba16aa94ce7c045eed0135cb123f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc83bb6ba17d5a9364a7f6a08bbe611c70dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73f3caa1735d6ef805e3fd8351446148738e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d4b65f193f4908ebdc0bfffeec674dc5027;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6296abed07784fb56b3f7c05fcccdbf3939f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75762e63a904cb9d0be0a193d9f3bf7dcf78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8b87630938f199613d75b69cdae8b99280d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4d72ee3362810d9c08ec0e8eee30809de7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdccb302843d6d985096ba733b3863c3c27d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e6bdcc3c60935adde42bf0be6a8ec8c84d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cbf3987fabb2eb8215ca1fca726449775fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35960b98955ac29c638a8d0b7996cbe79b11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cf111f23e82c4688356b2a91ff3b57ada55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb947794f6a48360c05de1926466364c47028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4a84f30844b1393cadb1fae6209cd821471;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9bafa2bb7d6056f07800e4906eb24921fe6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h213a5a53ae808e183a36e2e29abd394b0ec0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e21fd9f0dc58e4d999e75d2b5e9f28e1538;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd1501843fce16a433f2139933dfdc59a8d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd98680129da5b98662ac8ecc70a5cfe71ff2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a798a871adc2733207c98fbc082055485d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcc814df59244742cd75123646af952bfdd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57fd5a0895575fc3e8a464e9ff502bb5b29c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4340ac982ec10356e82f18570c09c7b8483f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8afbc542e87c0654c4d4d869c02de9c5552d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1432eee3649882b4c7860a21f0bfa748966;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3536159613b1b0a053db65140cfda47e9bb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa7bee785113f91d0fbb35afd255db8edd1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf6e481543c0ea65ab998ab1cc5a21cb28e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h804de10565440db07a5e023011fe20be3d71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ab584ce6cb5e11b152b3a8f3a6390a81fa4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd2f9e71eca93cffc91f1d50f85001d91162;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h631627dabe109c27e6f3909f2f473154f458;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd34330d549cdbafafa28a1ca5210f6704aaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdeee1c83e714005f74d4ba49034051a702f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95df36c1ffdd1bf33b3178ffd3cded628505;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff438533a2cafce6cbbace3253e5ccc82e06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa5c128006bbcdc6a9e718c1b4e143bde9e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5366f112c13859467316fef523e317cfa971;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd54a79c3dac608b9ea4020994ab63ac2e1b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecf913aab3cc0dd9bb319f9f092a79aab859;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20908080911fc91d46c5cdb9714e6ad95bdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h831887d34bdc17f7af9250770e483c6ba98c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5b6dc82685438528dd8417dff266cbe3cd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3857974be544edc38ecf6684de884621507;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he366cbad01da98fefabea4c70ebad4dc1216;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebc32a09e2184920e3bdb615d0adb3e90498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd72809f25ca6b8b8de8a63c1869ba5d5ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef03cb1f08e6dcd489faf58458712d5fee8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h749243390a1b1f7714b95eeddb6b64127d3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h682ea0d6bf00baa369f2af62d07e3c932c0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea6dca05fd1c98e1266022c9f9cd85e8e6b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h741c3c408e7bc392fd035424460bee2b0f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56aed63f36d94aa172772c340d0b504477fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f3c02515d43a4377007e888084104567e32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h785ca3092039ba46bf2518fda59cd7641cfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfab687184a0d973234e00a8cc589f8ed32b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h647d92d36f72bdfb9ff26b270aacce68140e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c9c3b8c75f06fc24631e6273334966dc031;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c4786198dda6d1198e4d35ff5bba41851eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6f91e85d09601e53ac121dddec267c1a183;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6ae42184255d602457bc4deef4da25a78f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f7823b946fd034b0069078cd67018b72099;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h889cb905ede2035c4ac63a18ef79246febda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cbf95591dd8ceb582f2b677b7b1d51f9770;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4074637c30b844b694c347a0b388bcdc3c2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d4edcbda115dd0886fadb52f0be601218c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d41335cfadbad154b4697305a8b46ff2b38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2efed82633faebdad720cc126fd3acb6163;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa0fee6e6abb107fc1113380ef2c7b3e169e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he88cb30f524af0c7ef3cb752779004dfe8fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1051fe5b54e95da50eb8ada3ce692e256fa4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1798ba3322c7886db042d8d13d51831b13ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd80699b32604cf495cb27b785ea427d553f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94ec5b690b990d04977a08417dd2ee447902;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22031e3fcb938f2cb65c3b19e9e368a8e95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3340e9c01b3869ae1c6d14b46a21aad969e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f5e068f36d92f50196a455bd5c59f0cf42f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30623bf2d6b29357fefab39af0bc531b7b46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6ae6b99690f22dd5ca651d724bf152e175c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7480f00416ca6e96421bf12a789bbd3c86e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ca42eb4dc70ead6deeea70b619d820a269c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa54f9bbcaea6bc6474bb21cb9cd325164bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e1b2de508288dd69183e7c96808618435f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d46179e4dbfa8987b73425c0bc6930ff580;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd3e9b07f5f5ade5ba5747493d033805487f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a6f752c16912d39db374dd399d766cd87a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ac324baad6c75430ac1f0d8abe1e0e9b5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f3573d777ea26c84ebb39b26978873778a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98af6638efe2a2d23a265878ca9b9fae4f03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30bc5a57a3398a5def8090fddeed1dbaf081;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4acfca5d3158a883b4230cb3fda67ac5e394;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h844ee6022748e3beb9b3b4f34459ba89d485;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ffe84bd4c2150d4954c3d59fc8c59bfcc9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ea5cda56f55d200b4657914c9f7e6131bcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3293790ebffaf24da7deaf82b52eb1836fe0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e1f4d326dda463bd5853038b24550601afc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd133828ff13b6c835eb820ca54a63914c09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa4dae19840b28ae0d0cdfc71802d66a3f79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cd047414d56c8e4c9da783f6acc2aa175cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34c63963428c1b0ce689537e3e6ae1ac54e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h478bad84dc20eda860b1386c8afcfc4b3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h764cbd3dd914097db269ce7bca924a1aedd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he19caf222b7fd977aa98fc60c7999d87cc3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f04b028b3087f403bcaab643a2c7f5af761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46458a3b2d8be19185c2337897ec4e4afb3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h963a352dcc7478ecf5222d26081cc7c008c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99fda91362eb077b37d29a0e2cc88ea93871;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h927e37a2a773ed344804097eec5daeb41aa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b9c1a812dbcc8bf8c8da56eb243e6b0ef6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea019087b911659db8f62a45d610466ca1d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2958fff839f8883c57d41ff9ffc0a07a781;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfac5c9f7e5f47c2521cea7ddcf41198af0ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50483e1dee1780d21c271d3e9b78a543df7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb6bcbb25ae109e1251687be91cb3f7a613a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3426b82bd2f025b3c6b6012475d878e02c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d2f9c169e4d55901c21a4cab8d0b03dbbf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bca836d1770dd87282ac9af08e0e8c9b6c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d6b5383a71d6e7b418235fa93885bce8039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16f5c927a7111051bb9f89069c6c0d5255c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd67aa484c35e4ff1cda34d4349468c0d36e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbd9c4fd06e99236e083b370c740d5f1ead2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7e661ab6a524f439ffb683cdf32c7b0b58f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb330e0d2904051af44d7acc1e79de9c78657;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfba0a37aad7c5584e390e4f088c4409ff19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had30d050c41f59d095d9e6ce9e0a86982ad9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4f2400b9e01e1b6881a2e004558602398a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ed99f90975f399e93ebbdeb707bf1380e3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38649421b050cbb144697d97decb75a2c7c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfa484155ae3e36d3fb4dfbe20adc7d715ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb377db0c8a3e1c8744001718c4b00cf6c5eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5602ec958985e88edc28918209eb485f54f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91804abf99487975ad2f5b924eaf0e9c00ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d0a66ed8a95e9864caf63fe63491c4e0a34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23fac8e13f19d93c761c50dd7f93002e83ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e9287a9381b02d922f0d373848faebf4a31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39630ac5dc1ea77716c6956f91f60b46f540;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfec61796d31b49d0dc28b18d43f45ea71061;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h481a69ba7adcdf7e739b885a7f08848a8141;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3df717a203d0932552c466c80007adf2b2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10a798cfb9ea1d090131e5ce76cd9aa07050;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf4c2b3364fa96cf424de62fcc8d8fecae35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52e6741b92fbd8d1129221be93b3b368255b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b413ddab43b4418c25a6010127ea6c25b05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56c1be1d801db3be32ad4091cf951a830d55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b7c9557ebf51fc573836907e2c9a2f09940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69200fa5058c738d106f856d6545aea9a3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54647fe3fac8e4c50115c46c82cdc23a4ecd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc874bffce05c55bddaad37b5050372076aff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0936dbbcee53cb283d8e4ab7d750964fb46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61d7d055e56532ff7052dc004f88649da456;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h427e7e45c69fb5ec775f592b5e56131e6f18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10331f35741d09098302c7cfad26f8430413;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45921fcc3ad8caa21efb521caf5d73a35cf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc66841d4c198db1fde2cff2633b2b31f753b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffec990e9a64f8e267a3f80871e5fc9889c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had972821642f09cb059aef645a17d63401b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h616750983e77f81ac7e2d84edf95ec468c5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h598658af9fffaeda6a6ed2d817d68eece0eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc1e5937eac5dbfec200f699c7dc3b182529;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b8580f8c8894394219795f42674a72a5b36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb65d60970d27a18f0973303e0ff42422d824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h359628d5f368c44c4242df70d8ab40f6d562;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5874ede8df4b88ec16e3c301ff61a15ca2d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26167cb2d48918f48d7b499cb35a3dd050d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92a77c045b5b79d71a470f96a7d663c018fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h284bda9908190596b9999ae668f2ac323ba5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2794f16de278f4e84b3145ebd0f94fe314aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fdefe997da5223754dc74ec6a4ebaa6bd14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96a4093e3f22625eb0e1ab6fbfd88d012401;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78165a9de297f61abd8d6171e2012289235e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4cfa70e61f82e486e4fe69977a5dcb95523;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf974df95e261e0e1263c94a4d1398918b882;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ff2864e0755e7860f7e8f6324356a505749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a130f4f3e1e955325eed1db9992f7f92c19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8366670081cec1ddc8800065b46af29b0e55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96686f6c158e790e95b81d531a2f10b8f005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4136d8f2f372545f9b9e0d1f518124624e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haed30ba7d5a9b414dcedec5d59180cf6c271;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48fd0a5318bf9794ac58aab761b59c1f6445;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e331269b21b977a165b8c8f3078dd8bf14b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27c590968fad2daa70339abbb04a20148c96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e5909936171a708009e7b3e2b2af750d83e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f54814371f2e2cced5849908c7ce2aa8c48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87cf3dfcdbe5aef3727e99ea0605c5f3eef1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8ff6e19f057981729e4e34cb7219ae7a085;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd4edd7ac4816c2aad661f58943ad5e10094;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95a1d158975cee93c591f1d01ad4741fb598;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a087f90d47fcb7003941a5112fd21381253;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habee74620d2a257042bf07850d83fb224394;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa883edc794e4a099f2a9ec08d3bbf35ef8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f4eb779dd0631d88a136d26d203834d4fa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd91ef99e2b844e4e8686fd79712d19f1f863;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb8e3a289e23899ab87a220c4168090be524;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc58550aaa459a67f56cfc38cc308042dc524;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74f5bf3e146bbc631c5eae79ebf4fef720b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2dcd9477faaa3d22612d914c05af89eef287;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h946ec2159e147c4496e113cf749a9516146e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cc69e83021488378e17fd18266793f3d2af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3b34c7dc7a95f4ed678135df25b039ba74b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3592d15a0abf90a6091597ed21cbd4a26a93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1397f04ce26197239276c4f1f16360f1f948;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ff10107290019786b6502e8e101bdb17138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0548c5e0261c4ea6e70270afba37f3129d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98729fe134643701678f9f8ad3d877c9e6aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82b4d5fd9be537ca52009a8aea5ba86edc95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h261935351dfa95f808d7a8760fed7aa6a9ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2ce52ebbb1d2799ba92ab4ada8c90ca845e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f0fbda66b9652992680a128db6f9ba2db88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4986aec5beab0a2acd2ef93708f28ac6e572;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec2bcccf5887c2a67a05b767faeedc5b6306;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c539d1c249c37dbe2035a23ce752f2ce371;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h577ce97153f5dfadb22777e628f88160ca08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4e4ce0039dacd1c28c82763f0b6aaa041a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf00157a12af74da288f5f21bd5ae98d7287e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c141b97ccd56145f96d5cf82798743373e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ce0214e9af763cd81fdcc9924beef6aa859;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43dffc1ebc53ce79fde4bcabcf6faf48d438;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9990b00e77cf6b498e1deb0a937fd1006e2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b2e2a83d1fea4bebf13f99caef56543339a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h986a3e5430e0a05de54b5ee9805faa6bb9d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0a73501bb17e08069bc1828302dbf00c979;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72df7b9a2780ad2e7c54da42bac07e86cc94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7406c60529c71e8f90b0ca89a50048c876b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h415b370dd90bc94f81968a7a3931156e8aa3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3a3d5e12d62a4187a8cf72601cf2b9e622a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa12b8f132f88b64ba4587347304e10ba12d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8eee67694f8492e71a42730615edf2861c39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18b4184c63d4a9f5fae157daa28e1a1308bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b87163537489216558b2920a6d73858bab4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89b30c1bf9d08f418bd542cfaacb259030a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfa3eecb2576622b5aafa96cebe63bd5a8d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef383e59f2e3fb2d458f75d0866abed32bd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h360b566c837fd15eb19889a156e40a02b024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9367b7c74292286b8ab0bfdb6a30ffccbc2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h736895838540dd3c4a8a49277ae4be73e7f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f57c6a0ccb7acd0a6a6da0bd37d7f91f389;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0c33b6009e3fcbb774b3f824f4c23818440;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6e73ed2f89f4487344425f20fa0322b50ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb95b25f985febdc7ad8c1522ac32182659d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65614aa0fd421909e4ef32b84510cb9fcb9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb613c0950cacac7c3faf19184abe4f5e4fbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7ba89e513d2b3901e0fee4403953b317178;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8edd4c6c5dd2508741c905d63b8f0dca1fa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h223523be9f72f706846d8c17f26f8b5000e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a9f78806a05cc2edd4633da10246f1ad4d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ccb321613803a94cf7b00396a39afa04376;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6942248523cf2ac149b05f51007cb0a287bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19afae278f6f211bf9424078723195455a8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83ab03fac58154a9cd3212ef0fe6b9b23f12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he93284b75b5ed2c79b8f1577cd04a9440b3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fbfbf6852ad2dbf5e77d7cce226af10670b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f11a79350ea550a207620c4088b635be92e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h594f46d58604bae9e11b0fda4f623038de30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7eb2bf1ff13e73974e5f3ac8072b522786b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6373e9b4ecc116543053bb14918ec80d45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0375bdc1bb521b8ced8b6a32bb4d6b5968f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h838ab4d1b038716fea93abfe1fc719ad617a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0a334c9d383edd813e6a3fb8fb608739c15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he810fc5f9809e95c9136e465a86d68c2e4c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdde085007a388a2d9fbee24e650d58111f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6b1ed603b2c5657e02a0f86f349a92b8664;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc2307c63d95a27733114db672611c5f09dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ce4614ddf8092a3afbb268a55e8ea80423f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73ca5888a519da571dbedcdab42afb581cfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4167f445468fe385fdf7f02301077bd7e2ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha22930074f356cd4f66b9af78cd168f25a27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he47517d0350c5f4c602017ba37b68079c9c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3685812aa69298d71ca6bd41040bc1458b5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3aaf0bebf61b5d0d2dd925bc7664154a0d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fee8f447a6a084f15e00d9d320248dc1f9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a3cd07e107328471d8dcd8099877578b52c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15a762cecea8369e42cf5e272a281e2d61b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0459d881149ff21b08ecafa58c58c4fa345;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafc6e95459b5e32193b7f403c17ad017fa15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55abae8613521c0cf1e0eb1f149d9638f841;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37a5b8d138b4ce16442ea77390c524c380fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h101b1a11c6f0546c061df786850ee77a99e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20375f77670e75eeccd02b056f416e7f3b62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc10168521c66d60d7cda9691fbe6721b486d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h640d5f5206445ecfa0f567a2fb9bc54625e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h881fb480291fb4400f7a56928b939729d53c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf45bd8553a5fda17ab0a5fde2ba2ede21940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b429208ab3b0a89beb3a48effebbf4455a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32c80e69afbff821099bd30092b9bc7f4e90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27fa86a417c2b012375f68ccaa4eacb670f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81022766c33b3400de9bd0396897e2ba3792;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6eca9b5627bd40bc13a24ef674f575b4f25c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9364cd32899025da37abc06907ef7623bcb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h382ac5c30376cbe6cdadeeca70e7b028899f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c89df13a4e67f6ae02cf1f5a1b7b5dca425;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8a8d381af9a8e775b9a570d9e20eb8c5ec9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf12589f8fb96225a15ca25824d7e26f28159;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bcdd0948bb34bfeab5b5aa8a42e118eabdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5709fc83fedc13ef3c6f5689e6486ca83fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h400d39ea5d8b044aef623a9c921124a973f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cce3427a80f55c11eb5a058a06346879a27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d2f206b6d8be3240e636f0d9bb05f96c648;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4bc21fa3bd7dd64a75bc229002b9fdff49b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc3569400ab6fa04dd8070c6eaa3ba5e85ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4db881bbd05fece4a8e5b42e24f13f06bdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h294121ecd30c30bd4c8117bba8245886560c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98692ab929d343d81a2589ac15fa2ed872b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha15e7aa4f6df01494b7d8a2bc29be9160a55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b95c031efe080fc64cf217fed6dbb580efc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb65020929ca032d77fad40d7007e5679b6bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dd8f2bbee78732d9cf51847fe5a00f5964f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1d8c26231955a72d179fd03d7264afc113d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h668fc401fa3e60ea4fdc3e393ed71b90497b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f49144e9c5ae19c034b704501522fc59ed8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e38475e4000b78fc0c9362440e1e922b73e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97767ee38e98c70b0284fb705df0aae03063;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13893ce3212085a41cc9b1b70ae9321267cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd27eb916f9521af75b93c655af7ce686e7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcc227ca6bfd26cee214a2483a4aadf7a0f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3783b1e09a939e3d71dbd7744d1be4e739c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e6881150902088ea9dc0a892f2115e5a547;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8a97ab506e72ec1a4ffb6170a687d61d2f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8716b0ece9ed2a402b2d69c712ad31ea28bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6454995e5ef70fcbe6da1f8504382ca65bbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46672395c85ee8e76f23b57674845def8b3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85e2b5f8e63a1b2b3f8ad9df12fef2805723;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefff1ca86254c712c311a52c86d2a4b7ff85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h361a55ce9bec01e4fbde7e625c16feb8aa9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc3e07c312ba76a27fcb8d6bcec92c45968b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h755c98ed0322d453bf43ab9219b5b610aa07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f89ed72785348f2a5d2a4f9e916f10845e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe8c94cc142136973a3833364b7e300c79de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d91539be7b56d06dcb94972d37c977707ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6e7915b76244ebac866a1bc521c7a1a5e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22d460f9e794b72c9d9be657d3200ed506b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dc3472bae25945a7c577de764608b4dbb03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86d141e455bfe86ebf9c8f9e86d9cc8743ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5126ec0e283fb6a5e4d67b9afd665e7de633;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h683b41c1cb6258b19c8f7229cb083ebbb056;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc04f33229f8944ff97dea847185abde81e4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4099a31e7b02c468b2ec35d8e57c4c526d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77b4dbe1ffb353c62a0cd459fbe0bc602da2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cf12a5b00085356309617d68ea86f5aabe3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbea8b3c552f74e60ea2abae4cea7d31a657a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5da4be7b2e3028913f4363178a32fcbedac5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46b95d90bfbde4bc674ddfdc1065aabc6a80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd364a160e4d63863ca1222ba7721b2487e8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fa0b85a69ea99079fa2a0db1a935b8e8b7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h169fc494076290be0a7007c5bf8e3c5c9ff6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21518a20d7af4aed1510b6c66177d7e71fa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e075cb0a6d8e299a4de382f4e009b9eb6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d8b45c4a76a4c790ba15a3e4c121c91fd34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h326c288d045c172ed6c164654c2b1b95a704;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bc4f6a8b5d091fb1189d25c5de5fbc3feca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff20877b7f0aadaddc95be7b8f65ab1ad05d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e408f1c80d8444d86de97bd28d502289af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73b782e762a74090358fe507ebc44795517f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64613ea5b82e93dff06e64a10400929bc88b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60acc45ec7fb3904f3d7a44477b5c3eb54b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8743659d75847e12cec244d78f05daf2b268;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef6055422a9d49308f047bd5cb815a41441f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c823e6f1d226647e157b09493f033561b7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9da4a3377174df9637a73aa53a39eea06dd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf13cb7c435de9ee2981c821e11d6cf9a575b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cc202573ac65c034856bd87c5295b1ec89c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha04800905114dac5f905995611af61d75e07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba2f23271256428675e5d681f046b279628b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h393a0881f52dbfb75ca053fb4e3b4ddcb972;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacee9d94d9b9d4d8f10868dc8d96d8db6b06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2466d3222e52a60e8264950852e1f92f13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc77833d787802374193961a187977e3acd78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he92c39ecf63241b92d4c6e985692bb5f6bbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d654f9eba40b8fa472f07cf383c609e2fe3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1828d7c73941b314ab96a70e8002d5fb10d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f70cee2042ad46340188acb3b59f14aa8ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e14693abaeac1d6cd7c3e5a5a780b9df6c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha81e9d9b36ad337ae5a61beb036ee4d1f60a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35422954142b248cf80ddd26b995c7f12c77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf13f58f87d5d3f14b8311095dd38c4dc2ccc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h654e8998c791e3646bfd6089ab478ed206c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h265826a55d1e5e8d338116b2c80a35682eb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6760115da57aa08840d56899d756144628f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bfceaee0e3c06f60cc89d2f87df7bdf3337;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99ec1876ef4495bd3820827756e7c3c216d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fca3a84700ba7b558e32c3d27e591f6ab9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h282bc22e01e9bc42209ec956cc5b3060997c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8eb78b347e8a5761f726f233412e19b0950;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7709b83ec86d25beeb650ea0b1ee37b2133;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39f5a35f65bb28103f1d9ab904367f3870f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h369fcceebaaca01cd7efbdc0ab29631c20d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd823c7bd5521289e9cf25a3db314602b35e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82429d2c5b5dc0a7cb547ff57201f1d592b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h452e785de42bf73918a7139fdc8841b34113;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6df437c83c096a279c8ba8a5cdc0feb2261;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heda63b5791e89748c9814e537eb41b19aef9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3405c22155c0b0b70b0f3953d7a683115d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6f7c20c1459430cc2118a7e73f4d4a24ec7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had212c6a67aa8b91b4918a60af18193e3c56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc944f60180bdfc9b270e4158c5e5f8ddffdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56e873ddfc5a4955605c14004a6e46118c79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffe6815691c3ea23b59e0cbd217f3f11acd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h186b3237d943cf5e0bc327c07bab4b5fa1f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6254ead93bde9cf5e91567b6ebf8dcbc174c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76fe6883b86863d8e442543f935f37c1ed63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h410988dbf71af80f81ce8aafdb3e0ee50818;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf85eee2e8e333cb2916e6c6d3c842c8c7d17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31b21678b911749d7696a3bb7f008399018f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a769dc8b18531a476e670452564df909b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76fb051e9357ac2f2c5cfd451af2b07b2db0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he50674ed9e86ea294e146011fe5a36778c79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he07485de260a7c119ce8e317d99ac5fac5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82f3395603c45374ca911ade66d92152c187;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c1d3c782020da5f9961354be9b35e4d7d2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h121f5488b17745c046c091649e97ccf553ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb5c65399931ea976d81f22a401c3b9ba01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdefb554917b17b525a36145793392f225a9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefed19197273ebbe055bc284912519b9c717;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40e96d3a38513840c4e1003f1ced56d99b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b5401fd1651575c59d3e50629802ce71226;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h426ced3e3313f947f9bd8c2e93c810077a62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79bb91eafb0f94c7abee8349f1855f527f10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5f22a1bacbdf71fae6ed46b845dc786a6e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf8ee1f8a0f8b7eb9bd56cd384349b6cfb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48db61c31855e71f4fddd0daa528c7d26e6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29c6d1c1dedd18807bf66b0fb07db60f533a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h413f6928f0e720ce133e6278b896473ff53b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7176e2692c1997b9ea6c908ccc772a7c5439;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h289c48f69345f2a3b768801e3be21e94c86a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2277ab0b777a08497acbc12bc5f314de8686;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc5d006045f54227845d5843dea406548cc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfe3118d219cf0ee60eb362f4b8915768a6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6182b0c64d9d5874091f5c9c208e436a2774;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h359c5faf78c4ef0866008f2f9064bdf707f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h985b5f704e2975d1c09bdc3e219570178d4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77e7e42687e70c30904c55d94517495546ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf09712b54bea657b537e3929ffa7f7fe881c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9923ea6ebae4028a7075f4e1c681ef3e1a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4208b11c9092efd38191c183fd6cc2463066;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87b2a24c8428cb218dfbca108d08be91ba00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h469947fa8fc17cde73d92490a87fb9761da9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ea8769bf03046b72443516f91afb725ec27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1f907656e9c09f5c2574f384eb3db0fe04d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a439db13485402265a9070a197dc38bba67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21b5edecb811f11e5046384baf88faab8609;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85c30522b3a1438ec9c2e737facb684dbcfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8bed8517849885e17e331d9484b37d0dec1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h624b5d72db63840a962974db0ad59dff6a4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbf0aef84e5be34bdf6099576df1e8e8ef37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ed63283c1f57bfe7a7c41e9db47b24c3959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b4f0edcf2d57135adbdea401cf173135ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b81a6c79e81e5257a343513e3d231e6c39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccf006aa82f81d1ec36ae3d627ada02583ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e30a931b9f8251a9d0508b94b4b4affc5f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h794f3d9f6b7aea9e542dc3d9a47bbbb43f4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h571c7163e7745ddc90f29eae1a5aa61b18d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71418cb28e203a76c03138bd5969611893e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7afeb7b801bf056fe93cad3d98f19bd1df5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf647623744fdda8a942e02dcb465479e4462;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4dfcd4eaa2a39736af69a577ad36647e233;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f62fdcb2fb65e247b979c0568bac61557b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h300d43033ee389edd408d6063f4b37d28b3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf24b5991d671d701b35847cb0326c80f3fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ae136b8e99e7206bc77e5c31397413d2e57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86f14c696ba53738c5a95e81bcbaa9c4e2d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7642614194e99a9286e585f8ee331d848dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfa30fda5c8c310f870826ac37921511a40d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc089abff4b39f7773f8175d671c068ff3df3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd542a0b92e83db9b42e6c50707580b1c2de4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74b1f2897fd55e74a0b1662809c6059097de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3021ef1a71157506aad071c6b8465fc96e0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3b8ccce48b4085068d4a8ef2dadb6103a4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had5f7b0dea8e764569cd5dc58f0c6a15952f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde72245db44e9890ecaa395ae9abb7387386;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h906ec650ce09f696ed48a8d79724c0ef64a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadaaf349d24427a8da9802ab8dcf5570e3ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63fe4f762379afa952a7da1c9494ab47c01e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ee0cf11f8f4fc5f8e41ece965e73f81f4a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcc7d7f91f93bd0ecc4a1cf951e1dd537145;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73c652baa55d449ce91aa4fbe85a2ffbbc03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8be93903ab3a724a05a22eb6fe41cc3710f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc5eb6dc2b97012873782e3185c361458c21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h446bf278e707fba42f71774683fcd531766c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32eb13e0d3c57ad878915c9e8646b623cdf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87c3c231955335d9c16660e61420a79ba739;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93e71ef98ca03e7ee2800dfefbc9ff603901;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29d09809df7feff29560618a82476ef29232;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e8fb6dda151d8427b8473ec7982c700e8bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf80c31d8ea9e04ee4998d66c1a252716b4d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6b9459dd9ef157c7c23b1f00f354f39cfd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4c2466cb37ef22bbf392c3b9cff3eb02cc2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5ae4d82754b8f5d22d62b8a85d7c4074b14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd04d1a4d17149cfeafdcc2b7253f7b939ac7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85203a0e6843c28824350545f1d5fa8da058;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdc8ebf145a5ab451c1256da8eabed375306;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2849f8bc4b4457759b23ce358fad6f217b5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebf2ea634ec8e0b90dbb7de7ba2d429aad78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea94df286b7ec0560e596efcd62d85d52dd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79aa33d3ef77e4b0094a2bf643bad684e8e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h195ae8b0c4daf68bc5ebdb204182b024a877;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ae23a627a7c26eebf0e730169e90ac1394c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e4b1447853b8ce271abc6ed08742ec08c6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31ac1ff7b683651b1b9e2e8500b35f49b27f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b99c47a2f016bcbacc0624c36ec9e00989;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h546059231e8b9ad2590966526747152c6562;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h828af5207c25466824709f51ced723a3cacd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdafa8988b3657419d68f0238debaa6026336;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb54009cfd2103dffcc2abfa003026ff3e1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd6b77281b9e82b644b4c4dbab114916ce1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83c31495ea39e451ee17cb70f43b20b187a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89d8f89b385368ab320a7d7c628881471b63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha05e6362347acecf1dfb1c3676b4fc8fd4e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc424997677fde96fde140feb5b5d66c2762;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a41819d6cf4f34b52493212784c158f70a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc56884569fdd1ca6064d4b4eb4c1a1774f7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e3d72efab137cebadf2dcfa31fc9c74e1f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2d514becedabe4cbbf07b6179b317fa1073;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a24b36870ecca9893e2aeac967b8fce3098;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5409e7c36e114ca13a884e81e1655fdef3b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d3010be59d92e2e0b49a96deece0605efc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17f68fe3ac0ebe9a1a78d68e4ffe3d30a11e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h274206474d8802bc9d917ce3f55f35f24c6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20ea56c9ba4ab96284c42b5928bc5492b344;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5362c35fb3218dd77364b86a9728cf043e03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb53bdae20ade41371e07b2196727ce8ff70a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6705570f233722e2de38292ba10fafe94fd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1793c485fb07c9d92f8cdb07794ff516193;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fd8260632ed5ec4697076f0507991dd568b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4cd70608bcfa50f8e0dd5b44af3eeb7d998;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8230d64fbc5571a7e443ac7dcce5f41a0a64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8500a769e3307a0d53ff51363889e58ba76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f61b263b5698d5ce8618f638d1ad229e4ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b41164a1bacb166cbd7c0089aa1bb943718;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd628e49fc68a8d1770cb782d0ec8b8ff9a81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc51556a8eab061190028a8314ac17cfb862a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d0d68b0f5b0732c46aff1af7862573e024f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3da77d11cba58b6c9ad4ad803f9a31344124;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60817bb3ee255add0bfcece90b37a433393f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b2a6083ee37e862778278c067756ffe900e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a0a95a28cca3bd80b3058ee24d23028442b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc88a7c4b7528468663daeb72f17490bf73d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7564148bd69cbcfb57036c6570a49b9b91e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12b37ab71360cab9c08ea45ed82281c96a88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbf3c79f48cb6af699278db8294b940f77b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80ea2b19ac43d6b0030bfb02f45df723c727;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ba8c9c1c1260c3854cf11ac44d87fb73cda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8077aa6bd2f2a1ef0d72b97c5100f36a6a10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha794cb8c408ea071d8b8baad5a162f18cdfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha95b0df7bda95446dee0f8fa03d69cd17474;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h746395544070745c07acffecff155c8d76dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fbcce5b10fad144ec302ed5a665343af3bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h407779399cd9313e9b64e4e41c7f15834a78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30cad130ef32f6ce43772a0e4157db0a2b06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3641fcdba38848fd64d84b850802f368c7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5239e0118f96deed21aeafc79009e1ffa414;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haeed17d415f48b9e3ef090545eb1beed46ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6867a1e46cdd10e636833bcccac351711508;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2ecb0e1bdb49644e4776b1b4cb01c9685bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89506dd464b733e96214fd3bb9c06e3441c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had48ac1c0ffa4eba5930e2d150466102a0e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fecab3835272c169bea629433919eb91ebe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20d352f6d4517b20328102b2253ea181d8f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6572a752e1f7706825c1553f71296c5feff1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h739a456ddd14dbaae8f3c68b29bb34214935;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha61efb4e7aa98ff3ce29351c9e8b78f9c79f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a7981e4f792093d5c5be6ffdfcf6cad63fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e56e48359086a5bb9b9ee6f26bd5054e09e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20539ff95262eee748851abf77345f7aa961;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e7d7e096019e22bc072e88f46c39a350966;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h514e62c2e79ad554bb958f9a2d3623bbf170;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h945badd95d2b3a4be9f80de553b2cf7c1609;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5812c203ed7534cc1cea5b41f02c3e21c3c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he693edf87f9a0ec70fb5cd5592a1b4cb2f53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd168d1d33efad8602a98b737fd5a692f141;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf39e536b05e3341136ad9e2e7b6f3ae10988;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c9226410dd539ea8832ba292ca07cfef67b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6e5424b1c4ed2d55289e2f100abd78e88c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe5a8aeea9785839773cf53e86aebcfadb99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h626b7887b6767f6b6319f549b8c3d261edc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0c3c527a0bd112b15d8d7a2fadde88654e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aad5ba34ca9803286474298e651e3d43539;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h364acb6bc47729ea1e79971d6749e855245e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaf3dcf52aeae70c04283e788361a66a66a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf80536e30c484d91b7bdbc6db3472581291;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1ef2bb228ce00074983d2097e4e512a39c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c5a5eaa78302f857c6b467b05effa57472;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce70903da61435b56faee9741bac934252b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90a891cfa7dc4c29ce486706a829df42366d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62e75fdacd9d4bb14dc44212ab56da470a89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9af823baab66ea397951ed8b68cbc4686f57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8159c1c98f7aa1b568302f7af069c7970818;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e3f57519f7a72f655b33c0075ad740be68b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h900513dbda19f437aef59ae5895efed2e70d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4573d6b619d113e6f83bd276ddb04986b03f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc495ba3a2ce6d52f896d1434e96f69cc22c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53a724b7341aec7aadcb7b4d175900b42ba9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h535820fe018d12e2cf9c87457616c160a378;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ab75e400d9e907b34f7c6eec0a2ea5725ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f3ef9295cff4bff1b09892233c66d3fea65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1282e83fe55880e58316b419024f754dc11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf3d0f46f07b545ac71e39026d60f8b42766;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63367b8656460700bdf738ae93e2f21d508d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9281a2f7dd2ca3eea1090f7407d7922ca7f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14d0a31761544c7ec7a28e48c7d6b39c1a55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h732ca33a2802faee1a57a1fcffa5b4086ed5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2ee6a7804e1168e0ec8f9a53df390bbaedb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf229371ee3e911efa68bf9849fb617246360;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he079aca13b27869ada1345a9e7c2b2458725;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd81c30a6afcdd93c9cddf5d433972924e964;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcba440d7e54c6923e24254d0afb92092d3d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h389237b82fd5144168486547172bbda50dd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h303a7f449b8473f82d915b99e1a0220bc9d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcab9de5f4223151e244028d43659509a7005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c46f52abe33403a1cc43dbb7829a7e70160;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12d87a0b042331ac03083da52cde6fbe1dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7259a136ac77b0978f947e72735c5459024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11162efa482872b6e69fc502881139a7aefa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7b4abba1a99998109d2aaa171be56b46eeb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfe2e7fa250c8787ee1f7f873998b5833156;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98f7ae570900f32585eb53c4539617bf6366;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e000a80f616736d4ae16d870ebc834c29ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6e71d690de1af6133acaca41407ca3624a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7b9358c8a56e9b4172be81a6ad7bbb332be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bdb479e478814c249b189b5be792449ad50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h464207269ddfdfd7ae3de72428634cd8a84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e3ac1424abfc87b0f12c2696b4a060c6f40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ef6c0485386a0618bef8718ef26c24b4f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6f61158374d9fe22b9f30ac7fd515669df2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0ec8526619d35088c51da0aefc9598ca8be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2efd8d80dab1f82ccb07fa314369deca17ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4f243d4b3f0009944e1ac0d9444150d27d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha05cc65412fda3184e4f98a3cf5f943ed191;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31c3fab3514bba17b98e25d17add97370571;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50fe19dd4363e82162f005c3ab33bf19188;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb3248293f04a55c2e56015813df8d81fe26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d6fd054d930ad77c4fbdc0f572ffe73159d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec888872cf8b09d7641727b9db34f04e057b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd91eb229f552c5aaa7664034e466a3f9ac76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ceb5c2b80f4c96ab59b40c3d7a789ef7597;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf46b6adb32582d00cb23c7b0ec76865a1bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5f0f07690aaadf70fd8b0b2b8b1e8d444d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57d562bfbe1c32c5b5121029dd1c8c5c1f7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee8914474d4eeec977e5c11d70f7f91b850b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90abf097973e84217b5f66ccb27c64504ba6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h434554529b809c43841580e28c3d599f25dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h115a8a5cd0e95692f6309117d46325402415;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd11c1517ef49f4db57d63ac790b9757d8484;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc59200521abd1eb79ddf727f1062eda238a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0949cc161d49fe8c554c6254dbf1b9cb34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86cb56d5b7304cb28b58a68b2034da8cd7d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h340caaad798842c9e48a55616809ba923f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8190957332512c113176c1c7f352a879b8a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aecf9242695183f40f4ed84f61507a7a77e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd174ac9b6f7785841f4779341adcad9d8ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h379cf39ab4f2736cdf858b8dd3a0621b1266;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf115f2e8c1926a0ec5fc2fc2e53f1f24af1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53289fd881ee1b806a3f8ccd16e1033aa753;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbadadbc2ee3ea6f83f48b66493e83907c52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14f6d0ba97e898c721b79f36f3d0bb8056c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb35e4b05b3903038521992718bb3fb0ef03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ffc595813a8cf39306197aa2188ef4b4d70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h759dce09fbc748185efd63018cc7c1a2269;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h656ef4c25ac252d62fc7381ea1d5f392e5ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h711a1ce87157e16098bf6d7a692a5fb3c846;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a8a482be4fc3cdcc5d28ddcedb15e7fff43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2502e991c6c0b373f8f9a2af3738b31d51d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32a1142e7b09ef9d60a08b793fa44775fef9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he33751ec036a2bd7d641524db400847ebcb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h878eff828b7b790c20bdf5975909426e2f77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d152eb31cf571bafb3d8d1a2c78c5e55842;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13080bb5960cd5f2f8e72bdae01ceda2a91b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e7b7065dd4895621de7cb22a975724704c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77c38808da5ca461030b316688d013adfd06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfcf97d844b9f48b154a8439808092109bea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a12ada5ac5ccb254aec3470e01e89759cac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h639592a6892120bff80c41701101b1f43c51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8165eed56674b52bd0e88495c5113606cdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed66858075cc14f7618c95ece5f294259bf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7f375d3315f34af4b5ced883508dd6d9d33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8238b0e0c4f14c94f7deba062b54fcb9c682;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb8f0ba764abec6e2ccbea071e1902b7ab38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57d2aabc43dfdb2a551c94eecfffc2205523;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd4aa5e5ea8c03e98e2074fa5f76d7e48f79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3fb4f6c58a0ea684ecf8deaaee4cf61b61e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ef21e9b6206310acd24c09230626c76577a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdf491e73a4e1894892b078453e3aa6b8f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcea57220915875d64dbb8af4e7e871593bf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h288481e77be6e32615f16c410142357eef7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6dd9a3c34f6f5d2f815a4c0d3957b6b0223;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a59b20579de28ab5e13842954b6b58baf1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he058aa54ad07b65ffd602005ad49c924fa47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d03a46f7664340273c8ce89f772740fd531;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2490b9bd4b506481e3e35695a9b5302528c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdab4a2f29bb85c0072a05eac72e9113f086a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fb4ac0db24b0799d4fdbfe56a0c9a1e5e9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24da99bc228d3bc8f22ff112a9f31d52d8af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29ca5763e88e520588dcc4a6555ac439dc1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19a6f763cd16c1636519f8d36b2c57f03f37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4829559f33166a93c02a16482fb180b63542;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b2c65b4b5d33cec44d817e7b6936a7a102b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcee3721fb0320ed4408fc210ecb34410d51c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3e2b71a8c558094e628715c254aae4faca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heaa678e416e68837cac9109cf18db5999b05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2b6b631a5f2427b4f2622d0d13c7ec7a82f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58981f481a62285e99717ba8f0887be8efaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd00ef92fa0f077e6fcd1d28c83352c2d78e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf22005ea9c13b14d45d2f44f7e5f315d3b60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h320fc0b0fba18212b7f3612adc97755d4cac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa48c2d82aff1a67ee187308525b3d10ba55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8dfa025f7c0f2b80bc0d4b196b41c646a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc86882893898db086dfa7d1d3b98d0aaa62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc4ed7ae968d6122ce05dcfff17f8226ffe9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd5a6c69338e7540bed510031c26fdf024b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h298eee1efb78d31df9087715fe5973b66e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae893057c0cc934dee6e31af12e280f92b04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e2879d4ab10ab57c972795fb2e78aad6ba8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ef097ec407ccdd687a4a7ef32bb8747f58b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8257e8512f3fe76bb019a6b277196d69cec3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f0987a30c76c5228c8e9f29b84f428922f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5624ecc541c98efa8399c214d6891a51ccb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c5c3de13236dc60807319f2d2433ee0f2ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64563e7c595cc11d3b27afe20ad6ed3f93f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee3482332abcd0c7e5b6932b3704de2d1f34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46fbad2e8467359d663c52375c7ff35813c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3eace73542c90714fd6128a7e4e3ecadbbbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfb5c7e8ebc517f05f0b1382a50adf15bd71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebeca5c9858ab40a4e24cede2056b8bd789f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf58892f93f73667e6e96b6b621b9dd0c33d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a63865d74726fa4a925a21bf58bd5436814;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39a0117e7c8d2b9bdcb0d2e0223195e68f92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8545a9e1237db85e9b8902b12a95aa3ebe74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88e6d8a90c3490b5ef0860042b26b9bec5d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h243b89601f78ef19d3c3bdaa5de44dc40c7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d2d5687ea04d596e6b39ef1fd7b30ccf3e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8536406848c542533aaf29dee2abd411e1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h350fe94d718987b8de59c419fedb97526e40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50137265044e1f98129c874da588b68305a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94e1f8a30d8d3c980d06af2f2faca0552c14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd116db1132b6e69e7657a7e3af1478519116;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9beffce77db3630df531d66cfc66459500cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83d7fdf980817e8a4769bb7d38cf1aa81aea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1570d309f063b11f9f0371b8fae9a1e814b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6fda582725bca7a5c7243104d3fb64edd5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h859a57a3de35ed775805b6d1cb8282d17417;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb005726c415a7fc059e68c359b1a60589909;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94f9f1234a7f2a967a086573d7e9892c9480;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff5615734c8525117b04565f3f45df81604a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80bcf4519bc34d5b198fa1d6a63c7d6f5347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11979b7e5431c948ad95e5d740d75107d5b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf55c55ceba15c60ee8b5f8ed75b9916a0c04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb48a538129ad851aad4644f62bb93a1e427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a683eff060b8a8cec5380d42e53dafb7684;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b74f0fa47c90754d15a378e8939aaaf1356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63a1a8204c4a757cc6bef7d11dd308a3dccc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9a7cfb430cf4bf58b8bb8c9eaf5bb8e9945;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha45c8a93a48972c243086a209ba0a575c86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfd3e8ce9e7f48560187486cf3a95600dd8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h488aad4a64eb74096e7dbbaa7d26ea41b1c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c5c7e4416674c9d3e9864e1e2586e7d15f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb20fd6801a875454ddc0b7bac32cc9d8ada2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e17da4e444b33196d4fb85958336a3f5de2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heafe11ebd099b5e70e330bca039131e59f04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb301bd8575344c76590b2fb669fc2f01f6b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46efa8cb826d602d18004b6e0ea30b75a69e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f70beb5d0fcbd093faea803aab5d2fd9dd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0972647ad8bae356859fcfd0bb16ca8ee2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ebc972a35a71245bbe81592075105b45b4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb28ce2fc19dfaacdc9c3c415b117753f2212;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d91c3c569d7566f16d51feb70d927c5a030;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcffd0e41294b22122806f59d186540d4d6c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he84ac595e09749c7a1d0a631961290eaac4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bc9ced7b12a9bb8aff65339f8f64aad81b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc316c5531e81f391fd19f5cbc22966d8220e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20e01d9eb8badcb84fb9d4249e193b87c962;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h861e25fe29d016327268281b7241a4fe4565;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab6567d3b39678ac0377f0a83617f057ce76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecdf2bd600636b90390f78044a091deb207b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h406685535e841f8957c7ac8a28ac8147c005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda1ef3cdf5396c8dce6f744ae95cde6ea14a;
        #1
        $finish();
    end
endmodule
